//
//					\\\ Sapere Aude ///
//
// -----------------------------------------------------------------------------
// Copyright (c) 2014-2020 All rights reserved
// -----------------------------------------------------------------------------
// Author : Angione Francesco s262620@studenti.polito.it franout@Github.com
// File   : tb_cu.sv
// Create : 2020-07-27 15:16:34
// Revise : 2020-07-27 15:18:09
// Editor : sublime text3, tab size (4)
// Description: 
// -----------------------------------------------------------------------------


module tb_cu ();

endmodule