
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, n554, 
      boothmul_pipelined_i_muxes_in_7_233_port, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_201_port, 
      boothmul_pipelined_i_muxes_in_7_200_port, 
      boothmul_pipelined_i_muxes_in_7_199_port, 
      boothmul_pipelined_i_muxes_in_7_198_port, 
      boothmul_pipelined_i_muxes_in_7_197_port, 
      boothmul_pipelined_i_muxes_in_7_196_port, 
      boothmul_pipelined_i_muxes_in_7_195_port, 
      boothmul_pipelined_i_muxes_in_7_194_port, 
      boothmul_pipelined_i_muxes_in_7_193_port, 
      boothmul_pipelined_i_muxes_in_7_192_port, 
      boothmul_pipelined_i_muxes_in_7_191_port, 
      boothmul_pipelined_i_muxes_in_7_190_port, 
      boothmul_pipelined_i_muxes_in_7_189_port, 
      boothmul_pipelined_i_muxes_in_7_188_port, 
      boothmul_pipelined_i_muxes_in_7_187_port, 
      boothmul_pipelined_i_muxes_in_7_186_port, 
      boothmul_pipelined_i_muxes_in_7_77_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_7_47_port, 
      boothmul_pipelined_i_muxes_in_7_46_port, 
      boothmul_pipelined_i_muxes_in_7_45_port, 
      boothmul_pipelined_i_muxes_in_7_44_port, 
      boothmul_pipelined_i_muxes_in_7_43_port, 
      boothmul_pipelined_i_muxes_in_7_42_port, 
      boothmul_pipelined_i_muxes_in_7_41_port, 
      boothmul_pipelined_i_muxes_in_7_40_port, 
      boothmul_pipelined_i_muxes_in_7_39_port, 
      boothmul_pipelined_i_muxes_in_7_38_port, 
      boothmul_pipelined_i_muxes_in_7_37_port, 
      boothmul_pipelined_i_muxes_in_7_36_port, 
      boothmul_pipelined_i_muxes_in_7_35_port, 
      boothmul_pipelined_i_muxes_in_7_34_port, 
      boothmul_pipelined_i_muxes_in_7_33_port, 
      boothmul_pipelined_i_muxes_in_7_32_port, 
      boothmul_pipelined_i_muxes_in_7_31_port, 
      boothmul_pipelined_i_muxes_in_6_219_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_189_port, 
      boothmul_pipelined_i_muxes_in_6_188_port, 
      boothmul_pipelined_i_muxes_in_6_187_port, 
      boothmul_pipelined_i_muxes_in_6_186_port, 
      boothmul_pipelined_i_muxes_in_6_185_port, 
      boothmul_pipelined_i_muxes_in_6_184_port, 
      boothmul_pipelined_i_muxes_in_6_183_port, 
      boothmul_pipelined_i_muxes_in_6_182_port, 
      boothmul_pipelined_i_muxes_in_6_181_port, 
      boothmul_pipelined_i_muxes_in_6_180_port, 
      boothmul_pipelined_i_muxes_in_6_179_port, 
      boothmul_pipelined_i_muxes_in_6_178_port, 
      boothmul_pipelined_i_muxes_in_6_177_port, 
      boothmul_pipelined_i_muxes_in_6_176_port, 
      boothmul_pipelined_i_muxes_in_6_175_port, 
      boothmul_pipelined_i_muxes_in_6_174_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_6_45_port, 
      boothmul_pipelined_i_muxes_in_6_44_port, 
      boothmul_pipelined_i_muxes_in_6_43_port, 
      boothmul_pipelined_i_muxes_in_6_42_port, 
      boothmul_pipelined_i_muxes_in_6_41_port, 
      boothmul_pipelined_i_muxes_in_6_40_port, 
      boothmul_pipelined_i_muxes_in_6_39_port, 
      boothmul_pipelined_i_muxes_in_6_38_port, 
      boothmul_pipelined_i_muxes_in_6_37_port, 
      boothmul_pipelined_i_muxes_in_6_36_port, 
      boothmul_pipelined_i_muxes_in_6_35_port, 
      boothmul_pipelined_i_muxes_in_6_34_port, 
      boothmul_pipelined_i_muxes_in_6_33_port, 
      boothmul_pipelined_i_muxes_in_6_32_port, 
      boothmul_pipelined_i_muxes_in_6_31_port, 
      boothmul_pipelined_i_muxes_in_6_30_port, 
      boothmul_pipelined_i_muxes_in_6_29_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_177_port, 
      boothmul_pipelined_i_muxes_in_5_176_port, 
      boothmul_pipelined_i_muxes_in_5_175_port, 
      boothmul_pipelined_i_muxes_in_5_174_port, 
      boothmul_pipelined_i_muxes_in_5_173_port, 
      boothmul_pipelined_i_muxes_in_5_172_port, 
      boothmul_pipelined_i_muxes_in_5_171_port, 
      boothmul_pipelined_i_muxes_in_5_170_port, 
      boothmul_pipelined_i_muxes_in_5_169_port, 
      boothmul_pipelined_i_muxes_in_5_168_port, 
      boothmul_pipelined_i_muxes_in_5_167_port, 
      boothmul_pipelined_i_muxes_in_5_166_port, 
      boothmul_pipelined_i_muxes_in_5_165_port, 
      boothmul_pipelined_i_muxes_in_5_164_port, 
      boothmul_pipelined_i_muxes_in_5_163_port, 
      boothmul_pipelined_i_muxes_in_5_162_port, 
      boothmul_pipelined_i_muxes_in_5_69_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_5_43_port, 
      boothmul_pipelined_i_muxes_in_5_42_port, 
      boothmul_pipelined_i_muxes_in_5_41_port, 
      boothmul_pipelined_i_muxes_in_5_40_port, 
      boothmul_pipelined_i_muxes_in_5_39_port, 
      boothmul_pipelined_i_muxes_in_5_38_port, 
      boothmul_pipelined_i_muxes_in_5_37_port, 
      boothmul_pipelined_i_muxes_in_5_36_port, 
      boothmul_pipelined_i_muxes_in_5_35_port, 
      boothmul_pipelined_i_muxes_in_5_34_port, 
      boothmul_pipelined_i_muxes_in_5_33_port, 
      boothmul_pipelined_i_muxes_in_5_32_port, 
      boothmul_pipelined_i_muxes_in_5_31_port, 
      boothmul_pipelined_i_muxes_in_5_30_port, 
      boothmul_pipelined_i_muxes_in_5_29_port, 
      boothmul_pipelined_i_muxes_in_5_28_port, 
      boothmul_pipelined_i_muxes_in_5_27_port, 
      boothmul_pipelined_i_muxes_in_4_191_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_165_port, 
      boothmul_pipelined_i_muxes_in_4_164_port, 
      boothmul_pipelined_i_muxes_in_4_163_port, 
      boothmul_pipelined_i_muxes_in_4_162_port, 
      boothmul_pipelined_i_muxes_in_4_161_port, 
      boothmul_pipelined_i_muxes_in_4_160_port, 
      boothmul_pipelined_i_muxes_in_4_159_port, 
      boothmul_pipelined_i_muxes_in_4_158_port, 
      boothmul_pipelined_i_muxes_in_4_157_port, 
      boothmul_pipelined_i_muxes_in_4_156_port, 
      boothmul_pipelined_i_muxes_in_4_155_port, 
      boothmul_pipelined_i_muxes_in_4_154_port, 
      boothmul_pipelined_i_muxes_in_4_153_port, 
      boothmul_pipelined_i_muxes_in_4_152_port, 
      boothmul_pipelined_i_muxes_in_4_151_port, 
      boothmul_pipelined_i_muxes_in_4_150_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_4_41_port, 
      boothmul_pipelined_i_muxes_in_4_40_port, 
      boothmul_pipelined_i_muxes_in_4_39_port, 
      boothmul_pipelined_i_muxes_in_4_38_port, 
      boothmul_pipelined_i_muxes_in_4_37_port, 
      boothmul_pipelined_i_muxes_in_4_36_port, 
      boothmul_pipelined_i_muxes_in_4_35_port, 
      boothmul_pipelined_i_muxes_in_4_34_port, 
      boothmul_pipelined_i_muxes_in_4_33_port, 
      boothmul_pipelined_i_muxes_in_4_32_port, 
      boothmul_pipelined_i_muxes_in_4_31_port, 
      boothmul_pipelined_i_muxes_in_4_30_port, 
      boothmul_pipelined_i_muxes_in_4_29_port, 
      boothmul_pipelined_i_muxes_in_4_28_port, 
      boothmul_pipelined_i_muxes_in_4_27_port, 
      boothmul_pipelined_i_muxes_in_4_26_port, 
      boothmul_pipelined_i_muxes_in_4_25_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_153_port, 
      boothmul_pipelined_i_muxes_in_3_152_port, 
      boothmul_pipelined_i_muxes_in_3_151_port, 
      boothmul_pipelined_i_muxes_in_3_150_port, 
      boothmul_pipelined_i_muxes_in_3_149_port, 
      boothmul_pipelined_i_muxes_in_3_148_port, 
      boothmul_pipelined_i_muxes_in_3_147_port, 
      boothmul_pipelined_i_muxes_in_3_146_port, 
      boothmul_pipelined_i_muxes_in_3_145_port, 
      boothmul_pipelined_i_muxes_in_3_144_port, 
      boothmul_pipelined_i_muxes_in_3_143_port, 
      boothmul_pipelined_i_muxes_in_3_142_port, 
      boothmul_pipelined_i_muxes_in_3_141_port, 
      boothmul_pipelined_i_muxes_in_3_140_port, 
      boothmul_pipelined_i_muxes_in_3_139_port, 
      boothmul_pipelined_i_muxes_in_3_138_port, 
      boothmul_pipelined_i_muxes_in_3_61_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_muxes_in_3_39_port, 
      boothmul_pipelined_i_muxes_in_3_38_port, 
      boothmul_pipelined_i_muxes_in_3_37_port, 
      boothmul_pipelined_i_muxes_in_3_36_port, 
      boothmul_pipelined_i_muxes_in_3_35_port, 
      boothmul_pipelined_i_muxes_in_3_34_port, 
      boothmul_pipelined_i_muxes_in_3_33_port, 
      boothmul_pipelined_i_muxes_in_3_32_port, 
      boothmul_pipelined_i_muxes_in_3_31_port, 
      boothmul_pipelined_i_muxes_in_3_30_port, 
      boothmul_pipelined_i_muxes_in_3_29_port, 
      boothmul_pipelined_i_muxes_in_3_28_port, 
      boothmul_pipelined_i_muxes_in_3_27_port, 
      boothmul_pipelined_i_muxes_in_3_26_port, 
      boothmul_pipelined_i_muxes_in_3_25_port, 
      boothmul_pipelined_i_muxes_in_3_24_port, 
      boothmul_pipelined_i_muxes_in_3_23_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_1_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_6_28_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_5_26_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_4_24_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_3_22_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_7_15_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517_port, n2518_port, n2519_port, n2520_port, n2521_port, n2522_port, 
      n2523_port, n2524_port, n2525_port, n2526_port, n2527_port, n2528_port, 
      n2529_port, n2530_port, n2531_port, n2532_port, n2533_port, n2534_port, 
      n2535_port, n2536_port, n2537_port, n2538_port, n2539_port, n2540_port, 
      n2541_port, n2542_port, n2543_port, n2544_port, n2545_port, n2546_port, 
      n2547_port, n2548_port, n2549, n2550, n2551, n2552, n2553, n2554, n2555, 
      n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, 
      n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, 
      n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
      n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
      n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
      n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, 
      n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
      n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, 
      n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, 
      n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, 
      n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, 
      n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, 
      n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, 
      n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, 
      n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, 
      n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, 
      n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
      n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, 
      n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, 
      n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, 
      n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, 
      n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, 
      n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
      n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
      n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, 
      n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, 
      n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, 
      n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, 
      n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, 
      n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, 
      n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, 
      n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
      n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, 
      n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, 
      n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
      n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, 
      n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, 
      n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, 
      n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, 
      n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, 
      n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
      n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, 
      n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, 
      n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
      n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
      n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
      n3036, n3037, n3038, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526 : std_logic;

begin
   
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n3038, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n3038, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n3038, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n554, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n554, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n554, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n3038, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n554, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n554, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n3038, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n554, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n554, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n554, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n3038, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n554, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n554, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n554, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n554, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n554, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n554, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n554, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n554, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n554, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n554, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n554, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n3038, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n554, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n554, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n3038, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n554, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n3038, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => DATA1(3), GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, QN 
                           => n3019);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3024);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3023);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3021);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3025);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, QN => 
                           n_1060);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => rst_BAR, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3035, CK => clk, RN => rst_BAR, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => rst_BAR, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => rst_BAR, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_219_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_29_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_31_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_218_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_30_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_32_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_217_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_31_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_33_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_216_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_32_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_34_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_215_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_33_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_35_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_214_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_34_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_36_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_213_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_35_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_37_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_212_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_36_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_38_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_211_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_37_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_39_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_210_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_38_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_40_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_209_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_39_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_41_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_208_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_40_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_42_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_207_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_41_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_43_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_42_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_44_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_43_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_45_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_44_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_46_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_45_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_47_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1106);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_175_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_77_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_174_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_186_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_175_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_187_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_176_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_188_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_177_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_189_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_178_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_190_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_179_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_191_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_180_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_192_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_181_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_193_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_182_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_194_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_183_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_195_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_184_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_196_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_185_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_197_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_186_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_198_port, QN => 
                           n_1120);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_187_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_199_port, QN => 
                           n_1121);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_188_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_200_port, QN => 
                           n_1122);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_189_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_201_port, QN => 
                           n_1123);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1124);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1125);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1126);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1127);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1128);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1129);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1130);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1131);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1132);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1133);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_219_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_233_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1156
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3034, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1157
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_9_port, QN => n_1158)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_8_port, QN => n_1159)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_7_port, QN => n_1160)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_6_port, QN => n_1161)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_5_port, QN => n_1162)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_4_port, QN => n_1163)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_3_port, QN => n_1164)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_2_port, QN => n_1165)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_1_port, QN => n_1166)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_0_port, QN => n_1167)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_221_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_27_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_29_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_220_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_28_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_30_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_219_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_29_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_31_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_218_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_30_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_32_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_217_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_31_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_33_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_216_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_32_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_34_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_215_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_33_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_35_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_214_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_34_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_36_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_213_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_35_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_37_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_212_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_36_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_38_port, QN => 
                           n_1177);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_211_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_37_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_39_port, QN => 
                           n_1178);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_210_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_38_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_40_port, QN => 
                           n_1179);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_209_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_39_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_41_port, QN => 
                           n_1180);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_208_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_40_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_42_port, QN => 
                           n_1181);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_207_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_41_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_43_port, QN => 
                           n_1182);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_42_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_44_port, QN => 
                           n_1183);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_43_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_45_port, QN => 
                           n_1184);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => 
                           n_1185);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1186);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1187);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1188);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1189);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1190);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1191);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_69_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_162_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_174_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_163_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_175_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_164_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_176_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_165_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_177_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_166_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_178_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_167_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_179_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_168_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_180_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_169_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_181_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_170_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_182_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_171_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_183_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_172_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_184_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_173_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_185_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_174_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_186_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_175_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_187_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_176_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_188_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_177_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_189_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1231);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1232);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_219_port, QN => 
                           n_1233);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1234);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1235);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1236);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1237);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1238);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1239);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1240);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1241);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1242);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1243);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1244);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1245);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1246);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_10_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_9_port, QN => n_1249)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3033, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1250)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_7_port, QN => n_1251)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_6_port, QN => n_1252)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_5_port, QN => n_1253)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_4_port, QN => n_1254)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_3_port, QN => n_1255)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_2_port, QN => n_1256)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_1_port, QN => n_1257)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_0_port, QN => n_1258)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_223_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_25_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_27_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_222_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_26_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_28_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_221_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_27_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_29_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_220_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_28_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_30_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_219_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_29_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_31_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_218_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_30_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_32_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_217_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_31_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_33_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_216_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_32_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_34_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_215_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_33_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_35_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_214_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_34_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_36_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_213_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_35_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_37_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_212_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_36_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_38_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_211_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_37_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_39_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_210_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_38_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_40_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_209_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_39_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_41_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_208_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_40_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_42_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_207_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_41_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_43_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1282);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1283);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1284);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1285);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1286);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1287);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1288);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1289);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1290);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_69_port, QN => 
                           n_1291);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_150_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_162_port, QN => 
                           n_1292);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_151_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_163_port, QN => 
                           n_1293);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_152_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_164_port, QN => 
                           n_1294);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_153_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_165_port, QN => 
                           n_1295);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_154_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_166_port, QN => 
                           n_1296);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_155_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_167_port, QN => 
                           n_1297);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_156_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_168_port, QN => 
                           n_1298);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_157_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_169_port, QN => 
                           n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_158_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_170_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_159_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_171_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_160_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_172_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_161_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_173_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_162_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_174_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_163_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_175_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_164_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_176_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_165_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_177_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_191_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1332);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1333);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1334);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1335);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1336);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1337);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1338
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, QN => n_1339
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_7_port, QN => n_1340)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3032, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1341)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_5_port, QN => n_1342)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_4_port, QN => n_1343)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_3_port, QN => n_1344)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_2_port, QN => n_1345)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_1_port, QN => n_1346)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_0_port, QN => n_1347)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_225_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_23_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_25_port, QN => 
                           n_1348);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_224_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_24_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_26_port, QN => 
                           n_1349);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_223_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_25_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_27_port, QN => 
                           n_1350);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_222_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_26_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_28_port, QN => 
                           n_1351);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_221_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_27_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_29_port, QN => 
                           n_1352);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_220_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_28_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_30_port, QN => 
                           n_1353);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_219_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_29_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_31_port, QN => 
                           n_1354);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_218_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_30_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_32_port, QN => 
                           n_1355);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_217_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_31_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_33_port, QN => 
                           n_1356);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_216_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_32_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_34_port, QN => 
                           n_1357);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_215_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_33_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_35_port, QN => 
                           n_1358);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_214_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_34_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_36_port, QN => 
                           n_1359);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_213_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_35_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_37_port, QN => 
                           n_1360);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_212_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_36_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_38_port, QN => 
                           n_1361);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_211_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_37_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_39_port, QN => 
                           n_1362);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_210_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_38_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_40_port, QN => 
                           n_1363);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_209_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_39_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_41_port, QN => 
                           n_1364);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => 
                           n_1365);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1366);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1367);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1368);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1369);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1370);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1371);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1372);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1373);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1374);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1375);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1376);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1377);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1378);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1379);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_61_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => 
                           n_1380);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_110_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_138_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_150_port, QN => 
                           n_1381);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_109_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_139_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_151_port, QN => 
                           n_1382);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_108_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_140_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_152_port, QN => 
                           n_1383);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_107_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_141_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_153_port, QN => 
                           n_1384);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_106_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_142_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_154_port, QN => 
                           n_1385);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_105_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_143_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_155_port, QN => 
                           n_1386);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_104_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_144_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_156_port, QN => 
                           n_1387);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_103_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_145_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_157_port, QN => 
                           n_1388);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_102_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_146_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_158_port, QN => 
                           n_1389);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_147_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_159_port, QN => 
                           n_1390);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_148_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_160_port, QN => 
                           n_1391);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_149_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_161_port, QN => 
                           n_1392);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_150_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_162_port, QN => 
                           n_1393);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_151_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_163_port, QN => 
                           n_1394);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_152_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_164_port, QN => 
                           n_1395);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_153_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_165_port, QN => 
                           n_1396);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1397);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1398);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1399);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1400);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1401);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1402);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1403);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1404);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1405);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1406);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1407);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1408);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1409);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1410);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1411);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1412);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_191_port, QN => 
                           n_1413);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1414);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1415);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1416);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1417);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1418);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1419);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1420);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1421);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1422);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1423);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1424);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1425
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1426
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1427
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_6_port, QN => n_1428
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_5_port, QN => n_1429)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3031, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1430)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_3_port, QN => n_1431)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_2_port, QN => n_1432)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_1_port, QN => n_1433)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_0_port, QN => n_1434)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_227_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_23_port, QN => 
                           n_1435);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_226_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_24_port, QN => 
                           n_1436);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_225_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_25_port, QN => 
                           n_1437);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_224_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_26_port, QN => 
                           n_1438);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_223_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_27_port, QN => 
                           n_1439);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_222_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_28_port, QN => 
                           n_1440);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_221_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_29_port, QN => 
                           n_1441);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_220_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_30_port, QN => 
                           n_1442);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_219_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_31_port, QN => 
                           n_1443);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_218_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_32_port, QN => 
                           n_1444);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_217_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_33_port, QN => 
                           n_1445);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_216_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_34_port, QN => 
                           n_1446);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_215_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_35_port, QN => 
                           n_1447);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_214_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_36_port, QN => 
                           n_1448);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_213_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_37_port, QN => 
                           n_1449);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_212_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_38_port, QN => 
                           n_1450);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_211_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_39_port, QN => 
                           n_1451);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => 
                           n_1452);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1453);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1454);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1455);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1456);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1457);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1458);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1459);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1460);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1461);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1462);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1463);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1464);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1465);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1466);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_61_port, QN => 
                           n_1467);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_122_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_138_port, QN => 
                           n_1468);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_121_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_139_port, QN => 
                           n_1469);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_120_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_140_port, QN => 
                           n_1470);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_119_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_141_port, QN => 
                           n_1471);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_118_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_142_port, QN => 
                           n_1472);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_117_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_143_port, QN => 
                           n_1473);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_116_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_144_port, QN => 
                           n_1474);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_115_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_145_port, QN => 
                           n_1475);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_114_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_146_port, QN => 
                           n_1476);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_113_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_147_port, QN => 
                           n_1477);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_112_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_148_port, QN => 
                           n_1478);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_111_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_149_port, QN => 
                           n_1479);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_110_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_150_port, QN => 
                           n_1480);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_109_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_151_port, QN => 
                           n_1481);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_108_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_152_port, QN => 
                           n_1482);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_107_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_153_port, QN => 
                           n_1483);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1484);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1485);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1486);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1487);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1488);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1489);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1490);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1491);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1492);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1493);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1494);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1495);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1496);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1497);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1498);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1499);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1500);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1501);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1502);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1503);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1504);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1505);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1506);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1507);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1508);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1509
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1510
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1511
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1512
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1513
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_4_port, QN => n_1514
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_2_3_port, QN => n_1515)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3037, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1516)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_1_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_2_1_port, QN => n_1517)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_2_0_port, QN => n_1518)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n_1519);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n554, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3036,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1520, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3026,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1521, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3030,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1522, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3029,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1523, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3028
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1524, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3027
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1525, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3020
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1526, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   U3 : INV_X2 port map( A => n2428, ZN => n2170);
   U4 : INV_X2 port map( A => n1068, ZN => n1721);
   U5 : NOR3_X2 port map( A1 => n2476, A2 => n1176, A3 => n1191, ZN => n2469);
   U6 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_7_15_port
                           , A2 => n2961, ZN => n2994);
   U7 : NOR2_X2 port map( A1 => n3025, A2 => n2773, ZN => n2807);
   U8 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_3_7_port,
                           A2 => n2813, ZN => n2845);
   U9 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_4_9_port,
                           A2 => n2850, ZN => n2882);
   U10 : NOR2_X2 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, A2 
                           => n2887, ZN => n2919);
   U11 : NOR2_X2 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, A2 
                           => n2924, ZN => n2956);
   U12 : NOR2_X2 port map( A1 => n2768, A2 => n2734, ZN => n2769);
   U13 : INV_X2 port map( A => n2121, ZN => n2440);
   U14 : NOR2_X2 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, A2 
                           => n1037, ZN => n2992);
   U15 : NOR2_X2 port map( A1 => n3023, A2 => n1040, ZN => n2920);
   U16 : NOR2_X2 port map( A1 => n3021, A2 => n1042, ZN => n2846);
   U17 : NOR2_X2 port map( A1 => n3024, A2 => n1044, ZN => n2957);
   U18 : NOR2_X2 port map( A1 => n3022, A2 => n1046, ZN => n2883);
   U19 : NOR2_X2 port map( A1 => n3019, A2 => n1037, ZN => n2993);
   U20 : NOR2_X2 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, A2 
                           => n1040, ZN => n2921);
   U21 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_3_7_port
                           , A2 => n1042, ZN => n2847);
   U22 : NOR2_X2 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, A2 
                           => n1044, ZN => n2958);
   U23 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_4_9_port
                           , A2 => n1046, ZN => n2884);
   U24 : OAI21_X2 port map( B1 => n2726, B2 => n1315, A => n1963, ZN => n2079);
   U25 : INV_X2 port map( A => n1750, ZN => n2461);
   U26 : INV_X2 port map( A => n1721, ZN => n2434);
   U27 : INV_X2 port map( A => n1678, ZN => n2431);
   U28 : NOR2_X2 port map( A1 => n1066, A2 => n1098, ZN => n2444);
   U29 : OAI21_X2 port map( B1 => n1175, B2 => n1174, A => n1907, ZN => n2472);
   U30 : AOI211_X4 port map( C1 => data2_mul_1_port, C2 => data2_mul_2_port, A 
                           => data2_mul_3_port, B => n2735, ZN => n2763);
   U31 : NOR3_X4 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           A3 => n3024, ZN => n2955);
   U32 : NOR3_X4 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           A3 => n3023, ZN => n2918);
   U33 : NOR3_X4 port map( A1 => boothmul_pipelined_i_multiplicand_pip_4_8_port
                           , A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => n3022, ZN => n2881);
   U34 : NOR3_X4 port map( A1 => boothmul_pipelined_i_multiplicand_pip_3_6_port
                           , A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => n3021, ZN => n2844);
   U35 : AOI211_X4 port map( C1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, C2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => boothmul_pipelined_i_multiplicand_pip_2_5_port, B
                           => n2774, ZN => n2802);
   U36 : NOR3_X4 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           A3 => n3019, ZN => n2995);
   U37 : NOR2_X2 port map( A1 => n1086, A2 => n2121, ZN => n2449);
   U38 : INV_X1 port map( A => n554, ZN => n2696);
   U39 : INV_X1 port map( A => data1_mul_0_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port);
   U40 : CLKBUF_X1 port map( A => n2731, Z => n2721);
   U41 : INV_X1 port map( A => data1_mul_2_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port);
   U42 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n1036);
   U43 : OAI21_X1 port map( B1 => data2_mul_1_port, B2 => data2_mul_2_port, A 
                           => n1036, ZN => n2734);
   U44 : NOR2_X1 port map( A1 => n2734, A2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           ZN => n1053);
   U45 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n3013);
   U46 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN => 
                           n2999);
   U47 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n2733);
   U48 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => n2733, ZN => n3012);
   U49 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n2998);
   U50 : OR2_X1 port map( A1 => n2733, A2 => data2_mul_1_port, ZN => n3018);
   U51 : OAI222_X1 port map( A1 => n3013, A2 => n2999, B1 => n3012, B2 => n2998
                           , C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, 
                           C2 => n3018, ZN => n1054);
   U52 : AND2_X1 port map( A1 => n1053, A2 => n1054, ZN => n3036);
   U53 : INV_X1 port map( A => data1_mul_15_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port);
   U54 : XOR2_X1 port map( A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => boothmul_pipelined_i_muxes_in_0_119_port);
   U55 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           ZN => n2961);
   U56 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           A => n2961, ZN => n1037);
   U57 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_233_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_47_port
                           , ZN => n1038);
   U58 : INV_X1 port map( A => n1038, ZN => n2312);
   U59 : AND2_X1 port map( A1 => n2312, A2 => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, ZN => n3020
                           );
   U60 : NOR2_X1 port map( A1 => FUNC(2), A2 => FUNC(0), ZN => n1063);
   U61 : INV_X1 port map( A => FUNC(1), ZN => n1890);
   U62 : NAND2_X1 port map( A1 => n1063, A2 => n1890, ZN => n554);
   U63 : INV_X1 port map( A => n2696, ZN => n3038);
   U64 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n1039);
   U65 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n1039, ZN => n2773);
   U66 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           A2 => n2773, ZN => n1048);
   U67 : AND2_X1 port map( A1 => n1048, A2 => 
                           boothmul_pipelined_i_sum_B_in_2_4_port, ZN => n3026)
                           ;
   U68 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n2887);
   U69 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, A
                           => n2887, ZN => n1040);
   U70 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_43_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_205_port, ZN
                           => n1041);
   U71 : INV_X1 port map( A => n1041, ZN => n1051);
   U72 : AND2_X1 port map( A1 => n1051, A2 => 
                           boothmul_pipelined_i_sum_B_in_5_10_port, ZN => n3028
                           );
   U73 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n2813);
   U74 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, A
                           => n2813, ZN => n1042);
   U75 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_39_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_177_port, ZN
                           => n1043);
   U76 : INV_X1 port map( A => n1043, ZN => n1049);
   U77 : AND2_X1 port map( A1 => n1049, A2 => 
                           boothmul_pipelined_i_sum_B_in_3_6_port, ZN => n3030)
                           ;
   U78 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n2924);
   U79 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           A => n2924, ZN => n1044);
   U80 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_45_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_219_port, ZN
                           => n1045);
   U81 : INV_X1 port map( A => n1045, ZN => n1052);
   U82 : AND2_X1 port map( A1 => n1052, A2 => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, ZN => n3027
                           );
   U83 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n2850);
   U84 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, A
                           => n2850, ZN => n1046);
   U85 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_41_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_191_port, ZN
                           => n1047);
   U86 : INV_X1 port map( A => n1047, ZN => n1050);
   U87 : AND2_X1 port map( A1 => n1050, A2 => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, ZN => n3029)
                           ;
   U88 : INV_X1 port map( A => data1_mul_1_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port);
   U89 : INV_X1 port map( A => data1_mul_3_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port);
   U90 : INV_X1 port map( A => data1_mul_4_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port);
   U91 : INV_X1 port map( A => data1_mul_5_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port);
   U92 : INV_X1 port map( A => data1_mul_6_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port);
   U93 : INV_X1 port map( A => data1_mul_7_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port);
   U94 : INV_X1 port map( A => data1_mul_8_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port);
   U95 : INV_X1 port map( A => data1_mul_9_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port);
   U96 : INV_X1 port map( A => data1_mul_10_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port);
   U97 : INV_X1 port map( A => data1_mul_11_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port);
   U98 : INV_X1 port map( A => data1_mul_12_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port);
   U99 : INV_X1 port map( A => data1_mul_13_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port);
   U100 : INV_X1 port map( A => data1_mul_14_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port);
   U101 : INV_X1 port map( A => FUNC(2), ZN => n2682);
   U102 : NOR2_X1 port map( A1 => n2682, A2 => FUNC(0), ZN => n1064);
   U103 : AND2_X1 port map( A1 => n1890, A2 => n1064, ZN => n1238);
   U104 : INV_X1 port map( A => FUNC(3), ZN => n2695);
   U105 : NAND2_X1 port map( A1 => n1238, A2 => n2695, ZN => n553);
   U106 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_2_4_port, B => 
                           n1048, Z => n3031);
   U107 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, B => 
                           n1049, Z => n3032);
   U108 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_4_8_port, B => 
                           n1050, Z => n3033);
   U109 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_5_10_port, B => 
                           n1051, Z => n3034);
   U110 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_6_12_port, B => 
                           n1052, Z => n3035);
   U111 : XOR2_X1 port map( A => n1054, B => n1053, Z => n3037);
   U112 : NOR4_X1 port map( A1 => DATA2(6), A2 => DATA2(7), A3 => DATA2(8), A4 
                           => DATA2(9), ZN => n1062);
   U113 : INV_X1 port map( A => DATA2(0), ZN => n2730);
   U114 : INV_X1 port map( A => DATA2(1), ZN => n2729);
   U115 : NAND2_X1 port map( A1 => n2730, A2 => n2729, ZN => n1175);
   U116 : INV_X1 port map( A => n1175, ZN => n1436);
   U117 : INV_X1 port map( A => DATA2(3), ZN => n2727);
   U118 : INV_X1 port map( A => DATA2(5), ZN => n2725);
   U119 : INV_X1 port map( A => DATA2(4), ZN => n2726);
   U120 : NAND2_X1 port map( A1 => n2725, A2 => n2726, ZN => n1907);
   U121 : INV_X1 port map( A => n1907, ZN => n2467);
   U122 : NAND2_X1 port map( A1 => n2727, A2 => n2467, ZN => n1086);
   U123 : NOR2_X1 port map( A1 => n1086, A2 => DATA2(2), ZN => n1518);
   U124 : CLKBUF_X1 port map( A => n1518, Z => n1678);
   U125 : NAND2_X1 port map( A1 => n1436, A2 => n1678, ZN => n2428);
   U126 : INV_X1 port map( A => DATA2(10), ZN => n2718);
   U127 : INV_X1 port map( A => DATA2(11), ZN => n2717);
   U128 : INV_X1 port map( A => DATA2(12), ZN => n2716);
   U129 : INV_X1 port map( A => DATA2(13), ZN => n2715);
   U130 : NAND4_X1 port map( A1 => n2718, A2 => n2717, A3 => n2716, A4 => n2715
                           , ZN => n1055);
   U131 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n2428, A4 
                           => n1055, ZN => n1061);
   U132 : NOR4_X1 port map( A1 => DATA1(15), A2 => DATA1(14), A3 => DATA1(13), 
                           A4 => DATA1(12), ZN => n1059);
   U133 : NOR4_X1 port map( A1 => DATA1(11), A2 => DATA1(10), A3 => DATA1(9), 
                           A4 => DATA1(8), ZN => n1058);
   U134 : NOR4_X1 port map( A1 => DATA1(7), A2 => DATA1(6), A3 => DATA1(5), A4 
                           => DATA1(4), ZN => n1057);
   U135 : NOR4_X1 port map( A1 => DATA1(3), A2 => DATA1(2), A3 => DATA1(1), A4 
                           => DATA1(0), ZN => n1056);
   U136 : AND4_X1 port map( A1 => n1059, A2 => n1058, A3 => n1057, A4 => n1056,
                           ZN => n1060);
   U137 : AOI211_X1 port map( C1 => n1062, C2 => n1061, A => n1060, B => n553, 
                           ZN => n1434);
   U138 : CLKBUF_X1 port map( A => n1434, Z => n2422);
   U139 : NAND2_X1 port map( A1 => FUNC(1), A2 => n1063, ZN => n2416);
   U140 : INV_X1 port map( A => n2416, ZN => n2393);
   U141 : INV_X1 port map( A => DATA2(9), ZN => n2719);
   U142 : NOR2_X1 port map( A1 => n2719, A2 => DATA1(9), ZN => n2626);
   U143 : INV_X1 port map( A => n2626, ZN => n2564);
   U144 : NAND2_X1 port map( A1 => DATA1(9), A2 => n2719, ZN => n2627);
   U145 : NAND2_X1 port map( A1 => n2564, A2 => n2627, ZN => n2520_port);
   U146 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_9_port, B1 => n2393
                           , B2 => n2520_port, ZN => n1256);
   U147 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(4), ZN => n1384);
   U148 : NOR2_X1 port map( A1 => n2729, A2 => n2727, ZN => n1066);
   U149 : INV_X1 port map( A => n1066, ZN => n1089);
   U150 : NOR2_X1 port map( A1 => n1384, A2 => n1089, ZN => n2507);
   U151 : NAND2_X1 port map( A1 => n1064, A2 => n2725, ZN => n1887);
   U152 : AOI211_X1 port map( C1 => n2507, C2 => DATA2(0), A => n1890, B => 
                           n1887, ZN => n1250);
   U153 : NAND2_X1 port map( A1 => FUNC(3), A2 => n1250, ZN => n2409);
   U154 : INV_X1 port map( A => n2409, ZN => n2688);
   U155 : NAND2_X1 port map( A1 => n1907, A2 => DATA2(3), ZN => n1961);
   U156 : NAND2_X1 port map( A1 => n2729, A2 => n1961, ZN => n1065);
   U157 : NAND2_X1 port map( A1 => n1384, A2 => n1961, ZN => n2476);
   U158 : NOR2_X1 port map( A1 => n2730, A2 => n1384, ZN => n1276);
   U159 : AOI21_X1 port map( B1 => n1065, B2 => n2476, A => n1276, ZN => n2481)
                           ;
   U160 : INV_X1 port map( A => n2481, ZN => n2375);
   U161 : NOR2_X1 port map( A1 => n2730, A2 => n1089, ZN => n1385);
   U162 : AOI21_X1 port map( B1 => DATA2(2), B2 => n1385, A => n1907, ZN => 
                           n1219);
   U163 : INV_X1 port map( A => n1219, ZN => n2463);
   U164 : NAND2_X1 port map( A1 => n2463, A2 => n2467, ZN => n2465);
   U165 : INV_X1 port map( A => DATA2(2), ZN => n2728);
   U166 : OAI21_X1 port map( B1 => n2727, B2 => n2728, A => n2467, ZN => n1098)
                           ;
   U167 : INV_X1 port map( A => n2444, ZN => n1896);
   U168 : INV_X1 port map( A => n1086, ZN => n1067);
   U169 : OAI21_X1 port map( B1 => n2729, B2 => n2728, A => n1067, ZN => n1068)
                           ;
   U170 : AOI21_X1 port map( B1 => DATA2(2), B2 => DATA2(0), A => n2434, ZN => 
                           n2176);
   U171 : INV_X1 port map( A => n2176, ZN => n2049);
   U172 : NAND3_X1 port map( A1 => n2730, A2 => DATA2(1), A3 => n1678, ZN => 
                           n1991);
   U173 : INV_X1 port map( A => DATA1(22), ZN => n2126);
   U174 : NOR2_X1 port map( A1 => n1991, A2 => n2126, ZN => n1520);
   U175 : NAND3_X1 port map( A1 => n2729, A2 => DATA2(0), A3 => n1518, ZN => 
                           n1937);
   U176 : INV_X1 port map( A => n1937, ZN => n2205);
   U177 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(21), ZN => n1513);
   U178 : NAND2_X1 port map( A1 => DATA1(20), A2 => n2170, ZN => n1500);
   U179 : OR3_X1 port map( A1 => n2730, A2 => n2729, A3 => n2431, ZN => n1660);
   U180 : INV_X1 port map( A => n1660, ZN => n2005);
   U181 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(23), ZN => n1547);
   U182 : NAND2_X1 port map( A1 => DATA1(24), A2 => n2431, ZN => n1069);
   U183 : NAND4_X1 port map( A1 => n1513, A2 => n1500, A3 => n1547, A4 => n1069
                           , ZN => n1070);
   U184 : NOR2_X1 port map( A1 => n1520, A2 => n1070, ZN => n1084);
   U185 : NOR4_X1 port map( A1 => n2728, A2 => n2730, A3 => n1086, A4 => 
                           DATA2(1), ZN => n1614);
   U186 : CLKBUF_X1 port map( A => n1614, Z => n2436);
   U187 : INV_X1 port map( A => n2436, ZN => n1723);
   U188 : INV_X1 port map( A => DATA1(23), ZN => n2093);
   U189 : NOR2_X1 port map( A1 => n1991, A2 => n2093, ZN => n1526);
   U190 : INV_X1 port map( A => DATA1(21), ZN => n2652);
   U191 : NOR2_X1 port map( A1 => n2428, A2 => n2652, ZN => n1495);
   U192 : AOI211_X1 port map( C1 => DATA1(25), C2 => n2431, A => n1526, B => 
                           n1495, ZN => n1071);
   U193 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(22), ZN => n1509);
   U194 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(24), ZN => n1557);
   U195 : AND3_X1 port map( A1 => n1071, A2 => n1509, A3 => n1557, ZN => n1105)
                           ;
   U196 : INV_X1 port map( A => n1660, ZN => n1801);
   U197 : INV_X1 port map( A => DATA1(24), ZN => n2661);
   U198 : NOR2_X1 port map( A1 => n1991, A2 => n2661, ZN => n1549);
   U199 : INV_X1 port map( A => DATA1(26), ZN => n2512);
   U200 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(23), ZN => n1516);
   U201 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(22), ZN => n1512);
   U202 : OAI211_X1 port map( C1 => n1678, C2 => n2512, A => n1516, B => n1512,
                           ZN => n1072);
   U203 : AOI211_X1 port map( C1 => DATA1(25), C2 => n1801, A => n1549, B => 
                           n1072, ZN => n1110);
   U204 : OAI222_X1 port map( A1 => n2049, A2 => n1084, B1 => n1723, B2 => 
                           n1105, C1 => n1721, C2 => n1110, ZN => n1197);
   U205 : OAI21_X1 port map( B1 => n1086, B2 => DATA2(0), A => n2434, ZN => 
                           n1745);
   U206 : CLKBUF_X1 port map( A => n1745, Z => n2121);
   U207 : INV_X1 port map( A => n1991, ZN => n2006);
   U208 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(20), ZN => n1514);
   U209 : NAND2_X1 port map( A1 => DATA1(21), A2 => n2005, ZN => n1517);
   U210 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(18), ZN => n1073);
   U211 : AND3_X1 port map( A1 => n1514, A2 => n1517, A3 => n1073, ZN => n1074)
                           ;
   U212 : NAND2_X1 port map( A1 => DATA1(19), A2 => n2205, ZN => n1501);
   U213 : OAI211_X1 port map( C1 => n1518, C2 => n2126, A => n1074, B => n1501,
                           ZN => n1075);
   U214 : INV_X1 port map( A => n1075, ZN => n1083);
   U215 : INV_X1 port map( A => DATA1(16), ZN => n2643);
   U216 : NOR2_X1 port map( A1 => n2428, A2 => n2643, ZN => n1077);
   U217 : INV_X1 port map( A => DATA1(20), ZN => n2653);
   U218 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(17), ZN => n1471);
   U219 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(18), ZN => n1502);
   U220 : OAI211_X1 port map( C1 => n1678, C2 => n2653, A => n1471, B => n1502,
                           ZN => n1076);
   U221 : AOI211_X1 port map( C1 => n2005, C2 => DATA1(19), A => n1077, B => 
                           n1076, ZN => n1095);
   U222 : INV_X1 port map( A => DATA1(17), ZN => n2253);
   U223 : NOR2_X1 port map( A1 => n2428, A2 => n2253, ZN => n1079);
   U224 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(18), ZN => n1491);
   U225 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(19), ZN => n1498);
   U226 : OAI211_X1 port map( C1 => n1678, C2 => n2652, A => n1491, B => n1498,
                           ZN => n1078);
   U227 : AOI211_X1 port map( C1 => n2005, C2 => DATA1(20), A => n1079, B => 
                           n1078, ZN => n1094);
   U228 : OAI222_X1 port map( A1 => n1083, A2 => n1721, B1 => n1095, B2 => 
                           n2049, C1 => n1094, C2 => n1723, ZN => n1122);
   U229 : INV_X1 port map( A => n1122, ZN => n1147);
   U230 : CLKBUF_X1 port map( A => n2176, Z => n2438);
   U231 : INV_X1 port map( A => n2438, ZN => n1725);
   U232 : INV_X1 port map( A => n2436, ZN => n2047);
   U233 : NAND2_X1 port map( A1 => DATA1(19), A2 => n2170, ZN => n1490);
   U234 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(20), ZN => n1497);
   U235 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(21), ZN => n1510);
   U236 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(22), ZN => n1524);
   U237 : AND3_X1 port map( A1 => n1497, A2 => n1510, A3 => n1524, ZN => n1080)
                           ;
   U238 : OAI211_X1 port map( C1 => n2093, C2 => n1518, A => n1490, B => n1080,
                           ZN => n1081);
   U239 : INV_X1 port map( A => n1081, ZN => n1085);
   U240 : OAI222_X1 port map( A1 => n1725, A2 => n1083, B1 => n2047, B2 => 
                           n1085, C1 => n1721, C2 => n1084, ZN => n1111);
   U241 : INV_X1 port map( A => n1111, ZN => n1082);
   U242 : NOR4_X1 port map( A1 => n2727, A2 => n1907, A3 => n1175, A4 => 
                           DATA2(2), ZN => n1762);
   U243 : CLKBUF_X1 port map( A => n1762, Z => n2125);
   U244 : INV_X1 port map( A => n2125, ZN => n2442);
   U245 : OAI22_X1 port map( A1 => n2440, A2 => n1147, B1 => n1082, B2 => n2442
                           , ZN => n1088);
   U246 : OAI222_X1 port map( A1 => n1085, A2 => n1721, B1 => n1094, B2 => 
                           n2049, C1 => n1083, C2 => n1723, ZN => n1121);
   U247 : INV_X1 port map( A => n1121, ZN => n1108);
   U248 : INV_X1 port map( A => n2449, ZN => n2178);
   U249 : CLKBUF_X1 port map( A => n2178, Z => n1687);
   U250 : OAI222_X1 port map( A1 => n1105, A2 => n1721, B1 => n1085, B2 => 
                           n2049, C1 => n1084, C2 => n2047, ZN => n1112);
   U251 : INV_X1 port map( A => n1112, ZN => n1132);
   U252 : NAND3_X1 port map( A1 => n1175, A2 => n1086, A3 => n2444, ZN => n2446
                           );
   U253 : OAI22_X1 port map( A1 => n1108, A2 => n1687, B1 => n1132, B2 => n2446
                           , ZN => n1087);
   U254 : AOI211_X1 port map( C1 => n1896, C2 => n1197, A => n1088, B => n1087,
                           ZN => n1212);
   U255 : NAND3_X1 port map( A1 => DATA2(0), A2 => DATA2(2), A3 => DATA2(3), ZN
                           => n1103);
   U256 : OAI21_X1 port map( B1 => n2728, B2 => n1089, A => n2467, ZN => n1102)
                           ;
   U257 : INV_X1 port map( A => n1102, ZN => n2456);
   U258 : NAND3_X1 port map( A1 => n1103, A2 => n2456, A3 => n1098, ZN => n2452
                           );
   U259 : OR2_X1 port map( A1 => n1385, A2 => n1098, ZN => n2454);
   U260 : INV_X1 port map( A => n2454, ZN => n1641);
   U261 : INV_X1 port map( A => DATA1(14), ZN => n2532_port);
   U262 : NOR2_X1 port map( A1 => n2428, A2 => n2532_port, ZN => n1091);
   U263 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(16), ZN => n1472);
   U264 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(15), ZN => n1482);
   U265 : OAI211_X1 port map( C1 => n1660, C2 => n2253, A => n1472, B => n1482,
                           ZN => n1090);
   U266 : AOI211_X1 port map( C1 => DATA1(18), C2 => n2431, A => n1091, B => 
                           n1090, ZN => n1142);
   U267 : NAND2_X1 port map( A1 => DATA1(19), A2 => n2431, ZN => n1092);
   U268 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(17), ZN => n1492);
   U269 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(16), ZN => n1476);
   U270 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(15), ZN => n1487);
   U271 : NAND4_X1 port map( A1 => n1092, A2 => n1492, A3 => n1476, A4 => n1487
                           , ZN => n1093);
   U272 : AOI21_X1 port map( B1 => n2005, B2 => DATA1(18), A => n1093, ZN => 
                           n1120);
   U273 : OAI222_X1 port map( A1 => n1725, A2 => n1142, B1 => n2047, B2 => 
                           n1120, C1 => n1721, C2 => n1095, ZN => n1167);
   U274 : INV_X1 port map( A => n1167, ZN => n1125);
   U275 : OAI22_X1 port map( A1 => n2440, A2 => n1125, B1 => n1147, B2 => n2442
                           , ZN => n1097);
   U276 : OAI222_X1 port map( A1 => n1725, A2 => n1120, B1 => n2047, B2 => 
                           n1095, C1 => n1721, C2 => n1094, ZN => n1157);
   U277 : INV_X1 port map( A => n1157, ZN => n1099);
   U278 : OAI22_X1 port map( A1 => n1099, A2 => n1687, B1 => n1108, B2 => n2446
                           , ZN => n1096);
   U279 : AOI211_X1 port map( C1 => n1896, C2 => n1111, A => n1097, B => n1096,
                           ZN => n1172);
   U280 : INV_X1 port map( A => n1172, ZN => n1158);
   U281 : OR2_X1 port map( A1 => n1098, A2 => n1641, ZN => n1750);
   U282 : INV_X1 port map( A => n2446, ZN => n2183);
   U283 : OAI22_X1 port map( A1 => n2440, A2 => n1099, B1 => n1108, B2 => n2442
                           , ZN => n1101);
   U284 : OAI22_X1 port map( A1 => n2444, A2 => n1132, B1 => n1147, B2 => n1687
                           , ZN => n1100);
   U285 : AOI211_X1 port map( C1 => n2183, C2 => n1111, A => n1101, B => n1100,
                           ZN => n1128);
   U286 : INV_X1 port map( A => n1128, ZN => n1159);
   U287 : AOI22_X1 port map( A1 => n1641, A2 => n1158, B1 => n2461, B2 => n1159
                           , ZN => n1116);
   U288 : CLKBUF_X1 port map( A => n1102, Z => n1902);
   U289 : NOR2_X1 port map( A1 => n1902, A2 => n1103, ZN => n2332);
   U290 : INV_X1 port map( A => n2332, ZN => n2458);
   U291 : INV_X1 port map( A => n2458, ZN => n1823);
   U292 : AOI22_X1 port map( A1 => n2125, A2 => n1112, B1 => n2449, B2 => n1111
                           , ZN => n1107);
   U293 : INV_X1 port map( A => DATA1(25), ZN => n2668);
   U294 : NOR2_X1 port map( A1 => n1991, A2 => n2668, ZN => n1559);
   U295 : INV_X1 port map( A => DATA1(27), ZN => n2025);
   U296 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(24), ZN => n1523);
   U297 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(23), ZN => n1508);
   U298 : OAI211_X1 port map( C1 => n1518, C2 => n2025, A => n1523, B => n1508,
                           ZN => n1104);
   U299 : AOI211_X1 port map( C1 => DATA1(26), C2 => n1801, A => n1559, B => 
                           n1104, ZN => n1131);
   U300 : OAI222_X1 port map( A1 => n1725, A2 => n1105, B1 => n2047, B2 => 
                           n1110, C1 => n1721, C2 => n1131, ZN => n1205);
   U301 : AOI22_X1 port map( A1 => n2183, A2 => n1197, B1 => n1896, B2 => n1205
                           , ZN => n1106);
   U302 : OAI211_X1 port map( C1 => n2440, C2 => n1108, A => n1107, B => n1106,
                           ZN => n1214);
   U303 : AOI22_X1 port map( A1 => DATA1(24), A2 => n2170, B1 => DATA1(28), B2 
                           => n2431, ZN => n1109);
   U304 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(25), ZN => n1546);
   U305 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(26), ZN => n1581);
   U306 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(27), ZN => n1677);
   U307 : AND4_X1 port map( A1 => n1109, A2 => n1546, A3 => n1581, A4 => n1677,
                           ZN => n1196);
   U308 : OAI222_X1 port map( A1 => n1196, A2 => n1721, B1 => n1110, B2 => 
                           n2049, C1 => n1131, C2 => n2047, ZN => n2120);
   U309 : INV_X1 port map( A => n2120, ZN => n1133);
   U310 : AOI22_X1 port map( A1 => n2125, A2 => n1197, B1 => n2121, B2 => n1111
                           , ZN => n1114);
   U311 : AOI22_X1 port map( A1 => n2183, A2 => n1205, B1 => n2449, B2 => n1112
                           , ZN => n1113);
   U312 : OAI211_X1 port map( C1 => n2444, C2 => n1133, A => n1114, B => n1113,
                           ZN => n2239);
   U313 : AOI22_X1 port map( A1 => n1823, A2 => n1214, B1 => n1902, B2 => n2239
                           , ZN => n1115);
   U314 : OAI211_X1 port map( C1 => n1212, C2 => n2452, A => n1116, B => n1115,
                           ZN => n1220);
   U315 : INV_X1 port map( A => n1220, ZN => n1190);
   U316 : AOI22_X1 port map( A1 => n2205, A2 => DATA1(14), B1 => n2005, B2 => 
                           DATA1(16), ZN => n1119);
   U317 : NAND2_X1 port map( A1 => DATA1(17), A2 => n2431, ZN => n1118);
   U318 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(15), ZN => n1477);
   U319 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(13), ZN => n1117);
   U320 : NAND4_X1 port map( A1 => n1119, A2 => n1118, A3 => n1477, A4 => n1117
                           , ZN => n1153);
   U321 : INV_X1 port map( A => n1153, ZN => n1143);
   U322 : OAI222_X1 port map( A1 => n1725, A2 => n1143, B1 => n2047, B2 => 
                           n1142, C1 => n1721, C2 => n1120, ZN => n1182);
   U323 : AOI22_X1 port map( A1 => n1762, A2 => n1157, B1 => n1745, B2 => n1182
                           , ZN => n1124);
   U324 : CLKBUF_X1 port map( A => n2183, Z => n1761);
   U325 : AOI22_X1 port map( A1 => n1761, A2 => n1122, B1 => n1896, B2 => n1121
                           , ZN => n1123);
   U326 : OAI211_X1 port map( C1 => n1125, C2 => n2178, A => n1124, B => n1123,
                           ZN => n1183);
   U327 : INV_X1 port map( A => n1183, ZN => n1162);
   U328 : OAI22_X1 port map( A1 => n1162, A2 => n2454, B1 => n1172, B2 => n1750
                           , ZN => n1127);
   U329 : OAI22_X1 port map( A1 => n1128, A2 => n2452, B1 => n1212, B2 => n2458
                           , ZN => n1126);
   U330 : AOI211_X1 port map( C1 => n1902, C2 => n1214, A => n1127, B => n1126,
                           ZN => n1189);
   U331 : INV_X1 port map( A => n2452, ZN => n2342);
   U332 : INV_X1 port map( A => n2239, ZN => n1217);
   U333 : OAI22_X1 port map( A1 => n1128, A2 => n2454, B1 => n1217, B2 => n2458
                           , ZN => n1138);
   U334 : AOI22_X1 port map( A1 => DATA1(25), A2 => n2170, B1 => DATA1(29), B2 
                           => n2431, ZN => n1130);
   U335 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(26), ZN => n1556);
   U336 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(27), ZN => n1594);
   U337 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(28), ZN => n1129);
   U338 : AND4_X1 port map( A1 => n1130, A2 => n1556, A3 => n1594, A4 => n1129,
                           ZN => n1204);
   U339 : OAI222_X1 port map( A1 => n1204, A2 => n1721, B1 => n1131, B2 => 
                           n2049, C1 => n1196, C2 => n2047, ZN => n2122);
   U340 : INV_X1 port map( A => n2122, ZN => n1200);
   U341 : OAI22_X1 port map( A1 => n2444, A2 => n1200, B1 => n2440, B2 => n1132
                           , ZN => n1136);
   U342 : INV_X1 port map( A => n1205, ZN => n1134);
   U343 : OAI22_X1 port map( A1 => n1134, A2 => n2442, B1 => n1133, B2 => n2446
                           , ZN => n1135);
   U344 : AOI211_X1 port map( C1 => n2449, C2 => n1197, A => n1136, B => n1135,
                           ZN => n1201);
   U345 : OAI22_X1 port map( A1 => n2456, A2 => n1201, B1 => n1212, B2 => n1750
                           , ZN => n1137);
   U346 : AOI211_X1 port map( C1 => n2342, C2 => n1214, A => n1138, B => n1137,
                           ZN => n1218);
   U347 : OAI222_X1 port map( A1 => n2465, A2 => n1190, B1 => n2463, B2 => 
                           n1189, C1 => n1218, C2 => n2467, ZN => n2348);
   U348 : INV_X1 port map( A => DATA1(15), ZN => n2531_port);
   U349 : NOR2_X1 port map( A1 => n1660, A2 => n2531_port, ZN => n1474);
   U350 : NOR2_X1 port map( A1 => n1991, A2 => n2532_port, ZN => n1484);
   U351 : NOR2_X1 port map( A1 => n1474, A2 => n1484, ZN => n1141);
   U352 : NAND2_X1 port map( A1 => DATA1(16), A2 => n2431, ZN => n1140);
   U353 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(13), ZN => n1571);
   U354 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(12), ZN => n1139);
   U355 : NAND4_X1 port map( A1 => n1141, A2 => n1140, A3 => n1571, A4 => n1139
                           , ZN => n1166);
   U356 : INV_X1 port map( A => n1166, ZN => n1144);
   U357 : OAI222_X1 port map( A1 => n1725, A2 => n1144, B1 => n2047, B2 => 
                           n1143, C1 => n1721, C2 => n1142, ZN => n1264);
   U358 : AOI22_X1 port map( A1 => n2125, A2 => n1167, B1 => n1745, B2 => n1264
                           , ZN => n1146);
   U359 : AOI22_X1 port map( A1 => n2183, A2 => n1157, B1 => n2449, B2 => n1182
                           , ZN => n1145);
   U360 : OAI211_X1 port map( C1 => n2444, C2 => n1147, A => n1146, B => n1145,
                           ZN => n1265);
   U361 : AOI22_X1 port map( A1 => n1641, A2 => n1265, B1 => n2461, B2 => n1183
                           , ZN => n1149);
   U362 : AOI22_X1 port map( A1 => n2342, A2 => n1158, B1 => n2332, B2 => n1159
                           , ZN => n1148);
   U363 : OAI211_X1 port map( C1 => n2456, C2 => n1212, A => n1149, B => n1148,
                           ZN => n1150);
   U364 : INV_X1 port map( A => n1150, ZN => n1188);
   U365 : INV_X1 port map( A => DATA1(11), ZN => n2366);
   U366 : NOR2_X1 port map( A1 => n2428, A2 => n2366, ZN => n1151);
   U367 : NOR2_X1 port map( A1 => n1660, A2 => n2532_port, ZN => n1479);
   U368 : AOI211_X1 port map( C1 => DATA1(15), C2 => n2431, A => n1151, B => 
                           n1479, ZN => n1152);
   U369 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(13), ZN => n1488);
   U370 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(12), ZN => n1612);
   U371 : NAND3_X1 port map( A1 => n1152, A2 => n1488, A3 => n1612, ZN => n1178
                           );
   U372 : AOI222_X1 port map( A1 => n1153, A2 => n2434, B1 => n1178, B2 => 
                           n2438, C1 => n1166, C2 => n2436, ZN => n1302);
   U373 : INV_X1 port map( A => n1264, ZN => n1179);
   U374 : OAI22_X1 port map( A1 => n2440, A2 => n1302, B1 => n1179, B2 => n1687
                           , ZN => n1156);
   U375 : AOI22_X1 port map( A1 => n1182, A2 => n2125, B1 => n1167, B2 => n1761
                           , ZN => n1154);
   U376 : INV_X1 port map( A => n1154, ZN => n1155);
   U377 : AOI211_X1 port map( C1 => n1896, C2 => n1157, A => n1156, B => n1155,
                           ZN => n1305);
   U378 : INV_X1 port map( A => n1305, ZN => n1266);
   U379 : INV_X1 port map( A => n2454, ZN => n2397);
   U380 : AOI22_X1 port map( A1 => n1266, A2 => n2397, B1 => n1265, B2 => n2461
                           , ZN => n1161);
   U381 : AOI22_X1 port map( A1 => n1902, A2 => n1159, B1 => n1158, B2 => n2332
                           , ZN => n1160);
   U382 : OAI211_X1 port map( C1 => n2452, C2 => n1162, A => n1161, B => n1160,
                           ZN => n1163);
   U383 : INV_X1 port map( A => n1163, ZN => n1187);
   U384 : INV_X1 port map( A => DATA1(10), ZN => n2516);
   U385 : NOR2_X1 port map( A1 => n2428, A2 => n2516, ZN => n1662);
   U386 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(13), ZN => n1481);
   U387 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(12), ZN => n1570);
   U388 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(11), ZN => n1631);
   U389 : NAND3_X1 port map( A1 => n1481, A2 => n1570, A3 => n1631, ZN => n1164
                           );
   U390 : AOI211_X1 port map( C1 => DATA1(14), C2 => n2431, A => n1662, B => 
                           n1164, ZN => n1165);
   U391 : INV_X1 port map( A => n1165, ZN => n1260);
   U392 : AOI222_X1 port map( A1 => n2176, A2 => n1260, B1 => n2436, B2 => 
                           n1178, C1 => n2434, C2 => n1166, ZN => n1261);
   U393 : INV_X1 port map( A => n1261, ZN => n1337);
   U394 : AOI22_X1 port map( A1 => n2125, A2 => n1264, B1 => n2121, B2 => n1337
                           , ZN => n1169);
   U395 : AOI22_X1 port map( A1 => n1761, A2 => n1182, B1 => n1896, B2 => n1167
                           , ZN => n1168);
   U396 : OAI211_X1 port map( C1 => n1302, C2 => n1687, A => n1169, B => n1168,
                           ZN => n1340);
   U397 : AOI22_X1 port map( A1 => n1641, A2 => n1340, B1 => n2342, B2 => n1265
                           , ZN => n1171);
   U398 : AOI22_X1 port map( A1 => n2461, A2 => n1266, B1 => n2332, B2 => n1183
                           , ZN => n1170);
   U399 : OAI211_X1 port map( C1 => n2456, C2 => n1172, A => n1171, B => n1170,
                           ZN => n1173);
   U400 : INV_X1 port map( A => n1173, ZN => n1270);
   U401 : OAI222_X1 port map( A1 => n1188, A2 => n2467, B1 => n1187, B2 => 
                           n2465, C1 => n1270, C2 => n2463, ZN => n1342);
   U402 : INV_X1 port map( A => n1342, ZN => n1312);
   U403 : NAND2_X1 port map( A1 => n2728, A2 => n2727, ZN => n1174);
   U404 : OAI21_X1 port map( B1 => n1174, B2 => DATA2(1), A => n1907, ZN => 
                           n1176);
   U405 : INV_X1 port map( A => n2472, ZN => n2283);
   U406 : NAND2_X1 port map( A1 => n1176, A2 => n2283, ZN => n2254);
   U407 : OAI222_X1 port map( A1 => n2465, A2 => n1188, B1 => n2463, B2 => 
                           n1187, C1 => n1189, C2 => n2467, ZN => n1309);
   U408 : INV_X1 port map( A => n1309, ZN => n1272);
   U409 : NOR3_X1 port map( A1 => n2730, A2 => n2726, A3 => n2729, ZN => n1191)
                           ;
   U410 : INV_X1 port map( A => n2469, ZN => n2230);
   U411 : OAI22_X1 port map( A1 => n1312, A2 => n2254, B1 => n1272, B2 => n2230
                           , ZN => n1193);
   U412 : INV_X1 port map( A => DATA1(13), ZN => n2602);
   U413 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(12), ZN => n1486);
   U414 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(11), ZN => n1611);
   U415 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(10), ZN => n1645);
   U416 : AND3_X1 port map( A1 => n1486, A2 => n1611, A3 => n1645, ZN => n1177)
                           ;
   U417 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(9), ZN => n1239);
   U418 : OAI211_X1 port map( C1 => n1518, C2 => n2602, A => n1177, B => n1239,
                           ZN => n1301);
   U419 : AOI222_X1 port map( A1 => n1178, A2 => n2434, B1 => n1301, B2 => 
                           n2176, C1 => n1260, C2 => n2436, ZN => n1367);
   U420 : OAI22_X1 port map( A1 => n2440, A2 => n1367, B1 => n1302, B2 => n2442
                           , ZN => n1181);
   U421 : OAI22_X1 port map( A1 => n1261, A2 => n1687, B1 => n1179, B2 => n2446
                           , ZN => n1180);
   U422 : AOI211_X1 port map( C1 => n1896, C2 => n1182, A => n1181, B => n1180,
                           ZN => n1370);
   U423 : OAI22_X1 port map( A1 => n2454, A2 => n1370, B1 => n2452, B2 => n1305
                           , ZN => n1186);
   U424 : AOI22_X1 port map( A1 => n1823, A2 => n1265, B1 => n1902, B2 => n1183
                           , ZN => n1184);
   U425 : INV_X1 port map( A => n1184, ZN => n1185);
   U426 : AOI211_X1 port map( C1 => n1340, C2 => n2461, A => n1186, B => n1185,
                           ZN => n1308);
   U427 : OAI222_X1 port map( A1 => n2465, A2 => n1270, B1 => n2463, B2 => 
                           n1308, C1 => n1187, C2 => n2467, ZN => n1376);
   U428 : INV_X1 port map( A => n1376, ZN => n1271);
   U429 : OAI222_X1 port map( A1 => n1190, A2 => n2467, B1 => n1189, B2 => 
                           n2465, C1 => n1188, C2 => n2463, ZN => n2347);
   U430 : INV_X1 port map( A => n2347, ZN => n1273);
   U431 : INV_X1 port map( A => n2476, ZN => n1957);
   U432 : NAND2_X1 port map( A1 => n1957, A2 => n1191, ZN => n2480);
   U433 : OAI22_X1 port map( A1 => n2283, A2 => n1271, B1 => n1273, B2 => n2480
                           , ZN => n1192);
   U434 : AOI211_X1 port map( C1 => n2476, C2 => n2348, A => n1193, B => n1192,
                           ZN => n1379);
   U435 : INV_X1 port map( A => n1961, ZN => n2487);
   U436 : NOR4_X2 port map( A1 => n1384, A2 => n2729, A3 => DATA2(0), A4 => 
                           n2487, ZN => n2483);
   U437 : INV_X1 port map( A => n2483, ZN => n2118);
   U438 : CLKBUF_X1 port map( A => n1896, Z => n1814);
   U439 : INV_X1 port map( A => DATA1(28), ZN => n2675);
   U440 : NOR2_X1 port map( A1 => n1991, A2 => n2675, ZN => n1680);
   U441 : INV_X1 port map( A => DATA1(30), ZN => n2535_port);
   U442 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(27), ZN => n1580);
   U443 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(26), ZN => n1194);
   U444 : OAI211_X1 port map( C1 => n1678, C2 => n2535_port, A => n1580, B => 
                           n1194, ZN => n1195);
   U445 : AOI211_X1 port map( C1 => DATA1(29), C2 => n2005, A => n1680, B => 
                           n1195, ZN => n2050);
   U446 : OAI222_X1 port map( A1 => n1725, A2 => n1196, B1 => n1723, B2 => 
                           n1204, C1 => n1721, C2 => n2050, ZN => n2124);
   U447 : AOI22_X1 port map( A1 => n2449, A2 => n1205, B1 => n1814, B2 => n2124
                           , ZN => n1199);
   U448 : AOI22_X1 port map( A1 => n2125, A2 => n2120, B1 => n2121, B2 => n1197
                           , ZN => n1198);
   U449 : OAI211_X1 port map( C1 => n1200, C2 => n2446, A => n1199, B => n1198,
                           ZN => n2236);
   U450 : INV_X1 port map( A => n2236, ZN => n1211);
   U451 : INV_X1 port map( A => n1201, ZN => n2237);
   U452 : INV_X1 port map( A => n2124, ZN => n1208);
   U453 : NOR2_X1 port map( A1 => n2428, A2 => n2025, ZN => n1203);
   U454 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(28), ZN => n1593);
   U455 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(29), ZN => n1802);
   U456 : OAI211_X1 port map( C1 => n1660, C2 => n2535_port, A => n1593, B => 
                           n1802, ZN => n1202);
   U457 : AOI211_X1 port map( C1 => DATA1(31), C2 => n2431, A => n1203, B => 
                           n1202, ZN => n2048);
   U458 : OAI222_X1 port map( A1 => n1725, A2 => n1204, B1 => n1723, B2 => 
                           n2050, C1 => n1721, C2 => n2048, ZN => n2123);
   U459 : AOI22_X1 port map( A1 => n2449, A2 => n2120, B1 => n1814, B2 => n2123
                           , ZN => n1207);
   U460 : AOI22_X1 port map( A1 => n2125, A2 => n2122, B1 => n2121, B2 => n1205
                           , ZN => n1206);
   U461 : OAI211_X1 port map( C1 => n1208, C2 => n2446, A => n1207, B => n1206,
                           ZN => n2238);
   U462 : AOI22_X1 port map( A1 => n2342, A2 => n2237, B1 => n1902, B2 => n2238
                           , ZN => n1210);
   U463 : AOI22_X1 port map( A1 => n1641, A2 => n1214, B1 => n2461, B2 => n2239
                           , ZN => n1209);
   U464 : OAI211_X1 port map( C1 => n1211, C2 => n2458, A => n1210, B => n1209,
                           ZN => n2269);
   U465 : OAI22_X1 port map( A1 => n2454, A2 => n1212, B1 => n2456, B2 => n1211
                           , ZN => n1213);
   U466 : INV_X1 port map( A => n1213, ZN => n1216);
   U467 : AOI22_X1 port map( A1 => n2461, A2 => n1214, B1 => n2332, B2 => n2237
                           , ZN => n1215);
   U468 : OAI211_X1 port map( C1 => n1217, C2 => n2452, A => n1216, B => n1215,
                           ZN => n2270);
   U469 : INV_X1 port map( A => n2465, ZN => n2281);
   U470 : INV_X1 port map( A => n1218, ZN => n1221);
   U471 : CLKBUF_X1 port map( A => n1219, Z => n2317);
   U472 : AOI222_X1 port map( A1 => n2269, A2 => n1907, B1 => n2270, B2 => 
                           n2281, C1 => n1221, C2 => n2317, ZN => n2303);
   U473 : INV_X1 port map( A => n2254, ZN => n2473);
   U474 : AOI22_X1 port map( A1 => n2473, A2 => n2347, B1 => n2469, B2 => n2348
                           , ZN => n1223);
   U475 : INV_X1 port map( A => n2480, ZN => n2345);
   U476 : AOI222_X1 port map( A1 => n2270, A2 => n1907, B1 => n1221, B2 => 
                           n2281, C1 => n1220, C2 => n2317, ZN => n1226);
   U477 : INV_X1 port map( A => n1226, ZN => n2346);
   U478 : AOI22_X1 port map( A1 => n2345, A2 => n2346, B1 => n2472, B2 => n1309
                           , ZN => n1222);
   U479 : OAI211_X1 port map( C1 => n1957, C2 => n2303, A => n1223, B => n1222,
                           ZN => n2385);
   U480 : INV_X1 port map( A => n2385, ZN => n2376);
   U481 : NAND3_X1 port map( A1 => n2729, A2 => n1961, A3 => n1276, ZN => n2492
                           );
   U482 : AOI22_X1 port map( A1 => n2469, A2 => n2347, B1 => n2472, B2 => n1342
                           , ZN => n1225);
   U483 : AOI22_X1 port map( A1 => n2473, A2 => n1309, B1 => n2345, B2 => n2348
                           , ZN => n1224);
   U484 : OAI211_X1 port map( C1 => n1957, C2 => n1226, A => n1225, B => n1224,
                           ZN => n2384);
   U485 : INV_X1 port map( A => n2384, ZN => n1296);
   U486 : OAI222_X1 port map( A1 => n2375, A2 => n1379, B1 => n2118, B2 => 
                           n2376, C1 => n2492, C2 => n1296, ZN => n1237);
   U487 : NOR2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n1233);
   U488 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n2391)
                           ;
   U489 : OAI21_X1 port map( B1 => DATA1(9), B2 => DATA2_I_9_port, A => n2391, 
                           ZN => n1851);
   U490 : NOR2_X1 port map( A1 => n1233, A2 => n1851, ZN => n2406);
   U491 : INV_X1 port map( A => DATA1(7), ZN => n2620);
   U492 : XNOR2_X1 port map( A => n2620, B => DATA2_I_7_port, ZN => n1322);
   U493 : INV_X1 port map( A => DATA1(5), ZN => n2553);
   U494 : XOR2_X1 port map( A => n2553, B => DATA2_I_5_port, Z => n1388);
   U495 : INV_X1 port map( A => n1388, ZN => n1390);
   U496 : INV_X1 port map( A => DATA1(3), ZN => n1433);
   U497 : XNOR2_X1 port map( A => n1433, B => DATA2_I_3_port, ZN => n1466);
   U498 : NAND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n1290)
                           ;
   U499 : OAI21_X1 port map( B1 => DATA1(2), B2 => DATA2_I_2_port, A => n1290, 
                           ZN => n1972);
   U500 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n1288)
                           ;
   U501 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n2207)
                           ;
   U502 : INV_X1 port map( A => n2207, ZN => n2414);
   U503 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n2413);
   U504 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n1288, 
                           ZN => n2206);
   U505 : NOR2_X1 port map( A1 => n2413, A2 => n2206, ZN => n2167);
   U506 : OAI21_X1 port map( B1 => cin, B2 => n2414, A => n2167, ZN => n1227);
   U507 : OAI221_X1 port map( B1 => n1972, B2 => n1288, C1 => n1972, C2 => 
                           n1227, A => n1290, ZN => n1228);
   U508 : AND2_X1 port map( A1 => DATA1(3), A2 => DATA2_I_3_port, ZN => n1292);
   U509 : AOI21_X1 port map( B1 => n1466, B2 => n1228, A => n1292, ZN => n1229)
                           ;
   U510 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n1293)
                           ;
   U511 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n1293, 
                           ZN => n1429);
   U512 : OAI21_X1 port map( B1 => n1229, B2 => n1429, A => n1293, ZN => n1230)
                           ;
   U513 : AND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n1294);
   U514 : AOI21_X1 port map( B1 => n1390, B2 => n1230, A => n1294, ZN => n1231)
                           ;
   U515 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n1295)
                           ;
   U516 : OAI21_X1 port map( B1 => DATA1(6), B2 => DATA2_I_6_port, A => n1295, 
                           ZN => n1353);
   U517 : OAI21_X1 port map( B1 => n1231, B2 => n1353, A => n1295, ZN => n1232)
                           ;
   U518 : AOI22_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, B1 => n1322,
                           B2 => n1232, ZN => n1852);
   U519 : NOR2_X1 port map( A1 => n3038, A2 => n1852, ZN => n2405);
   U520 : INV_X1 port map( A => n2405, ZN => n2307);
   U521 : AOI211_X1 port map( C1 => n1233, C2 => n1851, A => n2406, B => n2307,
                           ZN => n1236);
   U522 : NAND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n1257)
                           ;
   U523 : INV_X1 port map( A => DATA1(8), ZN => n2562);
   U524 : INV_X1 port map( A => DATA2_I_8_port, ZN => n1234);
   U525 : NOR3_X1 port map( A1 => n2562, A2 => n1851, A3 => n1234, ZN => n1855)
                           ;
   U526 : NAND2_X1 port map( A1 => n2696, A2 => n1852, ZN => n2388);
   U527 : AOI211_X1 port map( C1 => n1851, C2 => n1257, A => n1855, B => n2388,
                           ZN => n1235);
   U528 : AOI211_X1 port map( C1 => n2688, C2 => n1237, A => n1236, B => n1235,
                           ZN => n1255);
   U529 : OR2_X1 port map( A1 => n2416, A2 => FUNC(3), ZN => n2392);
   U530 : INV_X1 port map( A => n2392, ZN => n2365);
   U531 : NAND2_X1 port map( A1 => FUNC(3), A2 => n1238, ZN => n2412);
   U532 : INV_X1 port map( A => n2412, ZN => n2367);
   U533 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA1(9), B => 
                           DATA2(9), ZN => n1254);
   U534 : NOR2_X1 port map( A1 => n1991, A2 => n2620, ZN => n1362);
   U535 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(8), ZN => n1299);
   U536 : OAI211_X1 port map( C1 => n1678, C2 => n2553, A => n1239, B => n1299,
                           ZN => n1240);
   U537 : AOI211_X1 port map( C1 => DATA1(6), C2 => n2005, A => n1362, B => 
                           n1240, ZN => n1722);
   U538 : NOR2_X1 port map( A1 => n2428, A2 => n2562, ZN => n1258);
   U539 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(6), ZN => n1398);
   U540 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(5), ZN => n1942);
   U541 : OAI211_X1 port map( C1 => n2620, C2 => n1937, A => n1398, B => n1942,
                           ZN => n1241);
   U542 : AOI211_X1 port map( C1 => DATA1(4), C2 => n2431, A => n1258, B => 
                           n1241, ZN => n1720);
   U543 : INV_X1 port map( A => DATA1(6), ZN => n2534_port);
   U544 : NOR2_X1 port map( A1 => n1937, A2 => n2534_port, ZN => n1361);
   U545 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(7), ZN => n1297);
   U546 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(4), ZN => n2174);
   U547 : OAI211_X1 port map( C1 => n1518, C2 => n1433, A => n1297, B => n2174,
                           ZN => n1242);
   U548 : AOI211_X1 port map( C1 => DATA1(5), C2 => n2006, A => n1361, B => 
                           n1242, ZN => n1247);
   U549 : OAI222_X1 port map( A1 => n1725, A2 => n1722, B1 => n1723, B2 => 
                           n1720, C1 => n1721, C2 => n1247, ZN => n1763);
   U550 : INV_X1 port map( A => n1763, ZN => n1901);
   U551 : NOR2_X1 port map( A1 => n1937, A2 => n2553, ZN => n1401);
   U552 : INV_X1 port map( A => DATA1(2), ZN => n2611);
   U553 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(6), ZN => n1331);
   U554 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(3), ZN => n2426);
   U555 : OAI211_X1 port map( C1 => n1518, C2 => n2611, A => n1331, B => n2426,
                           ZN => n1243);
   U556 : AOI211_X1 port map( C1 => DATA1(4), C2 => n2006, A => n1401, B => 
                           n1243, ZN => n1249);
   U557 : OAI222_X1 port map( A1 => n1725, A2 => n1720, B1 => n1723, B2 => 
                           n1247, C1 => n1721, C2 => n1249, ZN => n1898);
   U558 : INV_X1 port map( A => n1898, ZN => n1244);
   U559 : OAI22_X1 port map( A1 => n2440, A2 => n1901, B1 => n1244, B2 => n1687
                           , ZN => n1252);
   U560 : INV_X1 port map( A => DATA1(1), ZN => n2604);
   U561 : INV_X1 port map( A => DATA1(4), ZN => n2613);
   U562 : NOR2_X1 port map( A1 => n1937, A2 => n2613, ZN => n1438);
   U563 : NOR2_X1 port map( A1 => n1991, A2 => n1433, ZN => n2172);
   U564 : AOI211_X1 port map( C1 => DATA1(2), C2 => n1801, A => n1438, B => 
                           n2172, ZN => n1245);
   U565 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(5), ZN => n1363);
   U566 : OAI211_X1 port map( C1 => n1518, C2 => n2604, A => n1245, B => n1363,
                           ZN => n1246);
   U567 : INV_X1 port map( A => n1246, ZN => n1355);
   U568 : OAI222_X1 port map( A1 => n1355, A2 => n1721, B1 => n1247, B2 => 
                           n2049, C1 => n1249, C2 => n2047, ZN => n1897);
   U569 : INV_X1 port map( A => n1897, ZN => n1285);
   U570 : NOR2_X1 port map( A1 => n1937, A2 => n1433, ZN => n1940);
   U571 : INV_X1 port map( A => DATA1(0), ZN => n2603);
   U572 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(4), ZN => n1399);
   U573 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(2), ZN => n2427);
   U574 : OAI211_X1 port map( C1 => n1518, C2 => n2603, A => n1399, B => n2427,
                           ZN => n1248);
   U575 : AOI211_X1 port map( C1 => DATA1(1), C2 => n2005, A => n1940, B => 
                           n1248, ZN => n1394);
   U576 : OAI222_X1 port map( A1 => n1725, A2 => n1249, B1 => n1723, B2 => 
                           n1355, C1 => n1721, C2 => n1394, ZN => n1895);
   U577 : INV_X1 port map( A => n1895, ZN => n1326);
   U578 : OAI22_X1 port map( A1 => n1285, A2 => n2442, B1 => n1326, B2 => n2446
                           , ZN => n1251);
   U579 : NAND2_X1 port map( A1 => n1250, A2 => n2695, ZN => n2382);
   U580 : INV_X1 port map( A => n2382, ZN => n2396);
   U581 : OAI21_X1 port map( B1 => n1252, B2 => n1251, A => n2396, ZN => n1253)
                           ;
   U582 : NAND4_X1 port map( A1 => n1256, A2 => n1255, A3 => n1254, A4 => n1253
                           , ZN => OUTALU(9));
   U583 : OAI21_X1 port map( B1 => DATA1(8), B2 => DATA2_I_8_port, A => n1257, 
                           ZN => n1850);
   U584 : INV_X1 port map( A => n1850, ZN => n1284);
   U585 : OAI22_X1 port map( A1 => n1379, A2 => n2492, B1 => n1296, B2 => n2118
                           , ZN => n1282);
   U586 : AOI21_X1 port map( B1 => DATA1(12), B2 => n2431, A => n1258, ZN => 
                           n1259);
   U587 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(11), ZN => n1569);
   U588 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(10), ZN => n1630);
   U589 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(9), ZN => n1659);
   U590 : NAND4_X1 port map( A1 => n1259, A2 => n1569, A3 => n1630, A4 => n1659
                           , ZN => n1334);
   U591 : AOI222_X1 port map( A1 => n1260, A2 => n2434, B1 => n1334, B2 => 
                           n2176, C1 => n1301, C2 => n2436, ZN => n1405);
   U592 : OAI22_X1 port map( A1 => n2440, A2 => n1405, B1 => n1261, B2 => n2442
                           , ZN => n1263);
   U593 : OAI22_X1 port map( A1 => n1302, A2 => n2446, B1 => n1367, B2 => n2178
                           , ZN => n1262);
   U594 : AOI211_X1 port map( C1 => n1896, C2 => n1264, A => n1263, B => n1262,
                           ZN => n1409);
   U595 : INV_X1 port map( A => n1409, ZN => n1373);
   U596 : AOI22_X1 port map( A1 => n1641, A2 => n1373, B1 => n2342, B2 => n1340
                           , ZN => n1268);
   U597 : AOI22_X1 port map( A1 => n1823, A2 => n1266, B1 => n1902, B2 => n1265
                           , ZN => n1267);
   U598 : OAI211_X1 port map( C1 => n1370, C2 => n1750, A => n1268, B => n1267,
                           ZN => n1269);
   U599 : INV_X1 port map( A => n1269, ZN => n1341);
   U600 : OAI222_X1 port map( A1 => n1270, A2 => n2467, B1 => n1308, B2 => 
                           n2465, C1 => n1341, C2 => n2463, ZN => n1375);
   U601 : INV_X1 port map( A => n1375, ZN => n1415);
   U602 : OAI22_X1 port map( A1 => n2283, A2 => n1415, B1 => n1271, B2 => n2254
                           , ZN => n1275);
   U603 : OAI22_X1 port map( A1 => n1957, A2 => n1273, B1 => n1272, B2 => n2480
                           , ZN => n1274);
   U604 : AOI211_X1 port map( C1 => n2469, C2 => n1342, A => n1275, B => n1274,
                           ZN => n1418);
   U605 : NAND3_X1 port map( A1 => DATA2(1), A2 => n1276, A3 => n1961, ZN => 
                           n2112);
   U606 : OAI22_X1 port map( A1 => n1418, A2 => n2375, B1 => n2376, B2 => n2112
                           , ZN => n1281);
   U607 : AOI222_X1 port map( A1 => n1898, A2 => n2121, B1 => n1897, B2 => 
                           n2449, C1 => n1895, C2 => n2125, ZN => n1279);
   U608 : INV_X1 port map( A => DATA2(8), ZN => n2720);
   U609 : OAI22_X1 port map( A1 => n2562, A2 => DATA2(8), B1 => n2720, B2 => 
                           DATA1(8), ZN => n2557);
   U610 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_8_port, B1 => n2393
                           , B2 => n2557, ZN => n1278);
   U611 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA1(8), B => 
                           DATA2(8), ZN => n1277);
   U612 : OAI211_X1 port map( C1 => n1279, C2 => n2382, A => n1278, B => n1277,
                           ZN => n1280);
   U613 : AOI221_X1 port map( B1 => n1282, B2 => n2688, C1 => n1281, C2 => 
                           n2688, A => n1280, ZN => n1283);
   U614 : OAI221_X1 port map( B1 => n1284, B2 => n2307, C1 => n1850, C2 => 
                           n2388, A => n1283, ZN => OUTALU(8));
   U615 : OAI22_X1 port map( A1 => n2440, A2 => n1285, B1 => n1326, B2 => n2178
                           , ZN => n1287);
   U616 : OAI221_X1 port map( B1 => DATA1(7), B2 => n2416, C1 => n2620, C2 => 
                           n2412, A => n2392, ZN => n1286);
   U617 : AOI22_X1 port map( A1 => n2396, A2 => n1287, B1 => DATA2(7), B2 => 
                           n1286, ZN => n1325);
   U618 : NOR2_X1 port map( A1 => DATA2(7), A2 => n2620, ZN => n2558);
   U619 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_7_port, B1 => n2393
                           , B2 => n2558, ZN => n1324);
   U620 : NOR2_X1 port map( A1 => cin, A2 => n3038, ZN => n2420);
   U621 : INV_X1 port map( A => n2420, ZN => n1938);
   U622 : INV_X1 port map( A => n2206, ZN => n2208);
   U623 : INV_X1 port map( A => n1288, ZN => n1289);
   U624 : AOI21_X1 port map( B1 => n2414, B2 => n2208, A => n1289, ZN => n1971)
                           ;
   U625 : OAI21_X1 port map( B1 => n1971, B2 => n1972, A => n1290, ZN => n1461)
                           ;
   U626 : AOI21_X1 port map( B1 => n1466, B2 => n1461, A => n1292, ZN => n1424)
                           ;
   U627 : OAI21_X1 port map( B1 => n1424, B2 => n1429, A => n1293, ZN => n1359)
                           ;
   U628 : AOI21_X1 port map( B1 => n1390, B2 => n1359, A => n1294, ZN => n1348)
                           ;
   U629 : OAI21_X1 port map( B1 => n1348, B2 => n1353, A => n1295, ZN => n1317)
                           ;
   U630 : NAND2_X1 port map( A1 => n2696, A2 => cin, ZN => n2415);
   U631 : NOR2_X1 port map( A1 => n1289, A2 => n2167, ZN => n1969);
   U632 : OAI21_X1 port map( B1 => n1969, B2 => n1972, A => n1290, ZN => n1465)
                           ;
   U633 : NAND2_X1 port map( A1 => n1466, A2 => n1465, ZN => n1464);
   U634 : INV_X1 port map( A => n1464, ZN => n1291);
   U635 : NOR2_X1 port map( A1 => n1292, A2 => n1291, ZN => n1423);
   U636 : OAI21_X1 port map( B1 => n1423, B2 => n1429, A => n1293, ZN => n1358)
                           ;
   U637 : AOI21_X1 port map( B1 => n1390, B2 => n1358, A => n1294, ZN => n1347)
                           ;
   U638 : OAI21_X1 port map( B1 => n1347, B2 => n1353, A => n1295, ZN => n1316)
                           ;
   U639 : OAI22_X1 port map( A1 => n1938, A2 => n1317, B1 => n2415, B2 => n1316
                           , ZN => n1321);
   U640 : OAI22_X1 port map( A1 => n1418, A2 => n2492, B1 => n1296, B2 => n2112
                           , ZN => n1314);
   U641 : INV_X1 port map( A => n1297, ZN => n1298);
   U642 : AOI21_X1 port map( B1 => DATA1(11), B2 => n2431, A => n1298, ZN => 
                           n1300);
   U643 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(10), ZN => n1610);
   U644 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(9), ZN => n1644);
   U645 : NAND4_X1 port map( A1 => n1300, A2 => n1610, A3 => n1644, A4 => n1299
                           , ZN => n1366);
   U646 : AOI222_X1 port map( A1 => n1301, A2 => n2434, B1 => n1366, B2 => 
                           n2438, C1 => n1334, C2 => n2436, ZN => n1442);
   U647 : OAI22_X1 port map( A1 => n2440, A2 => n1442, B1 => n1367, B2 => n2442
                           , ZN => n1304);
   U648 : OAI22_X1 port map( A1 => n2444, A2 => n1302, B1 => n1405, B2 => n2178
                           , ZN => n1303);
   U649 : AOI211_X1 port map( C1 => n2183, C2 => n1337, A => n1304, B => n1303,
                           ZN => n1445);
   U650 : OAI22_X1 port map( A1 => n1370, A2 => n2452, B1 => n1445, B2 => n2454
                           , ZN => n1307);
   U651 : OAI22_X1 port map( A1 => n2456, A2 => n1305, B1 => n1409, B2 => n1750
                           , ZN => n1306);
   U652 : AOI211_X1 port map( C1 => n1823, C2 => n1340, A => n1307, B => n1306,
                           ZN => n1374);
   U653 : OAI222_X1 port map( A1 => n1308, A2 => n2467, B1 => n1341, B2 => 
                           n2465, C1 => n1374, C2 => n2463, ZN => n1330);
   U654 : AOI22_X1 port map( A1 => n2473, A2 => n1375, B1 => n2472, B2 => n1330
                           , ZN => n1311);
   U655 : AOI22_X1 port map( A1 => n2469, A2 => n1376, B1 => n2476, B2 => n1309
                           , ZN => n1310);
   U656 : OAI211_X1 port map( C1 => n1312, C2 => n2480, A => n1311, B => n1310,
                           ZN => n1455);
   U657 : INV_X1 port map( A => n1455, ZN => n1419);
   U658 : OAI22_X1 port map( A1 => n1419, A2 => n2375, B1 => n1379, B2 => n2118
                           , ZN => n1313);
   U659 : AOI211_X1 port map( C1 => n2487, C2 => n2385, A => n1314, B => n1313,
                           ZN => n1383);
   U660 : NAND2_X1 port map( A1 => DATA2(0), A2 => DATA2(3), ZN => n1315);
   U661 : AOI211_X1 port map( C1 => n2728, C2 => n2729, A => n2727, B => n2726,
                           ZN => n2493);
   U662 : INV_X1 port map( A => n2493, ZN => n1963);
   U663 : NOR3_X1 port map( A1 => n1383, A2 => n2409, A3 => n2079, ZN => n1320)
                           ;
   U664 : INV_X1 port map( A => n2415, ZN => n1970);
   U665 : AOI22_X1 port map( A1 => n2420, A2 => n1317, B1 => n1970, B2 => n1316
                           , ZN => n1318);
   U666 : NOR2_X1 port map( A1 => n1318, A2 => n1322, ZN => n1319);
   U667 : AOI211_X1 port map( C1 => n1322, C2 => n1321, A => n1320, B => n1319,
                           ZN => n1323);
   U668 : NAND3_X1 port map( A1 => n1325, A2 => n1324, A3 => n1323, ZN => 
                           OUTALU(7));
   U669 : AOI22_X1 port map( A1 => n2420, A2 => n1348, B1 => n1970, B2 => n1347
                           , ZN => n1354);
   U670 : NOR3_X1 port map( A1 => n2440, A2 => n1326, A3 => n2382, ZN => n1329)
                           ;
   U671 : INV_X1 port map( A => DATA2(6), ZN => n2724);
   U672 : AOI22_X1 port map( A1 => DATA1(6), A2 => n2724, B1 => DATA2(6), B2 =>
                           n2534_port, ZN => n2617);
   U673 : AOI21_X1 port map( B1 => DATA1(6), B2 => n2367, A => n2365, ZN => 
                           n1327);
   U674 : OAI22_X1 port map( A1 => n2617, A2 => n2416, B1 => n1327, B2 => n2724
                           , ZN => n1328);
   U675 : AOI211_X1 port map( C1 => dataout_mul_6_port, C2 => n2422, A => n1329
                           , B => n1328, ZN => n1352);
   U676 : INV_X1 port map( A => n2079, ZN => n2496);
   U677 : NOR2_X1 port map( A1 => n2493, A2 => n2496, ZN => n2498);
   U678 : INV_X1 port map( A => n2498, ZN => n2066);
   U679 : OAI22_X1 port map( A1 => n1419, A2 => n2492, B1 => n1379, B2 => n2112
                           , ZN => n1346);
   U680 : INV_X1 port map( A => n1330, ZN => n1453);
   U681 : NAND2_X1 port map( A1 => DATA1(10), A2 => n2431, ZN => n1332);
   U682 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(9), ZN => n1629);
   U683 : NAND2_X1 port map( A1 => n2006, A2 => DATA1(8), ZN => n1658);
   U684 : AND4_X1 port map( A1 => n1332, A2 => n1629, A3 => n1658, A4 => n1331,
                           ZN => n1333);
   U685 : OAI21_X1 port map( B1 => n1937, B2 => n2620, A => n1333, ZN => n1403)
                           ;
   U686 : AOI222_X1 port map( A1 => n1334, A2 => n2434, B1 => n1403, B2 => 
                           n2176, C1 => n1366, C2 => n1614, ZN => n1945);
   U687 : OAI22_X1 port map( A1 => n2440, A2 => n1945, B1 => n1405, B2 => n2442
                           , ZN => n1336);
   U688 : OAI22_X1 port map( A1 => n1367, A2 => n2446, B1 => n1442, B2 => n2178
                           , ZN => n1335);
   U689 : AOI211_X1 port map( C1 => n1896, C2 => n1337, A => n1336, B => n1335,
                           ZN => n1949);
   U690 : OAI22_X1 port map( A1 => n1409, A2 => n2452, B1 => n1949, B2 => n2454
                           , ZN => n1339);
   U691 : OAI22_X1 port map( A1 => n1370, A2 => n2458, B1 => n1445, B2 => n1750
                           , ZN => n1338);
   U692 : AOI211_X1 port map( C1 => n1902, C2 => n1340, A => n1339, B => n1338,
                           ZN => n1413);
   U693 : OAI222_X1 port map( A1 => n1341, A2 => n2467, B1 => n1374, B2 => 
                           n2465, C1 => n1413, C2 => n2463, ZN => n1450);
   U694 : AOI22_X1 port map( A1 => n2469, A2 => n1375, B1 => n2472, B2 => n1450
                           , ZN => n1344);
   U695 : AOI22_X1 port map( A1 => n2345, A2 => n1376, B1 => n2476, B2 => n1342
                           , ZN => n1343);
   U696 : OAI211_X1 port map( C1 => n1453, C2 => n2254, A => n1344, B => n1343,
                           ZN => n1454);
   U697 : INV_X1 port map( A => n1454, ZN => n1962);
   U698 : OAI22_X1 port map( A1 => n1418, A2 => n2118, B1 => n1962, B2 => n2375
                           , ZN => n1345);
   U699 : AOI211_X1 port map( C1 => n2487, C2 => n2384, A => n1346, B => n1345,
                           ZN => n1422);
   U700 : OAI22_X1 port map( A1 => n1383, A2 => n2066, B1 => n1422, B2 => n2079
                           , ZN => n1350);
   U701 : OAI22_X1 port map( A1 => n1348, A2 => n1938, B1 => n1347, B2 => n2415
                           , ZN => n1349);
   U702 : AOI22_X1 port map( A1 => n2688, A2 => n1350, B1 => n1353, B2 => n1349
                           , ZN => n1351);
   U703 : OAI211_X1 port map( C1 => n1354, C2 => n1353, A => n1352, B => n1351,
                           ZN => OUTALU(6));
   U704 : OAI21_X1 port map( B1 => n2553, B2 => n2412, A => n2392, ZN => n1357)
                           ;
   U705 : OAI22_X1 port map( A1 => n1355, A2 => n2049, B1 => n1394, B2 => n2047
                           , ZN => n1356);
   U706 : AOI22_X1 port map( A1 => DATA2(5), A2 => n1357, B1 => n2396, B2 => 
                           n1356, ZN => n1393);
   U707 : AOI22_X1 port map( A1 => DATA2(5), A2 => DATA1(5), B1 => n2553, B2 =>
                           n2725, ZN => n2519_port);
   U708 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_5_port, B1 => n2393
                           , B2 => n2519_port, ZN => n1392);
   U709 : OAI22_X1 port map( A1 => n1938, A2 => n1359, B1 => n2415, B2 => n1358
                           , ZN => n1389);
   U710 : AOI22_X1 port map( A1 => n1359, A2 => n2420, B1 => n1358, B2 => n1970
                           , ZN => n1360);
   U711 : INV_X1 port map( A => n1360, ZN => n1387);
   U712 : OAI22_X1 port map( A1 => n1418, A2 => n2112, B1 => n1962, B2 => n2492
                           , ZN => n1382);
   U713 : INV_X1 port map( A => n1945, ZN => n1404);
   U714 : NOR2_X1 port map( A1 => n1362, A2 => n1361, ZN => n1365);
   U715 : NAND2_X1 port map( A1 => DATA1(9), A2 => n2431, ZN => n1364);
   U716 : NAND2_X1 port map( A1 => n2005, A2 => DATA1(8), ZN => n1643);
   U717 : NAND4_X1 port map( A1 => n1365, A2 => n1364, A3 => n1643, A4 => n1363
                           , ZN => n1441);
   U718 : AOI222_X1 port map( A1 => n1366, A2 => n2434, B1 => n1441, B2 => 
                           n2438, C1 => n1403, C2 => n2436, ZN => n2179);
   U719 : OAI22_X1 port map( A1 => n2440, A2 => n2179, B1 => n1442, B2 => n2442
                           , ZN => n1369);
   U720 : OAI22_X1 port map( A1 => n2444, A2 => n1367, B1 => n1405, B2 => n2446
                           , ZN => n1368);
   U721 : AOI211_X1 port map( C1 => n2449, C2 => n1404, A => n1369, B => n1368,
                           ZN => n2184);
   U722 : OAI22_X1 port map( A1 => n1445, A2 => n2452, B1 => n2184, B2 => n2454
                           , ZN => n1372);
   U723 : OAI22_X1 port map( A1 => n2456, A2 => n1370, B1 => n1949, B2 => n1750
                           , ZN => n1371);
   U724 : AOI211_X1 port map( C1 => n1823, C2 => n1373, A => n1372, B => n1371,
                           ZN => n1449);
   U725 : OAI222_X1 port map( A1 => n2465, A2 => n1413, B1 => n2463, B2 => 
                           n1449, C1 => n1374, C2 => n2467, ZN => n2189);
   U726 : AOI22_X1 port map( A1 => n2345, A2 => n1375, B1 => n2472, B2 => n2189
                           , ZN => n1378);
   U727 : AOI22_X1 port map( A1 => n2473, A2 => n1450, B1 => n2476, B2 => n1376
                           , ZN => n1377);
   U728 : OAI211_X1 port map( C1 => n1453, C2 => n2230, A => n1378, B => n1377,
                           ZN => n2192);
   U729 : INV_X1 port map( A => n2192, ZN => n1380);
   U730 : OAI22_X1 port map( A1 => n1380, A2 => n2375, B1 => n1379, B2 => n1961
                           , ZN => n1381);
   U731 : AOI211_X1 port map( C1 => n2483, C2 => n1455, A => n1382, B => n1381,
                           ZN => n1458);
   U732 : OAI222_X1 port map( A1 => n2066, A2 => n1422, B1 => n2079, B2 => 
                           n1458, C1 => n1383, C2 => n1963, ZN => n2199);
   U733 : INV_X1 port map( A => n2199, ZN => n1460);
   U734 : NOR2_X1 port map( A1 => n1384, A2 => n2727, ZN => n1798);
   U735 : AOI21_X1 port map( B1 => DATA2(4), B2 => n1385, A => n1798, ZN => 
                           n2503);
   U736 : INV_X1 port map( A => n2503, ZN => n1917);
   U737 : NOR3_X1 port map( A1 => n1460, A2 => n2409, A3 => n1917, ZN => n1386)
                           ;
   U738 : AOI221_X1 port map( B1 => n1390, B2 => n1389, C1 => n1388, C2 => 
                           n1387, A => n1386, ZN => n1391);
   U739 : NAND3_X1 port map( A1 => n1393, A2 => n1392, A3 => n1391, ZN => 
                           OUTALU(5));
   U740 : AOI22_X1 port map( A1 => n2420, A2 => n1424, B1 => n1970, B2 => n1423
                           , ZN => n1430);
   U741 : NOR3_X1 port map( A1 => n1394, A2 => n2049, A3 => n2382, ZN => n1397)
                           ;
   U742 : AOI22_X1 port map( A1 => DATA2(4), A2 => n2613, B1 => DATA1(4), B2 =>
                           n2726, ZN => n2550);
   U743 : AOI21_X1 port map( B1 => DATA1(4), B2 => n2367, A => n2365, ZN => 
                           n1395);
   U744 : OAI22_X1 port map( A1 => n2550, A2 => n2416, B1 => n1395, B2 => n2726
                           , ZN => n1396);
   U745 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n2422, A => n1397
                           , B => n1396, ZN => n1428);
   U746 : NOR2_X1 port map( A1 => n1798, A2 => n2503, ZN => n2198);
   U747 : INV_X1 port map( A => n2198, ZN => n2510);
   U748 : INV_X1 port map( A => n2492, ZN => n2386);
   U749 : INV_X1 port map( A => n2184, ZN => n1412);
   U750 : OAI211_X1 port map( C1 => n1518, C2 => n2562, A => n1399, B => n1398,
                           ZN => n1400);
   U751 : AOI211_X1 port map( C1 => DATA1(7), C2 => n2005, A => n1401, B => 
                           n1400, ZN => n1402);
   U752 : INV_X1 port map( A => n1402, ZN => n1944);
   U753 : AOI222_X1 port map( A1 => n2176, A2 => n1944, B1 => n2436, B2 => 
                           n1441, C1 => n2434, C2 => n1403, ZN => n2443);
   U754 : INV_X1 port map( A => n2443, ZN => n2182);
   U755 : AOI22_X1 port map( A1 => n2125, A2 => n1404, B1 => n1745, B2 => n2182
                           , ZN => n1408);
   U756 : OAI22_X1 port map( A1 => n2178, A2 => n2179, B1 => n2444, B2 => n1405
                           , ZN => n1406);
   U757 : INV_X1 port map( A => n1406, ZN => n1407);
   U758 : OAI211_X1 port map( C1 => n1442, C2 => n2446, A => n1408, B => n1407,
                           ZN => n1448);
   U759 : INV_X1 port map( A => n1448, ZN => n2455);
   U760 : OAI22_X1 port map( A1 => n2454, A2 => n2455, B1 => n2452, B2 => n1949
                           , ZN => n1411);
   U761 : OAI22_X1 port map( A1 => n2458, A2 => n1445, B1 => n2456, B2 => n1409
                           , ZN => n1410);
   U762 : AOI211_X1 port map( C1 => n1412, C2 => n2461, A => n1411, B => n1410,
                           ZN => n1953);
   U763 : OAI222_X1 port map( A1 => n1413, A2 => n2467, B1 => n1449, B2 => 
                           n2465, C1 => n1953, C2 => n2463, ZN => n2475);
   U764 : INV_X1 port map( A => n2475, ZN => n1414);
   U765 : INV_X1 port map( A => n1450, ZN => n1956);
   U766 : OAI22_X1 port map( A1 => n2283, A2 => n1414, B1 => n1956, B2 => n2230
                           , ZN => n1417);
   U767 : OAI22_X1 port map( A1 => n1957, A2 => n1415, B1 => n1453, B2 => n2480
                           , ZN => n1416);
   U768 : AOI211_X1 port map( C1 => n2473, C2 => n2189, A => n1417, B => n1416,
                           ZN => n1958);
   U769 : OAI22_X1 port map( A1 => n1962, A2 => n2118, B1 => n1958, B2 => n2375
                           , ZN => n1421);
   U770 : OAI22_X1 port map( A1 => n1419, A2 => n2112, B1 => n1418, B2 => n1961
                           , ZN => n1420);
   U771 : AOI211_X1 port map( C1 => n2386, C2 => n2192, A => n1421, B => n1420,
                           ZN => n1964);
   U772 : OAI222_X1 port map( A1 => n2066, A2 => n1458, B1 => n2079, B2 => 
                           n1964, C1 => n1422, C2 => n1963, ZN => n2506);
   U773 : INV_X1 port map( A => n2506, ZN => n1459);
   U774 : OAI22_X1 port map( A1 => n1460, A2 => n2510, B1 => n1459, B2 => n1917
                           , ZN => n1426);
   U775 : OAI22_X1 port map( A1 => n1424, A2 => n1938, B1 => n1423, B2 => n2415
                           , ZN => n1425);
   U776 : AOI22_X1 port map( A1 => n2688, A2 => n1426, B1 => n1429, B2 => n1425
                           , ZN => n1427);
   U777 : OAI211_X1 port map( C1 => n1430, C2 => n1429, A => n1428, B => n1427,
                           ZN => OUTALU(4));
   U778 : NOR2_X1 port map( A1 => n2428, A2 => n1433, ZN => n1437);
   U779 : NOR2_X1 port map( A1 => n1937, A2 => n2611, ZN => n2173);
   U780 : AOI211_X1 port map( C1 => DATA1(0), C2 => n2005, A => n1437, B => 
                           n2173, ZN => n1431);
   U781 : OAI21_X1 port map( B1 => n1991, B2 => n2604, A => n1431, ZN => n1432)
                           ;
   U782 : AOI22_X1 port map( A1 => DATA2(3), A2 => DATA1(3), B1 => n1433, B2 =>
                           n2727, ZN => n2525_port);
   U783 : AOI22_X1 port map( A1 => n2396, A2 => n1432, B1 => n2393, B2 => 
                           n2525_port, ZN => n1470);
   U784 : OAI21_X1 port map( B1 => n1433, B2 => n2412, A => n2392, ZN => n1435)
                           ;
   U785 : CLKBUF_X1 port map( A => n1434, Z => n2314);
   U786 : AOI22_X1 port map( A1 => DATA2(3), A2 => n1435, B1 => n2314, B2 => 
                           dataout_mul_3_port, ZN => n1469);
   U787 : NAND2_X1 port map( A1 => n1798, A2 => n1436, ZN => n2202);
   U788 : AOI211_X1 port map( C1 => DATA1(6), C2 => n1801, A => n1438, B => 
                           n1437, ZN => n1440);
   U789 : NAND2_X1 port map( A1 => DATA1(7), A2 => n2431, ZN => n1439);
   U790 : OAI211_X1 port map( C1 => n1991, C2 => n2553, A => n1440, B => n1439,
                           ZN => n2177);
   U791 : AOI222_X1 port map( A1 => n1441, A2 => n2434, B1 => n2177, B2 => 
                           n2438, C1 => n1944, C2 => n1614, ZN => n2445);
   U792 : OAI22_X1 port map( A1 => n2440, A2 => n2445, B1 => n2179, B2 => n2442
                           , ZN => n1444);
   U793 : OAI22_X1 port map( A1 => n2444, A2 => n1442, B1 => n1945, B2 => n2446
                           , ZN => n1443);
   U794 : AOI211_X1 port map( C1 => n2449, C2 => n2182, A => n1444, B => n1443,
                           ZN => n2457);
   U795 : OAI22_X1 port map( A1 => n2184, A2 => n2452, B1 => n2457, B2 => n2454
                           , ZN => n1447);
   U796 : OAI22_X1 port map( A1 => n2456, A2 => n1445, B1 => n1949, B2 => n2458
                           , ZN => n1446);
   U797 : AOI211_X1 port map( C1 => n2461, C2 => n1448, A => n1447, B => n1446,
                           ZN => n2188);
   U798 : OAI222_X1 port map( A1 => n2465, A2 => n1953, B1 => n2463, B2 => 
                           n2188, C1 => n1449, C2 => n2467, ZN => n2171);
   U799 : AOI22_X1 port map( A1 => n2473, A2 => n2475, B1 => n2472, B2 => n2171
                           , ZN => n1452);
   U800 : AOI22_X1 port map( A1 => n2469, A2 => n2189, B1 => n2345, B2 => n1450
                           , ZN => n1451);
   U801 : OAI211_X1 port map( C1 => n1957, C2 => n1453, A => n1452, B => n1451,
                           ZN => n2486);
   U802 : AOI22_X1 port map( A1 => n2481, A2 => n2486, B1 => n2483, B2 => n2192
                           , ZN => n1457);
   U803 : INV_X1 port map( A => n2112, ZN => n2485);
   U804 : AOI22_X1 port map( A1 => n2487, A2 => n1455, B1 => n2485, B2 => n1454
                           , ZN => n1456);
   U805 : OAI211_X1 port map( C1 => n1958, C2 => n2492, A => n1457, B => n1456,
                           ZN => n2196);
   U806 : INV_X1 port map( A => n2196, ZN => n1966);
   U807 : OAI222_X1 port map( A1 => n2066, A2 => n1964, B1 => n2079, B2 => 
                           n1966, C1 => n1458, C2 => n1963, ZN => n2504);
   U808 : INV_X1 port map( A => n2504, ZN => n2203);
   U809 : OAI222_X1 port map( A1 => n2202, A2 => n1460, B1 => n2510, B2 => 
                           n1459, C1 => n1917, C2 => n2203, ZN => n1463);
   U810 : XOR2_X1 port map( A => n1466, B => n1461, Z => n1462);
   U811 : AOI22_X1 port map( A1 => n2688, A2 => n1463, B1 => n2420, B2 => n1462
                           , ZN => n1468);
   U812 : OAI211_X1 port map( C1 => n1466, C2 => n1465, A => n1970, B => n1464,
                           ZN => n1467);
   U813 : NAND4_X1 port map( A1 => n1470, A2 => n1469, A3 => n1468, A4 => n1467
                           , ZN => OUTALU(3));
   U814 : OAI211_X1 port map( C1 => n1678, C2 => n2532_port, A => n1472, B => 
                           n1471, ZN => n1473);
   U815 : AOI211_X1 port map( C1 => DATA1(18), C2 => n2170, A => n1474, B => 
                           n1473, ZN => n1475);
   U816 : INV_X1 port map( A => n1475, ZN => n1505);
   U817 : OAI211_X1 port map( C1 => n1678, C2 => n2602, A => n1477, B => n1476,
                           ZN => n1478);
   U818 : AOI211_X1 port map( C1 => DATA1(17), C2 => n2170, A => n1479, B => 
                           n1478, ZN => n1480);
   U819 : INV_X1 port map( A => n1480, ZN => n1494);
   U820 : INV_X1 port map( A => DATA1(12), ZN => n2633);
   U821 : OAI211_X1 port map( C1 => n1518, C2 => n2633, A => n1482, B => n1481,
                           ZN => n1483);
   U822 : AOI211_X1 port map( C1 => DATA1(16), C2 => n2170, A => n1484, B => 
                           n1483, ZN => n1485);
   U823 : INV_X1 port map( A => n1485, ZN => n1573);
   U824 : AOI222_X1 port map( A1 => n2176, A2 => n1505, B1 => n2436, B2 => 
                           n1494, C1 => n2434, C2 => n1573, ZN => n1616);
   U825 : INV_X1 port map( A => n1616, ZN => n1636);
   U826 : AOI22_X1 port map( A1 => DATA1(14), A2 => n2205, B1 => DATA1(11), B2 
                           => n2431, ZN => n1489);
   U827 : NAND4_X1 port map( A1 => n1489, A2 => n1488, A3 => n1487, A4 => n1486
                           , ZN => n1615);
   U828 : AOI222_X1 port map( A1 => n1615, A2 => n2434, B1 => n1494, B2 => 
                           n2438, C1 => n1573, C2 => n2436, ZN => n1648);
   U829 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1801, B1 => DATA1(15), B2 
                           => n2431, ZN => n1493);
   U830 : NAND4_X1 port map( A1 => n1493, A2 => n1492, A3 => n1491, A4 => n1490
                           , ZN => n1504);
   U831 : AOI222_X1 port map( A1 => n1494, A2 => n2434, B1 => n1504, B2 => 
                           n2438, C1 => n1505, C2 => n2436, ZN => n1574);
   U832 : OAI22_X1 port map( A1 => n2444, A2 => n1648, B1 => n1574, B2 => n2442
                           , ZN => n1507);
   U833 : AOI22_X1 port map( A1 => DATA1(18), A2 => n1801, B1 => DATA1(17), B2 
                           => n2431, ZN => n1499);
   U834 : INV_X1 port map( A => n1495, ZN => n1496);
   U835 : NAND4_X1 port map( A1 => n1499, A2 => n1498, A3 => n1497, A4 => n1496
                           , ZN => n1530);
   U836 : AOI22_X1 port map( A1 => n1801, A2 => DATA1(17), B1 => DATA1(16), B2 
                           => n2431, ZN => n1503);
   U837 : NAND4_X1 port map( A1 => n1503, A2 => n1502, A3 => n1501, A4 => n1500
                           , ZN => n1528);
   U838 : AOI222_X1 port map( A1 => n1504, A2 => n2434, B1 => n1530, B2 => 
                           n2438, C1 => n1528, C2 => n2436, ZN => n1543);
   U839 : AOI222_X1 port map( A1 => n1505, A2 => n2434, B1 => n1528, B2 => 
                           n2438, C1 => n1504, C2 => n2436, ZN => n1568);
   U840 : OAI22_X1 port map( A1 => n1543, A2 => n2440, B1 => n1568, B2 => n2178
                           , ZN => n1506);
   U841 : AOI211_X1 port map( C1 => n2183, C2 => n1636, A => n1507, B => n1506,
                           ZN => n1651);
   U842 : AOI22_X1 port map( A1 => n1801, A2 => DATA1(20), B1 => DATA1(19), B2 
                           => n2431, ZN => n1511);
   U843 : NAND4_X1 port map( A1 => n1511, A2 => n1510, A3 => n1509, A4 => n1508
                           , ZN => n1521);
   U844 : AOI22_X1 port map( A1 => n1801, A2 => DATA1(19), B1 => DATA1(18), B2 
                           => n2431, ZN => n1515);
   U845 : NAND4_X1 port map( A1 => n1515, A2 => n1514, A3 => n1513, A4 => n1512
                           , ZN => n1529);
   U846 : AOI222_X1 port map( A1 => n1530, A2 => n2434, B1 => n1521, B2 => 
                           n2438, C1 => n1529, C2 => n2436, ZN => n1533);
   U847 : OAI211_X1 port map( C1 => n1518, C2 => n2653, A => n1517, B => n1516,
                           ZN => n1519);
   U848 : AOI211_X1 port map( C1 => n2170, C2 => DATA1(24), A => n1520, B => 
                           n1519, ZN => n1550);
   U849 : INV_X1 port map( A => n1521, ZN => n1527);
   U850 : INV_X1 port map( A => n1529, ZN => n1522);
   U851 : OAI222_X1 port map( A1 => n1725, A2 => n1550, B1 => n1723, B2 => 
                           n1527, C1 => n1721, C2 => n1522, ZN => n1585);
   U852 : OAI211_X1 port map( C1 => n1678, C2 => n2652, A => n1524, B => n1523,
                           ZN => n1525);
   U853 : AOI211_X1 port map( C1 => n2170, C2 => DATA1(25), A => n1526, B => 
                           n1525, ZN => n1560);
   U854 : OAI222_X1 port map( A1 => n1725, A2 => n1560, B1 => n1723, B2 => 
                           n1550, C1 => n1721, C2 => n1527, ZN => n1561);
   U855 : AOI22_X1 port map( A1 => n2449, A2 => n1585, B1 => n1745, B2 => n1561
                           , ZN => n1532);
   U856 : AOI222_X1 port map( A1 => n2436, A2 => n1530, B1 => n2176, B2 => 
                           n1529, C1 => n2434, C2 => n1528, ZN => n1539);
   U857 : INV_X1 port map( A => n1539, ZN => n1551);
   U858 : INV_X1 port map( A => n1543, ZN => n1536);
   U859 : AOI22_X1 port map( A1 => n1761, A2 => n1551, B1 => n1814, B2 => n1536
                           , ZN => n1531);
   U860 : OAI211_X1 port map( C1 => n1533, C2 => n2442, A => n1532, B => n1531,
                           ZN => n1588);
   U861 : INV_X1 port map( A => n1533, ZN => n1562);
   U862 : INV_X1 port map( A => n1574, ZN => n1619);
   U863 : AOI22_X1 port map( A1 => n1562, A2 => n2121, B1 => n1814, B2 => n1619
                           , ZN => n1535);
   U864 : INV_X1 port map( A => n1568, ZN => n1540);
   U865 : AOI22_X1 port map( A1 => n1761, A2 => n1540, B1 => n2449, B2 => n1551
                           , ZN => n1534);
   U866 : OAI211_X1 port map( C1 => n1543, C2 => n2442, A => n1535, B => n1534,
                           ZN => n1620);
   U867 : AOI22_X1 port map( A1 => n1641, A2 => n1588, B1 => n2342, B2 => n1620
                           , ZN => n1545);
   U868 : AOI22_X1 port map( A1 => n2449, A2 => n1562, B1 => n1745, B2 => n1585
                           , ZN => n1538);
   U869 : AOI22_X1 port map( A1 => n1761, A2 => n1536, B1 => n1814, B2 => n1540
                           , ZN => n1537);
   U870 : OAI211_X1 port map( C1 => n1539, C2 => n2442, A => n1538, B => n1537,
                           ZN => n1589);
   U871 : AOI22_X1 port map( A1 => n2125, A2 => n1540, B1 => n1551, B2 => n1745
                           , ZN => n1542);
   U872 : AOI22_X1 port map( A1 => n1761, A2 => n1619, B1 => n1814, B2 => n1636
                           , ZN => n1541);
   U873 : OAI211_X1 port map( C1 => n1543, C2 => n1687, A => n1542, B => n1541,
                           ZN => n1640);
   U874 : AOI22_X1 port map( A1 => n2461, A2 => n1589, B1 => n2332, B2 => n1640
                           , ZN => n1544);
   U875 : OAI211_X1 port map( C1 => n2456, C2 => n1651, A => n1545, B => n1544,
                           ZN => n1625);
   U876 : INV_X1 port map( A => n1588, ZN => n1604);
   U877 : INV_X1 port map( A => n1561, ZN => n1599);
   U878 : OAI211_X1 port map( C1 => n1678, C2 => n2126, A => n1547, B => n1546,
                           ZN => n1548);
   U879 : AOI211_X1 port map( C1 => n2170, C2 => DATA1(26), A => n1549, B => 
                           n1548, ZN => n1584);
   U880 : OAI222_X1 port map( A1 => n1725, A2 => n1584, B1 => n2047, B2 => 
                           n1560, C1 => n1721, C2 => n1550, ZN => n1684);
   U881 : AOI22_X1 port map( A1 => n1761, A2 => n1562, B1 => n2121, B2 => n1684
                           , ZN => n1553);
   U882 : AOI22_X1 port map( A1 => n2125, A2 => n1585, B1 => n1814, B2 => n1551
                           , ZN => n1552);
   U883 : OAI211_X1 port map( C1 => n1599, C2 => n2178, A => n1553, B => n1552,
                           ZN => n1688);
   U884 : AOI22_X1 port map( A1 => n1641, A2 => n1688, B1 => n2332, B2 => n1620
                           , ZN => n1555);
   U885 : AOI22_X1 port map( A1 => n2342, A2 => n1589, B1 => n1902, B2 => n1640
                           , ZN => n1554);
   U886 : OAI211_X1 port map( C1 => n1604, C2 => n1750, A => n1555, B => n1554,
                           ZN => n1608);
   U887 : INV_X1 port map( A => n1688, ZN => n1603);
   U888 : INV_X1 port map( A => n1684, ZN => n1565);
   U889 : OAI211_X1 port map( C1 => n1678, C2 => n2093, A => n1557, B => n1556,
                           ZN => n1558);
   U890 : AOI211_X1 port map( C1 => n2170, C2 => DATA1(27), A => n1559, B => 
                           n1558, ZN => n1592);
   U891 : OAI222_X1 port map( A1 => n1725, A2 => n1592, B1 => n1723, B2 => 
                           n1584, C1 => n1721, C2 => n1560, ZN => n1813);
   U892 : AOI22_X1 port map( A1 => n2125, A2 => n1561, B1 => n2121, B2 => n1813
                           , ZN => n1564);
   U893 : AOI22_X1 port map( A1 => n1761, A2 => n1585, B1 => n1562, B2 => n1896
                           , ZN => n1563);
   U894 : OAI211_X1 port map( C1 => n1565, C2 => n1687, A => n1564, B => n1563,
                           ZN => n1818);
   U895 : AOI22_X1 port map( A1 => n1641, A2 => n1818, B1 => n2342, B2 => n1588
                           , ZN => n1567);
   U896 : AOI22_X1 port map( A1 => n1823, A2 => n1589, B1 => n1902, B2 => n1620
                           , ZN => n1566);
   U897 : OAI211_X1 port map( C1 => n1603, C2 => n1750, A => n1567, B => n1566,
                           ZN => n1609);
   U898 : AOI222_X1 port map( A1 => n1625, A2 => n1907, B1 => n1608, B2 => 
                           n2281, C1 => n1609, C2 => n2317, ZN => n1829);
   U899 : INV_X1 port map( A => n1589, ZN => n1579);
   U900 : INV_X1 port map( A => n1651, ZN => n1621);
   U901 : AOI22_X1 port map( A1 => n1620, A2 => n2461, B1 => n1621, B2 => n1823
                           , ZN => n1578);
   U902 : OAI22_X1 port map( A1 => n2440, A2 => n1568, B1 => n1648, B2 => n2446
                           , ZN => n1576);
   U903 : AOI22_X1 port map( A1 => DATA1(14), A2 => n2170, B1 => DATA1(10), B2 
                           => n2431, ZN => n1572);
   U904 : NAND4_X1 port map( A1 => n1572, A2 => n1571, A3 => n1570, A4 => n1569
                           , ZN => n1633);
   U905 : AOI222_X1 port map( A1 => n1633, A2 => n2434, B1 => n1573, B2 => 
                           n2438, C1 => n1615, C2 => n1614, ZN => n1667);
   U906 : OAI22_X1 port map( A1 => n2444, A2 => n1667, B1 => n1574, B2 => n2178
                           , ZN => n1575);
   U907 : AOI211_X1 port map( C1 => n2125, C2 => n1636, A => n1576, B => n1575,
                           ZN => n1637);
   U908 : INV_X1 port map( A => n1637, ZN => n1669);
   U909 : AOI22_X1 port map( A1 => n1902, A2 => n1669, B1 => n1640, B2 => n2342
                           , ZN => n1577);
   U910 : OAI211_X1 port map( C1 => n2454, C2 => n1579, A => n1578, B => n1577,
                           ZN => n1672);
   U911 : AOI222_X1 port map( A1 => n2281, A2 => n1625, B1 => n2317, B2 => 
                           n1608, C1 => n1672, C2 => n1907, ZN => n1695);
   U912 : INV_X1 port map( A => n1695, ZN => n1701);
   U913 : INV_X1 port map( A => n1818, ZN => n1602);
   U914 : AOI22_X1 port map( A1 => DATA1(25), A2 => n1801, B1 => DATA1(24), B2 
                           => n2431, ZN => n1582);
   U915 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(28), ZN => n2008);
   U916 : NAND4_X1 port map( A1 => n1582, A2 => n1581, A3 => n1580, A4 => n2008
                           , ZN => n1682);
   U917 : INV_X1 port map( A => n1682, ZN => n1583);
   U918 : OAI222_X1 port map( A1 => n1584, A2 => n1721, B1 => n1583, B2 => 
                           n2049, C1 => n1592, C2 => n2047, ZN => n1598);
   U919 : AOI22_X1 port map( A1 => n2121, A2 => n1598, B1 => n1684, B2 => n2125
                           , ZN => n1587);
   U920 : AOI22_X1 port map( A1 => n1896, A2 => n1585, B1 => n1813, B2 => n2449
                           , ZN => n1586);
   U921 : OAI211_X1 port map( C1 => n2446, C2 => n1599, A => n1587, B => n1586,
                           ZN => n1822);
   U922 : AOI22_X1 port map( A1 => n1688, A2 => n2342, B1 => n1822, B2 => n1641
                           , ZN => n1591);
   U923 : AOI22_X1 port map( A1 => n1902, A2 => n1589, B1 => n1588, B2 => n1823
                           , ZN => n1590);
   U924 : OAI211_X1 port map( C1 => n1750, C2 => n1602, A => n1591, B => n1590,
                           ZN => n1692);
   U925 : INV_X1 port map( A => n1592, ZN => n1596);
   U926 : AOI22_X1 port map( A1 => DATA1(26), A2 => n1801, B1 => DATA1(25), B2 
                           => n2431, ZN => n1595);
   U927 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(29), ZN => n1989);
   U928 : NAND4_X1 port map( A1 => n1595, A2 => n1594, A3 => n1593, A4 => n1989
                           , ZN => n1806);
   U929 : AOI222_X1 port map( A1 => n1596, A2 => n2434, B1 => n1806, B2 => 
                           n2438, C1 => n1682, C2 => n2436, ZN => n1807);
   U930 : INV_X1 port map( A => n1813, ZN => n1597);
   U931 : OAI22_X1 port map( A1 => n2440, A2 => n1807, B1 => n1597, B2 => n2442
                           , ZN => n1601);
   U932 : INV_X1 port map( A => n1598, ZN => n1810);
   U933 : OAI22_X1 port map( A1 => n2444, A2 => n1599, B1 => n1810, B2 => n2178
                           , ZN => n1600);
   U934 : AOI211_X1 port map( C1 => n2183, C2 => n1684, A => n1601, B => n1600,
                           ZN => n1816);
   U935 : OAI22_X1 port map( A1 => n1602, A2 => n2452, B1 => n1816, B2 => n2454
                           , ZN => n1606);
   U936 : OAI22_X1 port map( A1 => n1604, A2 => n2456, B1 => n1603, B2 => n2458
                           , ZN => n1605);
   U937 : AOI211_X1 port map( C1 => n2461, C2 => n1822, A => n1606, B => n1605,
                           ZN => n1824);
   U938 : INV_X1 port map( A => n1824, ZN => n1691);
   U939 : AOI222_X1 port map( A1 => n2281, A2 => n1692, B1 => n2317, B2 => 
                           n1691, C1 => n1609, C2 => n1907, ZN => n1607);
   U940 : INV_X1 port map( A => n1607, ZN => n1828);
   U941 : AOI22_X1 port map( A1 => n2345, A2 => n1701, B1 => n2472, B2 => n1828
                           , ZN => n1628);
   U942 : AOI222_X1 port map( A1 => n2281, A2 => n1609, B1 => n2317, B2 => 
                           n1692, C1 => n1608, C2 => n1907, ZN => n1830);
   U943 : INV_X1 port map( A => n1640, ZN => n1624);
   U944 : AOI22_X1 port map( A1 => DATA1(13), A2 => n2170, B1 => DATA1(9), B2 
                           => n2431, ZN => n1613);
   U945 : NAND4_X1 port map( A1 => n1613, A2 => n1612, A3 => n1611, A4 => n1610
                           , ZN => n1647);
   U946 : AOI222_X1 port map( A1 => n1647, A2 => n2434, B1 => n1615, B2 => 
                           n2438, C1 => n1633, C2 => n1614, ZN => n1708);
   U947 : OAI22_X1 port map( A1 => n2444, A2 => n1708, B1 => n1648, B2 => n2442
                           , ZN => n1618);
   U948 : OAI22_X1 port map( A1 => n1616, A2 => n1687, B1 => n1667, B2 => n2446
                           , ZN => n1617);
   U949 : AOI211_X1 port map( C1 => n2121, C2 => n1619, A => n1618, B => n1617,
                           ZN => n1710);
   U950 : INV_X1 port map( A => n1710, ZN => n1668);
   U951 : AOI22_X1 port map( A1 => n1902, A2 => n1668, B1 => n1620, B2 => n1641
                           , ZN => n1623);
   U952 : AOI22_X1 port map( A1 => n1621, A2 => n2342, B1 => n1669, B2 => n1823
                           , ZN => n1622);
   U953 : OAI211_X1 port map( C1 => n1750, C2 => n1624, A => n1623, B => n1622,
                           ZN => n1673);
   U954 : AOI222_X1 port map( A1 => n2281, A2 => n1672, B1 => n2317, B2 => 
                           n1625, C1 => n1673, C2 => n1907, ZN => n1715);
   U955 : OAI22_X1 port map( A1 => n2254, A2 => n1830, B1 => n1957, B2 => n1715
                           , ZN => n1626);
   U956 : INV_X1 port map( A => n1626, ZN => n1627);
   U957 : OAI211_X1 port map( C1 => n1829, C2 => n2230, A => n1628, B => n1627,
                           ZN => n1835);
   U958 : OAI22_X1 port map( A1 => n1651, A2 => n1750, B1 => n1710, B2 => n2458
                           , ZN => n1639);
   U959 : AOI22_X1 port map( A1 => DATA1(12), A2 => n2170, B1 => DATA1(8), B2 
                           => n2431, ZN => n1632);
   U960 : NAND4_X1 port map( A1 => n1632, A2 => n1631, A3 => n1630, A4 => n1629
                           , ZN => n1656);
   U961 : AOI222_X1 port map( A1 => n1656, A2 => n2434, B1 => n1633, B2 => 
                           n2438, C1 => n1647, C2 => n2436, ZN => n1728);
   U962 : OAI22_X1 port map( A1 => n2444, A2 => n1728, B1 => n1667, B2 => n2442
                           , ZN => n1635);
   U963 : OAI22_X1 port map( A1 => n1648, A2 => n1687, B1 => n1708, B2 => n2446
                           , ZN => n1634);
   U964 : AOI211_X1 port map( C1 => n2121, C2 => n1636, A => n1635, B => n1634,
                           ZN => n1731);
   U965 : OAI22_X1 port map( A1 => n2456, A2 => n1731, B1 => n1637, B2 => n2452
                           , ZN => n1638);
   U966 : AOI211_X1 port map( C1 => n1641, C2 => n1640, A => n1639, B => n1638,
                           ZN => n1642);
   U967 : INV_X1 port map( A => n1642, ZN => n1674);
   U968 : INV_X1 port map( A => n1728, ZN => n1705);
   U969 : AOI22_X1 port map( A1 => DATA1(11), A2 => n2170, B1 => DATA1(7), B2 
                           => n2431, ZN => n1646);
   U970 : NAND4_X1 port map( A1 => n1646, A2 => n1645, A3 => n1644, A4 => n1643
                           , ZN => n1657);
   U971 : AOI222_X1 port map( A1 => n1657, A2 => n2434, B1 => n1647, B2 => 
                           n2176, C1 => n1656, C2 => n2436, ZN => n1655);
   U972 : OAI22_X1 port map( A1 => n2444, A2 => n1655, B1 => n1708, B2 => n2442
                           , ZN => n1650);
   U973 : OAI22_X1 port map( A1 => n2440, A2 => n1648, B1 => n1667, B2 => n1687
                           , ZN => n1649);
   U974 : AOI211_X1 port map( C1 => n2183, C2 => n1705, A => n1650, B => n1649,
                           ZN => n1709);
   U975 : OAI22_X1 port map( A1 => n2456, A2 => n1709, B1 => n1651, B2 => n2454
                           , ZN => n1653);
   U976 : OAI22_X1 port map( A1 => n1710, A2 => n2452, B1 => n1731, B2 => n2458
                           , ZN => n1652);
   U977 : AOI211_X1 port map( C1 => n2461, C2 => n1669, A => n1653, B => n1652,
                           ZN => n1654);
   U978 : INV_X1 port map( A => n1654, ZN => n1714);
   U979 : AOI222_X1 port map( A1 => n2281, A2 => n1674, B1 => n2317, B2 => 
                           n1673, C1 => n1714, C2 => n1907, ZN => n1733);
   U980 : INV_X1 port map( A => n1733, ZN => n1780);
   U981 : INV_X1 port map( A => n1655, ZN => n1744);
   U982 : AOI22_X1 port map( A1 => n2125, A2 => n1705, B1 => n1761, B2 => n1744
                           , ZN => n1666);
   U983 : INV_X1 port map( A => n1708, ZN => n1664);
   U984 : INV_X1 port map( A => n1656, ZN => n1663);
   U985 : INV_X1 port map( A => n1657, ZN => n1704);
   U986 : OAI211_X1 port map( C1 => n2620, C2 => n1660, A => n1659, B => n1658,
                           ZN => n1661);
   U987 : AOI211_X1 port map( C1 => DATA1(6), C2 => n2431, A => n1662, B => 
                           n1661, ZN => n1724);
   U988 : OAI222_X1 port map( A1 => n1725, A2 => n1663, B1 => n1723, B2 => 
                           n1704, C1 => n1721, C2 => n1724, ZN => n1743);
   U989 : AOI22_X1 port map( A1 => n2449, A2 => n1664, B1 => n1814, B2 => n1743
                           , ZN => n1665);
   U990 : OAI211_X1 port map( C1 => n2440, C2 => n1667, A => n1666, B => n1665,
                           ZN => n1752);
   U991 : AOI22_X1 port map( A1 => n2461, A2 => n1668, B1 => n1902, B2 => n1752
                           , ZN => n1671);
   U992 : INV_X1 port map( A => n1709, ZN => n1753);
   U993 : AOI22_X1 port map( A1 => n2397, A2 => n1669, B1 => n1823, B2 => n1753
                           , ZN => n1670);
   U994 : OAI211_X1 port map( C1 => n1731, C2 => n2452, A => n1671, B => n1670,
                           ZN => n1732);
   U995 : AOI222_X1 port map( A1 => n1732, A2 => n1907, B1 => n1714, B2 => 
                           n2281, C1 => n1674, C2 => n2317, ZN => n1777);
   U996 : AOI222_X1 port map( A1 => n1674, A2 => n1907, B1 => n1673, B2 => 
                           n2281, C1 => n1672, C2 => n2317, ZN => n1734);
   U997 : OAI22_X1 port map( A1 => n1957, A2 => n1777, B1 => n1734, B2 => n2230
                           , ZN => n1676);
   U998 : OAI22_X1 port map( A1 => n2283, A2 => n1695, B1 => n1715, B2 => n2254
                           , ZN => n1675);
   U999 : AOI211_X1 port map( C1 => n2345, C2 => n1780, A => n1676, B => n1675,
                           ZN => n1790);
   U1000 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(29), ZN => n2007);
   U1001 : OAI211_X1 port map( C1 => n1678, C2 => n2512, A => n1677, B => n2007
                           , ZN => n1679);
   U1002 : AOI211_X1 port map( C1 => n2170, C2 => DATA1(30), A => n1680, B => 
                           n1679, ZN => n1681);
   U1003 : INV_X1 port map( A => n1681, ZN => n1804);
   U1004 : AOI222_X1 port map( A1 => n2438, A2 => n1804, B1 => n2436, B2 => 
                           n1806, C1 => n2434, C2 => n1682, ZN => n1809);
   U1005 : OAI22_X1 port map( A1 => n2442, A2 => n1810, B1 => n2440, B2 => 
                           n1809, ZN => n1683);
   U1006 : INV_X1 port map( A => n1683, ZN => n1686);
   U1007 : AOI22_X1 port map( A1 => n1761, A2 => n1813, B1 => n1814, B2 => 
                           n1684, ZN => n1685);
   U1008 : OAI211_X1 port map( C1 => n1807, C2 => n1687, A => n1686, B => n1685
                           , ZN => n1817);
   U1009 : AOI22_X1 port map( A1 => n2397, A2 => n1817, B1 => n2342, B2 => 
                           n1822, ZN => n1690);
   U1010 : AOI22_X1 port map( A1 => n1823, A2 => n1818, B1 => n1902, B2 => 
                           n1688, ZN => n1689);
   U1011 : OAI211_X1 port map( C1 => n1816, C2 => n1750, A => n1690, B => n1689
                           , ZN => n1800);
   U1012 : AOI222_X1 port map( A1 => n1692, A2 => n1907, B1 => n1691, B2 => 
                           n2281, C1 => n1800, C2 => n2317, ZN => n1834);
   U1013 : OAI22_X1 port map( A1 => n1829, A2 => n2480, B1 => n2283, B2 => 
                           n1834, ZN => n1694);
   U1014 : OAI22_X1 port map( A1 => n1695, A2 => n1957, B1 => n1830, B2 => 
                           n2230, ZN => n1693);
   U1015 : AOI211_X1 port map( C1 => n2473, C2 => n1828, A => n1694, B => n1693
                           , ZN => n1838);
   U1016 : OAI22_X1 port map( A1 => n1790, A2 => n1961, B1 => n1838, B2 => 
                           n2375, ZN => n1703);
   U1017 : INV_X1 port map( A => n1830, ZN => n1698);
   U1018 : OAI22_X1 port map( A1 => n1695, A2 => n2230, B1 => n1829, B2 => 
                           n2254, ZN => n1697);
   U1019 : OAI22_X1 port map( A1 => n1715, A2 => n2480, B1 => n1957, B2 => 
                           n1734, ZN => n1696);
   U1020 : AOI211_X1 port map( C1 => n2472, C2 => n1698, A => n1697, B => n1696
                           , ZN => n1837);
   U1021 : OAI22_X1 port map( A1 => n1957, A2 => n1733, B1 => n1734, B2 => 
                           n2480, ZN => n1700);
   U1022 : OAI22_X1 port map( A1 => n2283, A2 => n1829, B1 => n1715, B2 => 
                           n2230, ZN => n1699);
   U1023 : AOI211_X1 port map( C1 => n2473, C2 => n1701, A => n1700, B => n1699
                           , ZN => n1842);
   U1024 : OAI22_X1 port map( A1 => n1837, A2 => n2118, B1 => n1842, B2 => 
                           n2112, ZN => n1702);
   U1025 : AOI211_X1 port map( C1 => n2386, C2 => n1835, A => n1703, B => n1702
                           , ZN => n1799);
   U1026 : INV_X1 port map( A => n1842, ZN => n1739);
   U1027 : AOI22_X1 port map( A1 => n1739, A2 => n2483, B1 => n1835, B2 => 
                           n2481, ZN => n1719);
   U1028 : INV_X1 port map( A => n1777, ZN => n1760);
   U1029 : OAI222_X1 port map( A1 => n1725, A2 => n1704, B1 => n1723, B2 => 
                           n1724, C1 => n1721, C2 => n1722, ZN => n1740);
   U1030 : AOI22_X1 port map( A1 => n2125, A2 => n1744, B1 => n1814, B2 => 
                           n1740, ZN => n1707);
   U1031 : AOI22_X1 port map( A1 => n1761, A2 => n1743, B1 => n2449, B2 => 
                           n1705, ZN => n1706);
   U1032 : OAI211_X1 port map( C1 => n2440, C2 => n1708, A => n1707, B => n1706
                           , ZN => n1768);
   U1033 : INV_X1 port map( A => n1768, ZN => n1751);
   U1034 : OAI22_X1 port map( A1 => n1750, A2 => n1731, B1 => n2456, B2 => 
                           n1751, ZN => n1712);
   U1035 : OAI22_X1 port map( A1 => n2454, A2 => n1710, B1 => n2452, B2 => 
                           n1709, ZN => n1711);
   U1036 : AOI211_X1 port map( C1 => n1752, C2 => n1823, A => n1712, B => n1711
                           , ZN => n1713);
   U1037 : INV_X1 port map( A => n1713, ZN => n1756);
   U1038 : AOI222_X1 port map( A1 => n1756, A2 => n1907, B1 => n1732, B2 => 
                           n2281, C1 => n1714, C2 => n2317, ZN => n1776);
   U1039 : OAI22_X1 port map( A1 => n1957, A2 => n1776, B1 => n1733, B2 => 
                           n2230, ZN => n1717);
   U1040 : OAI22_X1 port map( A1 => n2283, A2 => n1715, B1 => n1734, B2 => 
                           n2254, ZN => n1716);
   U1041 : AOI211_X1 port map( C1 => n2345, C2 => n1760, A => n1717, B => n1716
                           , ZN => n1791);
   U1042 : INV_X1 port map( A => n1791, ZN => n1786);
   U1043 : INV_X1 port map( A => n1790, ZN => n1783);
   U1044 : AOI22_X1 port map( A1 => n1786, A2 => n2487, B1 => n1783, B2 => 
                           n2485, ZN => n1718);
   U1045 : OAI211_X1 port map( C1 => n2492, C2 => n1837, A => n1719, B => n1718
                           , ZN => n1845);
   U1046 : INV_X1 port map( A => n1845, ZN => n1794);
   U1047 : OAI22_X1 port map( A1 => n1791, A2 => n2112, B1 => n1790, B2 => 
                           n2118, ZN => n1738);
   U1048 : INV_X1 port map( A => n1776, ZN => n1775);
   U1049 : AOI22_X1 port map( A1 => n1762, A2 => n1743, B1 => n2183, B2 => 
                           n1740, ZN => n1727);
   U1050 : OAI222_X1 port map( A1 => n1725, A2 => n1724, B1 => n1723, B2 => 
                           n1722, C1 => n1721, C2 => n1720, ZN => n1894);
   U1051 : AOI22_X1 port map( A1 => n2449, A2 => n1744, B1 => n1814, B2 => 
                           n1894, ZN => n1726);
   U1052 : OAI211_X1 port map( C1 => n2440, C2 => n1728, A => n1727, B => n1726
                           , ZN => n1767);
   U1053 : AOI22_X1 port map( A1 => n2461, A2 => n1753, B1 => n1902, B2 => 
                           n1767, ZN => n1730);
   U1054 : AOI22_X1 port map( A1 => n2342, A2 => n1752, B1 => n2332, B2 => 
                           n1768, ZN => n1729);
   U1055 : OAI211_X1 port map( C1 => n1731, C2 => n2454, A => n1730, B => n1729
                           , ZN => n1757);
   U1056 : AOI222_X1 port map( A1 => n1757, A2 => n1907, B1 => n1756, B2 => 
                           n2281, C1 => n1732, C2 => n2317, ZN => n1893);
   U1057 : OAI22_X1 port map( A1 => n1957, A2 => n1893, B1 => n1777, B2 => 
                           n2230, ZN => n1736);
   U1058 : OAI22_X1 port map( A1 => n2283, A2 => n1734, B1 => n1733, B2 => 
                           n2254, ZN => n1735);
   U1059 : AOI211_X1 port map( C1 => n2345, C2 => n1775, A => n1736, B => n1735
                           , ZN => n1785);
   U1060 : OAI22_X1 port map( A1 => n1785, A2 => n1961, B1 => n1837, B2 => 
                           n2375, ZN => n1737);
   U1061 : AOI211_X1 port map( C1 => n2386, C2 => n1739, A => n1738, B => n1737
                           , ZN => n1797);
   U1062 : OAI222_X1 port map( A1 => n2079, A2 => n1799, B1 => n2066, B2 => 
                           n1794, C1 => n1797, C2 => n1963, ZN => n1891);
   U1063 : INV_X1 port map( A => n1740, ZN => n1766);
   U1064 : AOI22_X1 port map( A1 => n1762, A2 => n1894, B1 => n1745, B2 => 
                           n1743, ZN => n1742);
   U1065 : AOI22_X1 port map( A1 => n1761, A2 => n1763, B1 => n1814, B2 => 
                           n1898, ZN => n1741);
   U1066 : OAI211_X1 port map( C1 => n1766, C2 => n2178, A => n1742, B => n1741
                           , ZN => n2343);
   U1067 : AOI22_X1 port map( A1 => n2342, A2 => n1767, B1 => n1902, B2 => 
                           n2343, ZN => n1749);
   U1068 : AOI22_X1 port map( A1 => n1761, A2 => n1894, B1 => n2449, B2 => 
                           n1743, ZN => n1747);
   U1069 : AOI22_X1 port map( A1 => n1814, A2 => n1763, B1 => n1745, B2 => 
                           n1744, ZN => n1746);
   U1070 : OAI211_X1 port map( C1 => n1766, C2 => n2442, A => n1747, B => n1746
                           , ZN => n2331);
   U1071 : AOI22_X1 port map( A1 => n2397, A2 => n1752, B1 => n2332, B2 => 
                           n2331, ZN => n1748);
   U1072 : OAI211_X1 port map( C1 => n1751, C2 => n1750, A => n1749, B => n1748
                           , ZN => n1906);
   U1073 : INV_X1 port map( A => n1767, ZN => n1905);
   U1074 : AOI22_X1 port map( A1 => n2342, A2 => n1768, B1 => n1902, B2 => 
                           n2331, ZN => n1755);
   U1075 : AOI22_X1 port map( A1 => n2397, A2 => n1753, B1 => n2461, B2 => 
                           n1752, ZN => n1754);
   U1076 : OAI211_X1 port map( C1 => n1905, C2 => n2458, A => n1755, B => n1754
                           , ZN => n1772);
   U1077 : AOI222_X1 port map( A1 => n1906, A2 => n1907, B1 => n1772, B2 => 
                           n2281, C1 => n1757, C2 => n2317, ZN => n2231);
   U1078 : OAI22_X1 port map( A1 => n1957, A2 => n2231, B1 => n1893, B2 => 
                           n2230, ZN => n1759);
   U1079 : AOI222_X1 port map( A1 => n1772, A2 => n1907, B1 => n1757, B2 => 
                           n2281, C1 => n1756, C2 => n2317, ZN => n2217);
   U1080 : OAI22_X1 port map( A1 => n1776, A2 => n2254, B1 => n2217, B2 => 
                           n2480, ZN => n1758);
   U1081 : AOI211_X1 port map( C1 => n2472, C2 => n1760, A => n1759, B => n1758
                           , ZN => n2119);
   U1082 : INV_X1 port map( A => n2119, ZN => n1784);
   U1083 : INV_X1 port map( A => n2343, ZN => n1771);
   U1084 : AOI22_X1 port map( A1 => n1896, A2 => n1897, B1 => n1894, B2 => 
                           n2449, ZN => n1765);
   U1085 : AOI22_X1 port map( A1 => n1763, A2 => n1762, B1 => n1898, B2 => 
                           n1761, ZN => n1764);
   U1086 : OAI211_X1 port map( C1 => n2440, C2 => n1766, A => n1765, B => n1764
                           , ZN => n2364);
   U1087 : AOI22_X1 port map( A1 => n1902, A2 => n2364, B1 => n2331, B2 => 
                           n2342, ZN => n1770);
   U1088 : AOI22_X1 port map( A1 => n1768, A2 => n2397, B1 => n1767, B2 => 
                           n2461, ZN => n1769);
   U1089 : OAI211_X1 port map( C1 => n2458, C2 => n1771, A => n1770, B => n1769
                           , ZN => n2282);
   U1090 : AOI222_X1 port map( A1 => n2281, A2 => n1906, B1 => n2317, B2 => 
                           n1772, C1 => n2282, C2 => n1907, ZN => n2255);
   U1091 : OAI22_X1 port map( A1 => n2230, A2 => n2217, B1 => n1957, B2 => 
                           n2255, ZN => n1774);
   U1092 : OAI22_X1 port map( A1 => n2254, A2 => n1893, B1 => n2480, B2 => 
                           n2231, ZN => n1773);
   U1093 : AOI211_X1 port map( C1 => n2472, C2 => n1775, A => n1774, B => n1773
                           , ZN => n2141);
   U1094 : OAI22_X1 port map( A1 => n2230, A2 => n1776, B1 => n1957, B2 => 
                           n2217, ZN => n1779);
   U1095 : OAI22_X1 port map( A1 => n2254, A2 => n1777, B1 => n2480, B2 => 
                           n1893, ZN => n1778);
   U1096 : AOI211_X1 port map( C1 => n2472, C2 => n1780, A => n1779, B => n1778
                           , ZN => n2111);
   U1097 : OAI22_X1 port map( A1 => n1961, A2 => n2141, B1 => n2118, B2 => 
                           n2111, ZN => n1782);
   U1098 : OAI22_X1 port map( A1 => n2492, A2 => n1785, B1 => n2375, B2 => 
                           n1791, ZN => n1781);
   U1099 : AOI211_X1 port map( C1 => n1784, C2 => n2485, A => n1782, B => n1781
                           , ZN => n2065);
   U1100 : AOI22_X1 port map( A1 => n2487, A2 => n1784, B1 => n2481, B2 => 
                           n1783, ZN => n1788);
   U1101 : INV_X1 port map( A => n1785, ZN => n1913);
   U1102 : AOI22_X1 port map( A1 => n2386, A2 => n1786, B1 => n2483, B2 => 
                           n1913, ZN => n1787);
   U1103 : OAI211_X1 port map( C1 => n2111, C2 => n2112, A => n1788, B => n1787
                           , ZN => n1789);
   U1104 : INV_X1 port map( A => n1789, ZN => n1914);
   U1105 : OAI22_X1 port map( A1 => n1961, A2 => n2111, B1 => n2492, B2 => 
                           n1790, ZN => n1793);
   U1106 : OAI22_X1 port map( A1 => n2118, A2 => n1791, B1 => n2375, B2 => 
                           n1842, ZN => n1792);
   U1107 : AOI211_X1 port map( C1 => n1913, C2 => n2485, A => n1793, B => n1792
                           , ZN => n1796);
   U1108 : OAI222_X1 port map( A1 => n2065, A2 => n1963, B1 => n1914, B2 => 
                           n2066, C1 => n1796, C2 => n2079, ZN => n2029);
   U1109 : OAI222_X1 port map( A1 => n1796, A2 => n1963, B1 => n1797, B2 => 
                           n2066, C1 => n1794, C2 => n2079, ZN => n1980);
   U1110 : INV_X1 port map( A => n2202, ZN => n2501);
   U1111 : AOI22_X1 port map( A1 => n2029, A2 => n2507, B1 => n1980, B2 => 
                           n2501, ZN => n1795);
   U1112 : INV_X1 port map( A => n1795, ZN => n1849);
   U1113 : OAI222_X1 port map( A1 => n1914, A2 => n1963, B1 => n1797, B2 => 
                           n2079, C1 => n1796, C2 => n2066, ZN => n2002);
   U1114 : INV_X1 port map( A => n2002, ZN => n1847);
   U1115 : INV_X1 port map( A => n2507, ZN => n1888);
   U1116 : NAND3_X1 port map( A1 => DATA2(0), A2 => n1798, A3 => n1888, ZN => 
                           n1892);
   U1117 : INV_X1 port map( A => n1799, ZN => n1844);
   U1118 : INV_X1 port map( A => n1800, ZN => n1826);
   U1119 : AOI22_X1 port map( A1 => DATA1(28), A2 => n1801, B1 => DATA1(27), B2
                           => n2431, ZN => n1803);
   U1120 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(30), ZN => n1990);
   U1121 : NAND2_X1 port map( A1 => n2170, A2 => DATA1(31), ZN => n1880);
   U1122 : NAND4_X1 port map( A1 => n1803, A2 => n1802, A3 => n1990, A4 => 
                           n1880, ZN => n1805);
   U1123 : AOI222_X1 port map( A1 => n1806, A2 => n2434, B1 => n1805, B2 => 
                           n2438, C1 => n1804, C2 => n2436, ZN => n1808);
   U1124 : OAI22_X1 port map( A1 => n2440, A2 => n1808, B1 => n1807, B2 => 
                           n2442, ZN => n1812);
   U1125 : OAI22_X1 port map( A1 => n1810, A2 => n2446, B1 => n1809, B2 => 
                           n2178, ZN => n1811);
   U1126 : AOI211_X1 port map( C1 => n1814, C2 => n1813, A => n1812, B => n1811
                           , ZN => n1815);
   U1127 : OAI22_X1 port map( A1 => n1816, A2 => n2452, B1 => n1815, B2 => 
                           n2454, ZN => n1821);
   U1128 : AOI22_X1 port map( A1 => n1902, A2 => n1818, B1 => n1817, B2 => 
                           n2461, ZN => n1819);
   U1129 : INV_X1 port map( A => n1819, ZN => n1820);
   U1130 : AOI211_X1 port map( C1 => n1823, C2 => n1822, A => n1821, B => n1820
                           , ZN => n1825);
   U1131 : OAI222_X1 port map( A1 => n2465, A2 => n1826, B1 => n2463, B2 => 
                           n1825, C1 => n1824, C2 => n2467, ZN => n1827);
   U1132 : AOI22_X1 port map( A1 => n2469, A2 => n1828, B1 => n2472, B2 => 
                           n1827, ZN => n1833);
   U1133 : OAI22_X1 port map( A1 => n2480, A2 => n1830, B1 => n1829, B2 => 
                           n1957, ZN => n1831);
   U1134 : INV_X1 port map( A => n1831, ZN => n1832);
   U1135 : OAI211_X1 port map( C1 => n1834, C2 => n2254, A => n1833, B => n1832
                           , ZN => n1836);
   U1136 : AOI22_X1 port map( A1 => n2481, A2 => n1836, B1 => n2483, B2 => 
                           n1835, ZN => n1841);
   U1137 : OAI22_X1 port map( A1 => n2492, A2 => n1838, B1 => n2112, B2 => 
                           n1837, ZN => n1839);
   U1138 : INV_X1 port map( A => n1839, ZN => n1840);
   U1139 : OAI211_X1 port map( C1 => n1842, C2 => n1961, A => n1841, B => n1840
                           , ZN => n1843);
   U1140 : AOI222_X1 port map( A1 => n1845, A2 => n2493, B1 => n1844, B2 => 
                           n2498, C1 => n1843, C2 => n2496, ZN => n1846);
   U1141 : OAI22_X1 port map( A1 => n1847, A2 => n1892, B1 => n1846, B2 => 
                           n1917, ZN => n1848);
   U1142 : AOI211_X1 port map( C1 => n2198, C2 => n1891, A => n1849, B => n1848
                           , ZN => n1921);
   U1143 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n1866);
   U1144 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => 
                           n1866, ZN => n2108);
   U1145 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n2109);
   U1146 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n1863);
   U1147 : INV_X1 port map( A => n1863, ZN => n2103);
   U1148 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n2099);
   U1149 : OAI21_X1 port map( B1 => DATA1(17), B2 => DATA2_I_17_port, A => 
                           n2099, ZN => n2259);
   U1150 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n2100);
   U1151 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => 
                           n2100, ZN => n2234);
   U1152 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n2101);
   U1153 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => 
                           n2101, ZN => n2227);
   U1154 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n2260);
   U1155 : OAI21_X1 port map( B1 => DATA1(16), B2 => DATA2_I_16_port, A => 
                           n2260, ZN => n2278);
   U1156 : NOR4_X1 port map( A1 => n2259, A2 => n2234, A3 => n2227, A4 => n2278
                           , ZN => n1862);
   U1157 : NAND2_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, ZN => 
                           n2289);
   U1158 : OAI21_X1 port map( B1 => DATA1(14), B2 => DATA2_I_14_port, A => 
                           n2289, ZN => n2323);
   U1159 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n1853);
   U1160 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => 
                           n1853, ZN => n2330);
   U1161 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n2329);
   U1162 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => 
                           n2329, ZN => n1854);
   U1163 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n2287);
   U1164 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n2287, ZN => n2373);
   U1165 : NOR4_X1 port map( A1 => n2323, A2 => n2330, A3 => n1854, A4 => n2373
                           , ZN => n1858);
   U1166 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n2286);
   U1167 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n2286, ZN => n2404);
   U1168 : NOR4_X1 port map( A1 => n1852, A2 => n1851, A3 => n2404, A4 => n1850
                           , ZN => n1857);
   U1169 : INV_X1 port map( A => n1853, ZN => n2311);
   U1170 : INV_X1 port map( A => n1854, ZN => n2360);
   U1171 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n1856);
   U1172 : INV_X1 port map( A => n1855, ZN => n2400);
   U1173 : AOI21_X1 port map( B1 => n2391, B2 => n2400, A => n2404, ZN => n2389
                           );
   U1174 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => DATA1(10), A => 
                           n2389, ZN => n2374);
   U1175 : OAI21_X1 port map( B1 => n1856, B2 => n2374, A => n2287, ZN => n2359
                           );
   U1176 : NAND2_X1 port map( A1 => n2360, A2 => n2359, ZN => n2357);
   U1177 : AOI21_X1 port map( B1 => n2329, B2 => n2357, A => n2330, ZN => n2306
                           );
   U1178 : NOR2_X1 port map( A1 => n2311, A2 => n2306, ZN => n2305);
   U1179 : OAI21_X1 port map( B1 => n2305, B2 => n2323, A => n2289, ZN => n2298
                           );
   U1180 : AOI21_X1 port map( B1 => n1858, B2 => n1857, A => n2298, ZN => n1860
                           );
   U1181 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n1859);
   U1182 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => 
                           n1859, ZN => n2297);
   U1183 : OAI21_X1 port map( B1 => n1860, B2 => n2297, A => n1859, ZN => n2098
                           );
   U1184 : NOR2_X1 port map( A1 => n2260, A2 => n2259, ZN => n2258);
   U1185 : AOI21_X1 port map( B1 => DATA2_I_17_port, B2 => DATA1(17), A => 
                           n2258, ZN => n2235);
   U1186 : NOR2_X1 port map( A1 => n2235, A2 => n2234, ZN => n2233);
   U1187 : AOI21_X1 port map( B1 => DATA2_I_18_port, B2 => DATA1(18), A => 
                           n2233, ZN => n2216);
   U1188 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n1861);
   U1189 : OAI21_X1 port map( B1 => n2216, B2 => n1861, A => n2101, ZN => n2152
                           );
   U1190 : AOI21_X1 port map( B1 => n1862, B2 => n2098, A => n2152, ZN => n1864
                           );
   U1191 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n2102);
   U1192 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n2102, ZN => n2164);
   U1193 : OAI21_X1 port map( B1 => DATA1(21), B2 => DATA2_I_21_port, A => 
                           n1863, ZN => n2149);
   U1194 : AOI221_X1 port map( B1 => n1864, B2 => n2102, C1 => n2164, C2 => 
                           n2102, A => n2149, ZN => n1865);
   U1195 : XOR2_X1 port map( A => n2126, B => DATA2_I_22_port, Z => n2135);
   U1196 : INV_X1 port map( A => n2135, ZN => n2137);
   U1197 : OAI21_X1 port map( B1 => n2103, B2 => n1865, A => n2137, ZN => n1867
                           );
   U1198 : OAI221_X1 port map( B1 => n2108, B2 => n2109, C1 => n2108, C2 => 
                           n1867, A => n1866, ZN => n1872);
   U1199 : NAND2_X1 port map( A1 => n2696, A2 => n1872, ZN => n2069);
   U1200 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n1877);
   U1201 : NAND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => 
                           n1870);
   U1202 : INV_X1 port map( A => n1870, ZN => n1932);
   U1203 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n1986);
   U1204 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n1869);
   U1205 : INV_X1 port map( A => n1869, ZN => n2019);
   U1206 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n2034);
   U1207 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n1868);
   U1208 : INV_X1 port map( A => n1868, ZN => n2059);
   U1209 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n2090);
   U1210 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => 
                           n1868, ZN => n2071);
   U1211 : NOR2_X1 port map( A1 => n2090, A2 => n2071, ZN => n2070);
   U1212 : XOR2_X1 port map( A => DATA1(26), B => DATA2_I_26_port, Z => n2058);
   U1213 : OAI21_X1 port map( B1 => n2059, B2 => n2070, A => n2058, ZN => n2023
                           );
   U1214 : OAI21_X1 port map( B1 => DATA1(27), B2 => DATA2_I_27_port, A => 
                           n1869, ZN => n2035);
   U1215 : AOI21_X1 port map( B1 => n2034, B2 => n2023, A => n2035, ZN => n2024
                           );
   U1216 : XNOR2_X1 port map( A => n2675, B => DATA2_I_28_port, ZN => n2018);
   U1217 : OAI21_X1 port map( B1 => n2019, B2 => n2024, A => n2018, ZN => n2003
                           );
   U1218 : OAI21_X1 port map( B1 => DATA1(29), B2 => DATA2_I_29_port, A => 
                           n1870, ZN => n1985);
   U1219 : AOI21_X1 port map( B1 => n1986, B2 => n2003, A => n1985, ZN => n1924
                           );
   U1220 : XOR2_X1 port map( A => DATA1(30), B => DATA2_I_30_port, Z => n1933);
   U1221 : OAI21_X1 port map( B1 => n1932, B2 => n1924, A => n1933, ZN => n1875
                           );
   U1222 : INV_X1 port map( A => n2071, ZN => n1871);
   U1223 : NAND3_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, A3 => 
                           n1871, ZN => n2062);
   U1224 : INV_X1 port map( A => n2062, ZN => n2068);
   U1225 : OAI21_X1 port map( B1 => n2059, B2 => n2068, A => n2058, ZN => n2031
                           );
   U1226 : AOI21_X1 port map( B1 => n2034, B2 => n2031, A => n2035, ZN => n2032
                           );
   U1227 : OAI21_X1 port map( B1 => n2019, B2 => n2032, A => n2018, ZN => n1982
                           );
   U1228 : AOI21_X1 port map( B1 => n1986, B2 => n1982, A => n1985, ZN => n1922
                           );
   U1229 : OAI21_X1 port map( B1 => n1932, B2 => n1922, A => n1933, ZN => n1876
                           );
   U1230 : NOR2_X1 port map( A1 => n3038, A2 => n1872, ZN => n2083);
   U1231 : INV_X1 port map( A => n2083, ZN => n2067);
   U1232 : AOI21_X1 port map( B1 => n1877, B2 => n1876, A => n2067, ZN => n1873
                           );
   U1233 : INV_X1 port map( A => n1873, ZN => n1874);
   U1234 : OAI221_X1 port map( B1 => n2069, B2 => n1877, C1 => n2069, C2 => 
                           n1875, A => n1874, ZN => n1886);
   U1235 : INV_X1 port map( A => DATA1(31), ZN => n2599);
   U1236 : XOR2_X1 port map( A => n2599, B => DATA2_I_31_port, Z => n1885);
   U1237 : INV_X1 port map( A => n2069, ZN => n2089);
   U1238 : NAND2_X1 port map( A1 => n2089, A2 => n1875, ZN => n1927);
   U1239 : NAND2_X1 port map( A1 => n2083, A2 => n1876, ZN => n1936);
   U1240 : NAND2_X1 port map( A1 => n1927, A2 => n1936, ZN => n1931);
   U1241 : NAND2_X1 port map( A1 => n1877, A2 => n1931, ZN => n1883);
   U1242 : OAI221_X1 port map( B1 => DATA1(31), B2 => n2416, C1 => n2599, C2 =>
                           n2412, A => n2392, ZN => n1878);
   U1243 : NOR2_X1 port map( A1 => DATA2(31), A2 => n2599, ZN => n2679);
   U1244 : AOI22_X1 port map( A1 => DATA2(31), A2 => n1878, B1 => n2679, B2 => 
                           n2393, ZN => n1879);
   U1245 : OAI21_X1 port map( B1 => n1880, B2 => n2409, A => n1879, ZN => n1881
                           );
   U1246 : AOI21_X1 port map( B1 => n2422, B2 => dataout_mul_31_port, A => 
                           n1881, ZN => n1882);
   U1247 : OAI21_X1 port map( B1 => n1883, B2 => n1885, A => n1882, ZN => n1884
                           );
   U1248 : AOI21_X1 port map( B1 => n1886, B2 => n1885, A => n1884, ZN => n1920
                           );
   U1249 : OR3_X1 port map( A1 => n2730, A2 => n1888, A3 => n1887, ZN => n1889)
                           ;
   U1250 : NOR2_X1 port map( A1 => n1890, A2 => n1889, ZN => n2690);
   U1251 : INV_X1 port map( A => n1891, ZN => n1918);
   U1252 : INV_X1 port map( A => n1892, ZN => n2505);
   U1253 : AOI22_X1 port map( A1 => n2505, A2 => n2029, B1 => n2198, B2 => 
                           n1980, ZN => n1916);
   U1254 : INV_X1 port map( A => n1893, ZN => n1910);
   U1255 : AOI22_X1 port map( A1 => n1896, A2 => n1895, B1 => n2121, B2 => 
                           n1894, ZN => n1900);
   U1256 : AOI22_X1 port map( A1 => n2125, A2 => n1898, B1 => n2183, B2 => 
                           n1897, ZN => n1899);
   U1257 : OAI211_X1 port map( C1 => n1901, C2 => n2178, A => n1900, B => n1899
                           , ZN => n2395);
   U1258 : AOI22_X1 port map( A1 => n2342, A2 => n2343, B1 => n1902, B2 => 
                           n2395, ZN => n1904);
   U1259 : AOI22_X1 port map( A1 => n2461, A2 => n2331, B1 => n2332, B2 => 
                           n2364, ZN => n1903);
   U1260 : OAI211_X1 port map( C1 => n1905, C2 => n2454, A => n1904, B => n1903
                           , ZN => n2316);
   U1261 : AOI222_X1 port map( A1 => n2316, A2 => n1907, B1 => n2282, B2 => 
                           n2281, C1 => n1906, C2 => n2317, ZN => n2268);
   U1262 : OAI22_X1 port map( A1 => n1957, A2 => n2268, B1 => n2231, B2 => 
                           n2230, ZN => n1909);
   U1263 : OAI22_X1 port map( A1 => n2217, A2 => n2254, B1 => n2255, B2 => 
                           n2480, ZN => n1908);
   U1264 : AOI211_X1 port map( C1 => n2472, C2 => n1910, A => n1909, B => n1908
                           , ZN => n2156);
   U1265 : OAI22_X1 port map( A1 => n2119, A2 => n2118, B1 => n2156, B2 => 
                           n1961, ZN => n1912);
   U1266 : OAI22_X1 port map( A1 => n2111, A2 => n2492, B1 => n2141, B2 => 
                           n2112, ZN => n1911);
   U1267 : AOI211_X1 port map( C1 => n2481, C2 => n1913, A => n1912, B => n1911
                           , ZN => n2080);
   U1268 : OAI222_X1 port map( A1 => n2066, A2 => n2065, B1 => n2079, B2 => 
                           n1914, C1 => n2080, C2 => n1963, ZN => n2046);
   U1269 : AOI22_X1 port map( A1 => n2507, A2 => n2046, B1 => n2501, B2 => 
                           n2002, ZN => n1915);
   U1270 : OAI211_X1 port map( C1 => n1918, C2 => n1917, A => n1916, B => n1915
                           , ZN => n1930);
   U1271 : NAND3_X1 port map( A1 => n2690, A2 => n2695, A3 => n1930, ZN => 
                           n1919);
   U1272 : OAI211_X1 port map( C1 => n1921, C2 => n2382, A => n1920, B => n1919
                           , ZN => OUTALU(31));
   U1273 : INV_X1 port map( A => n1922, ZN => n1981);
   U1274 : INV_X1 port map( A => DATA2(30), ZN => n2698);
   U1275 : AOI22_X1 port map( A1 => DATA1(30), A2 => n2698, B1 => DATA2(30), B2
                           => n2535_port, ZN => n2678);
   U1276 : AOI21_X1 port map( B1 => DATA1(30), B2 => n2367, A => n2365, ZN => 
                           n1923);
   U1277 : OAI22_X1 port map( A1 => n2678, A2 => n2416, B1 => n1923, B2 => 
                           n2698, ZN => n1929);
   U1278 : INV_X1 port map( A => n1924, ZN => n1983);
   U1279 : OAI22_X1 port map( A1 => n1937, A2 => n2599, B1 => n2428, B2 => 
                           n2535_port, ZN => n1925);
   U1280 : AOI22_X1 port map( A1 => n2688, A2 => n1925, B1 => n2314, B2 => 
                           dataout_mul_30_port, ZN => n1926);
   U1281 : OAI21_X1 port map( B1 => n1983, B2 => n1927, A => n1926, ZN => n1928
                           );
   U1282 : AOI211_X1 port map( C1 => n2396, C2 => n1930, A => n1929, B => n1928
                           , ZN => n1935);
   U1283 : OAI21_X1 port map( B1 => n1933, B2 => n1932, A => n1931, ZN => n1934
                           );
   U1284 : OAI211_X1 port map( C1 => n1936, C2 => n1981, A => n1935, B => n1934
                           , ZN => OUTALU(30));
   U1285 : NOR2_X1 port map( A1 => n2428, A2 => n2611, ZN => n1941);
   U1286 : NOR2_X1 port map( A1 => n1937, A2 => n2604, ZN => n2430);
   U1287 : AOI211_X1 port map( C1 => DATA1(0), C2 => n2006, A => n1941, B => 
                           n2430, ZN => n1979);
   U1288 : OAI22_X1 port map( A1 => n1969, A2 => n2415, B1 => n1971, B2 => 
                           n1938, ZN => n1939);
   U1289 : AOI22_X1 port map( A1 => dataout_mul_2_port, A2 => n2422, B1 => 
                           n1972, B2 => n1939, ZN => n1978);
   U1290 : OAI21_X1 port map( B1 => n2611, B2 => n2412, A => n2392, ZN => n1976
                           );
   U1291 : AOI22_X1 port map( A1 => n2501, A2 => n2506, B1 => n2198, B2 => 
                           n2504, ZN => n1968);
   U1292 : AOI22_X1 port map( A1 => n2386, A2 => n2486, B1 => n2485, B2 => 
                           n2192, ZN => n1960);
   U1293 : INV_X1 port map( A => n2457, ZN => n1952);
   U1294 : INV_X1 port map( A => n2179, ZN => n1948);
   U1295 : AOI211_X1 port map( C1 => DATA1(6), C2 => n2431, A => n1941, B => 
                           n1940, ZN => n1943);
   U1296 : OAI211_X1 port map( C1 => n1991, C2 => n2613, A => n1943, B => n1942
                           , ZN => n2433);
   U1297 : AOI222_X1 port map( A1 => n1944, A2 => n2434, B1 => n2433, B2 => 
                           n2438, C1 => n2177, C2 => n2436, ZN => n2441);
   U1298 : OAI22_X1 port map( A1 => n2440, A2 => n2441, B1 => n2443, B2 => 
                           n2442, ZN => n1947);
   U1299 : OAI22_X1 port map( A1 => n2444, A2 => n1945, B1 => n2445, B2 => 
                           n2178, ZN => n1946);
   U1300 : AOI211_X1 port map( C1 => n2183, C2 => n1948, A => n1947, B => n1946
                           , ZN => n2451);
   U1301 : OAI22_X1 port map( A1 => n2455, A2 => n2452, B1 => n2451, B2 => 
                           n2454, ZN => n1951);
   U1302 : OAI22_X1 port map( A1 => n2456, A2 => n1949, B1 => n2184, B2 => 
                           n2458, ZN => n1950);
   U1303 : AOI211_X1 port map( C1 => n2461, C2 => n1952, A => n1951, B => n1950
                           , ZN => n2468);
   U1304 : OAI222_X1 port map( A1 => n2465, A2 => n2188, B1 => n2463, B2 => 
                           n2468, C1 => n1953, C2 => n2467, ZN => n2470);
   U1305 : AOI22_X1 port map( A1 => n2345, A2 => n2189, B1 => n2472, B2 => 
                           n2470, ZN => n1955);
   U1306 : AOI22_X1 port map( A1 => n2473, A2 => n2171, B1 => n2469, B2 => 
                           n2475, ZN => n1954);
   U1307 : OAI211_X1 port map( C1 => n1957, C2 => n1956, A => n1955, B => n1954
                           , ZN => n2484);
   U1308 : INV_X1 port map( A => n1958, ZN => n2488);
   U1309 : AOI22_X1 port map( A1 => n2481, A2 => n2484, B1 => n2483, B2 => 
                           n2488, ZN => n1959);
   U1310 : OAI211_X1 port map( C1 => n1962, C2 => n1961, A => n1960, B => n1959
                           , ZN => n2494);
   U1311 : INV_X1 port map( A => n2494, ZN => n1965);
   U1312 : OAI222_X1 port map( A1 => n2066, A2 => n1966, B1 => n2079, B2 => 
                           n1965, C1 => n1964, C2 => n1963, ZN => n2500);
   U1313 : AOI22_X1 port map( A1 => n2503, A2 => n2500, B1 => n2505, B2 => 
                           n2199, ZN => n1967);
   U1314 : AOI21_X1 port map( B1 => n1968, B2 => n1967, A => n2409, ZN => n1975
                           );
   U1315 : AOI22_X1 port map( A1 => DATA2(2), A2 => n2611, B1 => DATA1(2), B2 
                           => n2728, ZN => n2606);
   U1316 : AOI22_X1 port map( A1 => n2420, A2 => n1971, B1 => n1970, B2 => 
                           n1969, ZN => n1973);
   U1317 : OAI22_X1 port map( A1 => n2606, A2 => n2416, B1 => n1973, B2 => 
                           n1972, ZN => n1974);
   U1318 : AOI211_X1 port map( C1 => DATA2(2), C2 => n1976, A => n1975, B => 
                           n1974, ZN => n1977);
   U1319 : OAI211_X1 port map( C1 => n1979, C2 => n2382, A => n1978, B => n1977
                           , ZN => OUTALU(2));
   U1320 : AOI22_X1 port map( A1 => n2503, A2 => n1980, B1 => n2501, B2 => 
                           n2029, ZN => n2001);
   U1321 : AOI22_X1 port map( A1 => n2198, A2 => n2002, B1 => n2505, B2 => 
                           n2046, ZN => n2000);
   U1322 : NAND2_X1 port map( A1 => n1981, A2 => n2083, ZN => n1984);
   U1323 : INV_X1 port map( A => n1984, ZN => n1998);
   U1324 : INV_X1 port map( A => n1982, ZN => n2015);
   U1325 : NAND2_X1 port map( A1 => n2089, A2 => n1983, ZN => n1995);
   U1326 : AOI22_X1 port map( A1 => n1986, A2 => n1985, B1 => n1984, B2 => 
                           n1995, ZN => n1997);
   U1327 : INV_X1 port map( A => DATA1(29), ZN => n1987);
   U1328 : NAND2_X1 port map( A1 => DATA2(29), A2 => n1987, ZN => n2677);
   U1329 : INV_X1 port map( A => DATA2(29), ZN => n2699);
   U1330 : NAND2_X1 port map( A1 => DATA1(29), A2 => n2699, ZN => n2674);
   U1331 : NAND2_X1 port map( A1 => n2677, A2 => n2674, ZN => n2522_port);
   U1332 : OAI21_X1 port map( B1 => n1987, B2 => n2412, A => n2392, ZN => n1988
                           );
   U1333 : AOI22_X1 port map( A1 => n2393, A2 => n2522_port, B1 => DATA2(29), 
                           B2 => n1988, ZN => n1994);
   U1334 : OAI211_X1 port map( C1 => n1991, C2 => n2599, A => n1990, B => n1989
                           , ZN => n1992);
   U1335 : AOI22_X1 port map( A1 => n2688, A2 => n1992, B1 => n2314, B2 => 
                           dataout_mul_29_port, ZN => n1993);
   U1336 : OAI211_X1 port map( C1 => n2003, C2 => n1995, A => n1994, B => n1993
                           , ZN => n1996);
   U1337 : AOI211_X1 port map( C1 => n1998, C2 => n2015, A => n1997, B => n1996
                           , ZN => n1999);
   U1338 : OAI221_X1 port map( B1 => n2382, B2 => n2001, C1 => n2382, C2 => 
                           n2000, A => n1999, ZN => OUTALU(29));
   U1339 : AOI222_X1 port map( A1 => n2002, A2 => n2503, B1 => n2046, B2 => 
                           n2501, C1 => n2029, C2 => n2198, ZN => n2022);
   U1340 : AND2_X1 port map( A1 => n2003, A2 => n2089, ZN => n2016);
   U1341 : INV_X1 port map( A => n2032, ZN => n2004);
   U1342 : NOR3_X1 port map( A1 => n2018, A2 => n2004, A3 => n2067, ZN => n2014
                           );
   U1343 : INV_X1 port map( A => DATA2(28), ZN => n2700);
   U1344 : AOI22_X1 port map( A1 => DATA1(28), A2 => n2700, B1 => DATA2(28), B2
                           => n2675, ZN => n2670);
   U1345 : AOI22_X1 port map( A1 => n2006, A2 => DATA1(30), B1 => n2005, B2 => 
                           DATA1(31), ZN => n2009);
   U1346 : NAND3_X1 port map( A1 => n2009, A2 => n2008, A3 => n2007, ZN => 
                           n2010);
   U1347 : AOI22_X1 port map( A1 => n2688, A2 => n2010, B1 => n2314, B2 => 
                           dataout_mul_28_port, ZN => n2012);
   U1348 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA2(28), B => 
                           DATA1(28), ZN => n2011);
   U1349 : OAI211_X1 port map( C1 => n2670, C2 => n2416, A => n2012, B => n2011
                           , ZN => n2013);
   U1350 : AOI211_X1 port map( C1 => n2016, C2 => n2024, A => n2014, B => n2013
                           , ZN => n2021);
   U1351 : NOR2_X1 port map( A1 => n2015, A2 => n2067, ZN => n2017);
   U1352 : OAI22_X1 port map( A1 => n2019, A2 => n2018, B1 => n2017, B2 => 
                           n2016, ZN => n2020);
   U1353 : OAI211_X1 port map( C1 => n2022, C2 => n2382, A => n2021, B => n2020
                           , ZN => OUTALU(28));
   U1354 : INV_X1 port map( A => n2023, ZN => n2045);
   U1355 : NOR2_X1 port map( A1 => n2024, A2 => n2069, ZN => n2036);
   U1356 : AOI22_X1 port map( A1 => n2045, A2 => n2036, B1 => n2314, B2 => 
                           dataout_mul_27_port, ZN => n2043);
   U1357 : INV_X1 port map( A => DATA2(27), ZN => n2701);
   U1358 : OAI21_X1 port map( B1 => n2412, B2 => n2701, A => n2392, ZN => n2028
                           );
   U1359 : NOR3_X1 port map( A1 => n2048, A2 => n2409, A3 => n2049, ZN => n2027
                           );
   U1360 : NAND2_X1 port map( A1 => n2025, A2 => DATA2(27), ZN => n2669);
   U1361 : NAND2_X1 port map( A1 => DATA1(27), A2 => n2701, ZN => n2594);
   U1362 : AOI21_X1 port map( B1 => n2669, B2 => n2594, A => n2416, ZN => n2026
                           );
   U1363 : AOI211_X1 port map( C1 => DATA1(27), C2 => n2028, A => n2027, B => 
                           n2026, ZN => n2042);
   U1364 : AOI22_X1 port map( A1 => n2046, A2 => n2198, B1 => n2029, B2 => 
                           n2503, ZN => n2030);
   U1365 : INV_X1 port map( A => n2030, ZN => n2033);
   U1366 : INV_X1 port map( A => n2031, ZN => n2044);
   U1367 : NOR2_X1 port map( A1 => n2032, A2 => n2067, ZN => n2037);
   U1368 : AOI22_X1 port map( A1 => n2396, A2 => n2033, B1 => n2044, B2 => 
                           n2037, ZN => n2041);
   U1369 : INV_X1 port map( A => n2034, ZN => n2039);
   U1370 : INV_X1 port map( A => n2035, ZN => n2038);
   U1371 : OAI22_X1 port map( A1 => n2039, A2 => n2038, B1 => n2037, B2 => 
                           n2036, ZN => n2040);
   U1372 : NAND4_X1 port map( A1 => n2043, A2 => n2042, A3 => n2041, A4 => 
                           n2040, ZN => OUTALU(27));
   U1373 : NOR2_X1 port map( A1 => n2067, A2 => n2044, ZN => n2057);
   U1374 : INV_X1 port map( A => n2057, ZN => n2063);
   U1375 : NOR2_X1 port map( A1 => n2045, A2 => n2069, ZN => n2056);
   U1376 : AND3_X1 port map( A1 => n2046, A2 => n2503, A3 => n2396, ZN => n2055
                           );
   U1377 : INV_X1 port map( A => DATA2(26), ZN => n2702);
   U1378 : OAI22_X1 port map( A1 => n2512, A2 => n2702, B1 => DATA2(26), B2 => 
                           DATA1(26), ZN => n2591);
   U1379 : OAI22_X1 port map( A1 => n2050, A2 => n2049, B1 => n2048, B2 => 
                           n2047, ZN => n2051);
   U1380 : AOI22_X1 port map( A1 => n2688, A2 => n2051, B1 => n2314, B2 => 
                           dataout_mul_26_port, ZN => n2053);
   U1381 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA2(26), B => 
                           DATA1(26), ZN => n2052);
   U1382 : OAI211_X1 port map( C1 => n2591, C2 => n2416, A => n2053, B => n2052
                           , ZN => n2054);
   U1383 : AOI211_X1 port map( C1 => n2056, C2 => n2070, A => n2055, B => n2054
                           , ZN => n2061);
   U1384 : OAI22_X1 port map( A1 => n2059, A2 => n2058, B1 => n2057, B2 => 
                           n2056, ZN => n2060);
   U1385 : OAI211_X1 port map( C1 => n2063, C2 => n2062, A => n2061, B => n2060
                           , ZN => OUTALU(26));
   U1386 : NAND2_X1 port map( A1 => DATA2(25), A2 => n2668, ZN => n2064);
   U1387 : OAI21_X1 port map( B1 => DATA2(25), B2 => n2668, A => n2064, ZN => 
                           n2521_port);
   U1388 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_25_port, B1 => 
                           n2393, B2 => n2521_port, ZN => n2078);
   U1389 : OAI22_X1 port map( A1 => n2080, A2 => n2066, B1 => n2065, B2 => 
                           n2079, ZN => n2074);
   U1390 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n2082);
   U1391 : AOI211_X1 port map( C1 => n2082, C2 => n2071, A => n2068, B => n2067
                           , ZN => n2073);
   U1392 : AOI211_X1 port map( C1 => n2090, C2 => n2071, A => n2070, B => n2069
                           , ZN => n2072);
   U1393 : AOI211_X1 port map( C1 => n2396, C2 => n2074, A => n2073, B => n2072
                           , ZN => n2077);
   U1394 : NAND3_X1 port map( A1 => n2688, A2 => n2121, A3 => n2123, ZN => 
                           n2076);
   U1395 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA2(25), B => 
                           DATA1(25), ZN => n2075);
   U1396 : NAND4_X1 port map( A1 => n2078, A2 => n2077, A3 => n2076, A4 => 
                           n2075, ZN => OUTALU(25));
   U1397 : AOI22_X1 port map( A1 => DATA2_I_24_port, A2 => n2089, B1 => n2367, 
                           B2 => DATA2(24), ZN => n2092);
   U1398 : NOR3_X1 port map( A1 => n2080, A2 => n2079, A3 => n2382, ZN => n2088
                           );
   U1399 : AOI22_X1 port map( A1 => n2449, A2 => n2123, B1 => n2121, B2 => 
                           n2124, ZN => n2086);
   U1400 : INV_X1 port map( A => DATA2(24), ZN => n2704);
   U1401 : OAI22_X1 port map( A1 => n2661, A2 => DATA2(24), B1 => n2704, B2 => 
                           DATA1(24), ZN => n2658);
   U1402 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_24_port, B1 => 
                           n2393, B2 => n2658, ZN => n2085);
   U1403 : INV_X1 port map( A => n2090, ZN => n2081);
   U1404 : NAND3_X1 port map( A1 => n2083, A2 => n2082, A3 => n2081, ZN => 
                           n2084);
   U1405 : OAI211_X1 port map( C1 => n2086, C2 => n2409, A => n2085, B => n2084
                           , ZN => n2087);
   U1406 : AOI211_X1 port map( C1 => n2090, C2 => n2089, A => n2088, B => n2087
                           , ZN => n2091);
   U1407 : OAI221_X1 port map( B1 => n2661, B2 => n2092, C1 => n2661, C2 => 
                           n2392, A => n2091, ZN => OUTALU(24));
   U1408 : NAND2_X1 port map( A1 => DATA2(23), A2 => n2093, ZN => n2664);
   U1409 : INV_X1 port map( A => DATA2(23), ZN => n2705);
   U1410 : NAND2_X1 port map( A1 => DATA1(23), A2 => n2705, ZN => n2587);
   U1411 : AOI21_X1 port map( B1 => n2664, B2 => n2587, A => n2416, ZN => n2097
                           );
   U1412 : AOI222_X1 port map( A1 => n2122, A2 => n2121, B1 => n2124, B2 => 
                           n2449, C1 => n2123, C2 => n2125, ZN => n2095);
   U1413 : AOI21_X1 port map( B1 => n2367, B2 => DATA2(23), A => n2365, ZN => 
                           n2094);
   U1414 : OAI22_X1 port map( A1 => n2095, A2 => n2409, B1 => n2094, B2 => 
                           n2093, ZN => n2096);
   U1415 : AOI211_X1 port map( C1 => n2422, C2 => dataout_mul_23_port, A => 
                           n2097, B => n2096, ZN => n2117);
   U1416 : NOR2_X1 port map( A1 => n3038, A2 => n2098, ZN => n2215);
   U1417 : INV_X1 port map( A => n2149, ZN => n2151);
   U1418 : INV_X1 port map( A => n2152, ZN => n2155);
   U1419 : OAI21_X1 port map( B1 => n2155, B2 => n2164, A => n2102, ZN => n2139
                           );
   U1420 : AOI21_X1 port map( B1 => n2151, B2 => n2139, A => n2103, ZN => n2105
                           );
   U1421 : NAND2_X1 port map( A1 => n2098, A2 => n2696, ZN => n2279);
   U1422 : INV_X1 port map( A => n2279, ZN => n2247);
   U1423 : INV_X1 port map( A => n2234, ZN => n2249);
   U1424 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n2257);
   U1425 : OAI21_X1 port map( B1 => n2257, B2 => n2259, A => n2099, ZN => n2248
                           );
   U1426 : NAND2_X1 port map( A1 => n2249, A2 => n2248, ZN => n2246);
   U1427 : AND2_X1 port map( A1 => n2100, A2 => n2246, ZN => n2214);
   U1428 : OAI21_X1 port map( B1 => n2227, B2 => n2214, A => n2101, ZN => n2153
                           );
   U1429 : INV_X1 port map( A => n2153, ZN => n2154);
   U1430 : OAI21_X1 port map( B1 => n2154, B2 => n2164, A => n2102, ZN => n2138
                           );
   U1431 : AOI21_X1 port map( B1 => n2151, B2 => n2138, A => n2103, ZN => n2104
                           );
   U1432 : AOI22_X1 port map( A1 => n2215, A2 => n2105, B1 => n2247, B2 => 
                           n2104, ZN => n2134);
   U1433 : AOI211_X1 port map( C1 => n2134, C2 => n2137, A => n2108, B => n3038
                           , ZN => n2110);
   U1434 : INV_X1 port map( A => n2215, ZN => n2277);
   U1435 : OAI22_X1 port map( A1 => n2277, A2 => n2105, B1 => n2279, B2 => 
                           n2104, ZN => n2106);
   U1436 : INV_X1 port map( A => n2106, ZN => n2136);
   U1437 : OAI22_X1 port map( A1 => n2136, A2 => n2135, B1 => n3038, B2 => 
                           n2109, ZN => n2107);
   U1438 : AOI22_X1 port map( A1 => n2110, A2 => n2109, B1 => n2108, B2 => 
                           n2107, ZN => n2116);
   U1439 : OAI22_X1 port map( A1 => n2111, A2 => n2375, B1 => n2119, B2 => 
                           n2492, ZN => n2114);
   U1440 : OAI22_X1 port map( A1 => n2141, A2 => n2118, B1 => n2156, B2 => 
                           n2112, ZN => n2113);
   U1441 : OAI21_X1 port map( B1 => n2114, B2 => n2113, A => n2396, ZN => n2115
                           );
   U1442 : NAND3_X1 port map( A1 => n2117, A2 => n2116, A3 => n2115, ZN => 
                           OUTALU(23));
   U1443 : OAI222_X1 port map( A1 => n2375, A2 => n2119, B1 => n2118, B2 => 
                           n2156, C1 => n2492, C2 => n2141, ZN => n2132);
   U1444 : INV_X1 port map( A => DATA2(22), ZN => n2706);
   U1445 : AOI211_X1 port map( C1 => n2392, C2 => n2412, A => n2126, B => n2706
                           , ZN => n2131);
   U1446 : AOI22_X1 port map( A1 => n2449, A2 => n2122, B1 => n2121, B2 => 
                           n2120, ZN => n2129);
   U1447 : AOI22_X1 port map( A1 => n2125, A2 => n2124, B1 => n2183, B2 => 
                           n2123, ZN => n2128);
   U1448 : OAI22_X1 port map( A1 => n2126, A2 => n2706, B1 => DATA2(22), B2 => 
                           DATA1(22), ZN => n2655);
   U1449 : INV_X1 port map( A => n2655, ZN => n2583);
   U1450 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_22_port, B1 => 
                           n2393, B2 => n2583, ZN => n2127);
   U1451 : OAI221_X1 port map( B1 => n2409, B2 => n2129, C1 => n2409, C2 => 
                           n2128, A => n2127, ZN => n2130);
   U1452 : AOI211_X1 port map( C1 => n2396, C2 => n2132, A => n2131, B => n2130
                           , ZN => n2133);
   U1453 : OAI221_X1 port map( B1 => n2137, B2 => n2136, C1 => n2135, C2 => 
                           n2134, A => n2133, ZN => OUTALU(22));
   U1454 : AOI22_X1 port map( A1 => n2215, A2 => n2139, B1 => n2247, B2 => 
                           n2138, ZN => n2150);
   U1455 : OAI22_X1 port map( A1 => n2277, A2 => n2139, B1 => n2279, B2 => 
                           n2138, ZN => n2140);
   U1456 : INV_X1 port map( A => n2140, ZN => n2148);
   U1457 : OAI22_X1 port map( A1 => n2141, A2 => n2375, B1 => n2156, B2 => 
                           n2492, ZN => n2146);
   U1458 : AOI21_X1 port map( B1 => n2367, B2 => DATA2(21), A => n2365, ZN => 
                           n2144);
   U1459 : NAND2_X1 port map( A1 => DATA2(21), A2 => n2652, ZN => n2654);
   U1460 : OAI21_X1 port map( B1 => DATA2(21), B2 => n2652, A => n2654, ZN => 
                           n2524_port);
   U1461 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_21_port, B1 => 
                           n2393, B2 => n2524_port, ZN => n2143);
   U1462 : NAND3_X1 port map( A1 => n2688, A2 => n2397, A3 => n2238, ZN => 
                           n2142);
   U1463 : OAI211_X1 port map( C1 => n2144, C2 => n2652, A => n2143, B => n2142
                           , ZN => n2145);
   U1464 : AOI21_X1 port map( B1 => n2396, B2 => n2146, A => n2145, ZN => n2147
                           );
   U1465 : OAI221_X1 port map( B1 => n2151, B2 => n2150, C1 => n2149, C2 => 
                           n2148, A => n2147, ZN => OUTALU(21));
   U1466 : INV_X1 port map( A => n2164, ZN => n2166);
   U1467 : AOI22_X1 port map( A1 => n2247, A2 => n2153, B1 => n2215, B2 => 
                           n2152, ZN => n2165);
   U1468 : AOI22_X1 port map( A1 => n2155, A2 => n2215, B1 => n2247, B2 => 
                           n2154, ZN => n2163);
   U1469 : INV_X1 port map( A => DATA2(20), ZN => n2708);
   U1470 : OAI21_X1 port map( B1 => n2412, B2 => n2708, A => n2392, ZN => n2161
                           );
   U1471 : NOR3_X1 port map( A1 => n2156, A2 => n2375, A3 => n2382, ZN => n2160
                           );
   U1472 : AOI22_X1 port map( A1 => n2397, A2 => n2236, B1 => n2461, B2 => 
                           n2238, ZN => n2158);
   U1473 : OAI22_X1 port map( A1 => n2653, A2 => DATA2(20), B1 => n2708, B2 => 
                           DATA1(20), ZN => n2648);
   U1474 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_20_port, B1 => 
                           n2393, B2 => n2648, ZN => n2157);
   U1475 : OAI21_X1 port map( B1 => n2158, B2 => n2409, A => n2157, ZN => n2159
                           );
   U1476 : AOI211_X1 port map( C1 => DATA1(20), C2 => n2161, A => n2160, B => 
                           n2159, ZN => n2162);
   U1477 : OAI221_X1 port map( B1 => n2166, B2 => n2165, C1 => n2164, C2 => 
                           n2163, A => n2162, ZN => OUTALU(20));
   U1478 : AOI22_X1 port map( A1 => DATA2(1), A2 => DATA1(1), B1 => n2604, B2 
                           => n2729, ZN => n2513);
   U1479 : AND2_X1 port map( A1 => n2393, A2 => n2513, ZN => n2169);
   U1480 : AOI211_X1 port map( C1 => n2413, C2 => n2206, A => n2167, B => n2415
                           , ZN => n2168);
   U1481 : AOI211_X1 port map( C1 => n2422, C2 => dataout_mul_1_port, A => 
                           n2169, B => n2168, ZN => n2212);
   U1482 : AOI21_X1 port map( B1 => n2396, B2 => n2170, A => n2365, ZN => n2411
                           );
   U1483 : OAI21_X1 port map( B1 => n2729, B2 => n2412, A => n2411, ZN => n2204
                           );
   U1484 : INV_X1 port map( A => n2484, ZN => n2195);
   U1485 : INV_X1 port map( A => n2171, ZN => n2479);
   U1486 : INV_X1 port map( A => n2451, ZN => n2187);
   U1487 : AOI211_X1 port map( C1 => DATA1(5), C2 => n2431, A => n2173, B => 
                           n2172, ZN => n2175);
   U1488 : OAI211_X1 port map( C1 => n2428, C2 => n2604, A => n2175, B => n2174
                           , ZN => n2435);
   U1489 : AOI222_X1 port map( A1 => n2177, A2 => n2434, B1 => n2435, B2 => 
                           n2176, C1 => n2433, C2 => n2436, ZN => n2425);
   U1490 : OAI22_X1 port map( A1 => n2440, A2 => n2425, B1 => n2445, B2 => 
                           n2442, ZN => n2181);
   U1491 : OAI22_X1 port map( A1 => n2444, A2 => n2179, B1 => n2441, B2 => 
                           n2178, ZN => n2180);
   U1492 : AOI211_X1 port map( C1 => n2183, C2 => n2182, A => n2181, B => n2180
                           , ZN => n2424);
   U1493 : OAI22_X1 port map( A1 => n2457, A2 => n2452, B1 => n2424, B2 => 
                           n2454, ZN => n2186);
   U1494 : OAI22_X1 port map( A1 => n2456, A2 => n2184, B1 => n2455, B2 => 
                           n2458, ZN => n2185);
   U1495 : AOI211_X1 port map( C1 => n2461, C2 => n2187, A => n2186, B => n2185
                           , ZN => n2466);
   U1496 : OAI222_X1 port map( A1 => n2465, A2 => n2468, B1 => n2463, B2 => 
                           n2466, C1 => n2188, C2 => n2467, ZN => n2474);
   U1497 : AOI22_X1 port map( A1 => n2345, A2 => n2475, B1 => n2472, B2 => 
                           n2474, ZN => n2191);
   U1498 : AOI22_X1 port map( A1 => n2473, A2 => n2470, B1 => n2476, B2 => 
                           n2189, ZN => n2190);
   U1499 : OAI211_X1 port map( C1 => n2479, C2 => n2230, A => n2191, B => n2190
                           , ZN => n2423);
   U1500 : AOI22_X1 port map( A1 => n2481, A2 => n2423, B1 => n2483, B2 => 
                           n2486, ZN => n2194);
   U1501 : AOI22_X1 port map( A1 => n2487, A2 => n2192, B1 => n2485, B2 => 
                           n2488, ZN => n2193);
   U1502 : OAI211_X1 port map( C1 => n2195, C2 => n2492, A => n2194, B => n2193
                           , ZN => n2497);
   U1503 : AOI222_X1 port map( A1 => n2196, A2 => n2493, B1 => n2494, B2 => 
                           n2498, C1 => n2497, C2 => n2496, ZN => n2511);
   U1504 : INV_X1 port map( A => n2511, ZN => n2197);
   U1505 : AOI22_X1 port map( A1 => n2503, A2 => n2197, B1 => n2505, B2 => 
                           n2506, ZN => n2201);
   U1506 : AOI22_X1 port map( A1 => n2507, A2 => n2199, B1 => n2198, B2 => 
                           n2500, ZN => n2200);
   U1507 : OAI211_X1 port map( C1 => n2203, C2 => n2202, A => n2201, B => n2200
                           , ZN => n2689);
   U1508 : AOI22_X1 port map( A1 => DATA1(1), A2 => n2204, B1 => n2688, B2 => 
                           n2689, ZN => n2211);
   U1509 : NAND3_X1 port map( A1 => n2205, A2 => DATA1(0), A3 => n2396, ZN => 
                           n2210);
   U1510 : OAI221_X1 port map( B1 => n2414, B2 => n2208, C1 => n2207, C2 => 
                           n2206, A => n2420, ZN => n2209);
   U1511 : NAND4_X1 port map( A1 => n2212, A2 => n2211, A3 => n2210, A4 => 
                           n2209, ZN => OUTALU(1));
   U1512 : INV_X1 port map( A => n2227, ZN => n2229);
   U1513 : OAI22_X1 port map( A1 => n2279, A2 => n2214, B1 => n2277, B2 => 
                           n2216, ZN => n2213);
   U1514 : INV_X1 port map( A => n2213, ZN => n2228);
   U1515 : AOI22_X1 port map( A1 => n2216, A2 => n2215, B1 => n2247, B2 => 
                           n2214, ZN => n2226);
   U1516 : OAI22_X1 port map( A1 => n2283, A2 => n2217, B1 => n2231, B2 => 
                           n2254, ZN => n2224);
   U1517 : OAI22_X1 port map( A1 => n2255, A2 => n2230, B1 => n2268, B2 => 
                           n2480, ZN => n2223);
   U1518 : AOI222_X1 port map( A1 => n2237, A2 => n2397, B1 => n2236, B2 => 
                           n2461, C1 => n2238, C2 => n2342, ZN => n2221);
   U1519 : INV_X1 port map( A => DATA2(19), ZN => n2709);
   U1520 : OAI21_X1 port map( B1 => n2412, B2 => n2709, A => n2392, ZN => n2218
                           );
   U1521 : AOI22_X1 port map( A1 => DATA1(19), A2 => n2218, B1 => n2314, B2 => 
                           dataout_mul_19_port, ZN => n2220);
   U1522 : NOR2_X1 port map( A1 => DATA1(19), A2 => n2709, ZN => n2649);
   U1523 : NAND2_X1 port map( A1 => DATA1(19), A2 => n2709, ZN => n2579);
   U1524 : INV_X1 port map( A => n2579, ZN => n2517_port);
   U1525 : OAI21_X1 port map( B1 => n2649, B2 => n2517_port, A => n2393, ZN => 
                           n2219);
   U1526 : OAI211_X1 port map( C1 => n2221, C2 => n2409, A => n2220, B => n2219
                           , ZN => n2222);
   U1527 : AOI221_X1 port map( B1 => n2224, B2 => n2396, C1 => n2223, C2 => 
                           n2396, A => n2222, ZN => n2225);
   U1528 : OAI221_X1 port map( B1 => n2229, B2 => n2228, C1 => n2227, C2 => 
                           n2226, A => n2225, ZN => OUTALU(19));
   U1529 : OAI222_X1 port map( A1 => n2231, A2 => n2283, B1 => n2268, B2 => 
                           n2230, C1 => n2255, C2 => n2254, ZN => n2232);
   U1530 : INV_X1 port map( A => n2232, ZN => n2252);
   U1531 : INV_X1 port map( A => DATA2(18), ZN => n2710);
   U1532 : OAI21_X1 port map( B1 => n2412, B2 => n2710, A => n2392, ZN => n2245
                           );
   U1533 : AOI211_X1 port map( C1 => n2235, C2 => n2234, A => n2233, B => n2277
                           , ZN => n2244);
   U1534 : AOI22_X1 port map( A1 => n2461, A2 => n2237, B1 => n2342, B2 => 
                           n2236, ZN => n2242);
   U1535 : AOI22_X1 port map( A1 => n2397, A2 => n2239, B1 => n2332, B2 => 
                           n2238, ZN => n2241);
   U1536 : INV_X1 port map( A => DATA1(18), ZN => n2537_port);
   U1537 : OAI22_X1 port map( A1 => n2537_port, A2 => n2710, B1 => DATA2(18), 
                           B2 => DATA1(18), ZN => n2645);
   U1538 : INV_X1 port map( A => n2645, ZN => n2576);
   U1539 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_18_port, B1 => 
                           n2393, B2 => n2576, ZN => n2240);
   U1540 : OAI221_X1 port map( B1 => n2409, B2 => n2242, C1 => n2409, C2 => 
                           n2241, A => n2240, ZN => n2243);
   U1541 : AOI211_X1 port map( C1 => DATA1(18), C2 => n2245, A => n2244, B => 
                           n2243, ZN => n2251);
   U1542 : OAI211_X1 port map( C1 => n2249, C2 => n2248, A => n2247, B => n2246
                           , ZN => n2250);
   U1543 : OAI211_X1 port map( C1 => n2252, C2 => n2382, A => n2251, B => n2250
                           , ZN => OUTALU(18));
   U1544 : NAND2_X1 port map( A1 => DATA2(17), A2 => n2253, ZN => n2644);
   U1545 : NOR2_X1 port map( A1 => n2253, A2 => DATA2(17), ZN => n2577);
   U1546 : INV_X1 port map( A => n2577, ZN => n2642);
   U1547 : NAND2_X1 port map( A1 => n2644, A2 => n2642, ZN => n2523_port);
   U1548 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_17_port, B1 => 
                           n2393, B2 => n2523_port, ZN => n2267);
   U1549 : OAI22_X1 port map( A1 => n2283, A2 => n2255, B1 => n2268, B2 => 
                           n2254, ZN => n2263);
   U1550 : NOR2_X1 port map( A1 => n2257, A2 => n2259, ZN => n2256);
   U1551 : AOI211_X1 port map( C1 => n2257, C2 => n2259, A => n2256, B => n2279
                           , ZN => n2262);
   U1552 : AOI211_X1 port map( C1 => n2260, C2 => n2259, A => n2258, B => n2277
                           , ZN => n2261);
   U1553 : AOI211_X1 port map( C1 => n2396, C2 => n2263, A => n2262, B => n2261
                           , ZN => n2266);
   U1554 : NAND3_X1 port map( A1 => n2688, A2 => n2317, A3 => n2269, ZN => 
                           n2265);
   U1555 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA1(17), B => 
                           DATA2(17), ZN => n2264);
   U1556 : NAND4_X1 port map( A1 => n2267, A2 => n2266, A3 => n2265, A4 => 
                           n2264, ZN => OUTALU(17));
   U1557 : INV_X1 port map( A => n2278, ZN => n2280);
   U1558 : INV_X1 port map( A => DATA2(16), ZN => n2712);
   U1559 : OAI21_X1 port map( B1 => n2412, B2 => n2712, A => n2392, ZN => n2275
                           );
   U1560 : NOR3_X1 port map( A1 => n2283, A2 => n2268, A3 => n2382, ZN => n2274
                           );
   U1561 : AOI22_X1 port map( A1 => n2317, A2 => n2270, B1 => n2281, B2 => 
                           n2269, ZN => n2272);
   U1562 : OAI22_X1 port map( A1 => n2643, A2 => DATA2(16), B1 => n2712, B2 => 
                           DATA1(16), ZN => n2638);
   U1563 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_16_port, B1 => 
                           n2393, B2 => n2638, ZN => n2271);
   U1564 : OAI21_X1 port map( B1 => n2272, B2 => n2409, A => n2271, ZN => n2273
                           );
   U1565 : AOI211_X1 port map( C1 => DATA1(16), C2 => n2275, A => n2274, B => 
                           n2273, ZN => n2276);
   U1566 : OAI221_X1 port map( B1 => n2280, B2 => n2279, C1 => n2278, C2 => 
                           n2277, A => n2276, ZN => OUTALU(16));
   U1567 : AOI22_X1 port map( A1 => n2317, A2 => n2282, B1 => n2281, B2 => 
                           n2316, ZN => n2302);
   U1568 : NOR3_X1 port map( A1 => n2283, A2 => n2303, A3 => n2409, ZN => n2295
                           );
   U1569 : INV_X1 port map( A => n2297, ZN => n2299);
   U1570 : INV_X1 port map( A => n2406, ZN => n2284);
   U1571 : AOI21_X1 port map( B1 => n2391, B2 => n2284, A => n2404, ZN => n2285
                           );
   U1572 : INV_X1 port map( A => n2285, ZN => n2387);
   U1573 : NAND2_X1 port map( A1 => n2286, A2 => n2387, ZN => n2370);
   U1574 : INV_X1 port map( A => n2370, ZN => n2288);
   U1575 : OAI21_X1 port map( B1 => n2373, B2 => n2288, A => n2287, ZN => n2352
                           );
   U1576 : NAND2_X1 port map( A1 => n2352, A2 => n2360, ZN => n2351);
   U1577 : AOI21_X1 port map( B1 => n2329, B2 => n2351, A => n2330, ZN => n2308
                           );
   U1578 : NOR2_X1 port map( A1 => n2311, A2 => n2308, ZN => n2304);
   U1579 : OAI21_X1 port map( B1 => n2304, B2 => n2323, A => n2289, ZN => n2290
                           );
   U1580 : XNOR2_X1 port map( A => n2299, B => n2290, ZN => n2293);
   U1581 : INV_X1 port map( A => DATA2(15), ZN => n2713);
   U1582 : NOR2_X1 port map( A1 => DATA1(15), A2 => n2713, ZN => n2639);
   U1583 : NOR2_X1 port map( A1 => DATA2(15), A2 => n2531_port, ZN => n2572);
   U1584 : OAI21_X1 port map( B1 => n2639, B2 => n2572, A => n2393, ZN => n2292
                           );
   U1585 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA2(15), B => 
                           DATA1(15), ZN => n2291);
   U1586 : OAI211_X1 port map( C1 => n2293, C2 => n2307, A => n2292, B => n2291
                           , ZN => n2294);
   U1587 : AOI211_X1 port map( C1 => n2422, C2 => dataout_mul_15_port, A => 
                           n2295, B => n2294, ZN => n2301);
   U1588 : INV_X1 port map( A => n2298, ZN => n2296);
   U1589 : INV_X1 port map( A => n2388, ZN => n2358);
   U1590 : OAI221_X1 port map( B1 => n2299, B2 => n2298, C1 => n2297, C2 => 
                           n2296, A => n2358, ZN => n2300);
   U1591 : OAI211_X1 port map( C1 => n2302, C2 => n2382, A => n2301, B => n2300
                           , ZN => OUTALU(15));
   U1592 : INV_X1 port map( A => n2303, ZN => n2344);
   U1593 : AOI22_X1 port map( A1 => n2473, A2 => n2344, B1 => n2472, B2 => 
                           n2346, ZN => n2325);
   U1594 : OAI22_X1 port map( A1 => n2305, A2 => n2388, B1 => n2304, B2 => 
                           n2307, ZN => n2322);
   U1595 : INV_X1 port map( A => n2306, ZN => n2310);
   U1596 : NOR2_X1 port map( A1 => n2308, A2 => n2307, ZN => n2309);
   U1597 : AOI21_X1 port map( B1 => n2358, B2 => n2310, A => n2309, ZN => n2328
                           );
   U1598 : NOR3_X1 port map( A1 => n2311, A2 => n2328, A3 => n2323, ZN => n2321
                           );
   U1599 : INV_X1 port map( A => DATA2(14), ZN => n2714);
   U1600 : AOI22_X1 port map( A1 => DATA1(14), A2 => n2714, B1 => DATA2(14), B2
                           => n2532_port, ZN => n2635);
   U1601 : OAI21_X1 port map( B1 => n2532_port, B2 => n2412, A => n2392, ZN => 
                           n2315);
   U1602 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_7_14_port, B =>
                           n2312, Z => n2313);
   U1603 : AOI22_X1 port map( A1 => DATA2(14), A2 => n2315, B1 => n2314, B2 => 
                           n2313, ZN => n2319);
   U1604 : NAND3_X1 port map( A1 => n2317, A2 => n2396, A3 => n2316, ZN => 
                           n2318);
   U1605 : OAI211_X1 port map( C1 => n2635, C2 => n2416, A => n2319, B => n2318
                           , ZN => n2320);
   U1606 : AOI211_X1 port map( C1 => n2323, C2 => n2322, A => n2321, B => n2320
                           , ZN => n2324);
   U1607 : OAI21_X1 port map( B1 => n2325, B2 => n2409, A => n2324, ZN => 
                           OUTALU(14));
   U1608 : AOI222_X1 port map( A1 => n2348, A2 => n2472, B1 => n2344, B2 => 
                           n2469, C1 => n2346, C2 => n2473, ZN => n2341);
   U1609 : NOR2_X1 port map( A1 => n2357, A2 => n2388, ZN => n2327);
   U1610 : INV_X1 port map( A => n2351, ZN => n2326);
   U1611 : OAI211_X1 port map( C1 => n2327, C2 => n2405, A => n2326, B => n2330
                           , ZN => n2340);
   U1612 : OAI21_X1 port map( B1 => n2715, B2 => n2412, A => n2392, ZN => n2338
                           );
   U1613 : AOI21_X1 port map( B1 => n2330, B2 => n2329, A => n2328, ZN => n2337
                           );
   U1614 : AOI22_X1 port map( A1 => n2397, A2 => n2331, B1 => n2461, B2 => 
                           n2343, ZN => n2335);
   U1615 : AOI22_X1 port map( A1 => n2342, A2 => n2364, B1 => n2332, B2 => 
                           n2395, ZN => n2334);
   U1616 : NAND2_X1 port map( A1 => DATA2(13), A2 => n2602, ZN => n2634);
   U1617 : OAI21_X1 port map( B1 => DATA2(13), B2 => n2602, A => n2634, ZN => 
                           n2526_port);
   U1618 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_13_port, B1 => 
                           n2393, B2 => n2526_port, ZN => n2333);
   U1619 : OAI221_X1 port map( B1 => n2382, B2 => n2335, C1 => n2382, C2 => 
                           n2334, A => n2333, ZN => n2336);
   U1620 : AOI211_X1 port map( C1 => DATA1(13), C2 => n2338, A => n2337, B => 
                           n2336, ZN => n2339);
   U1621 : OAI211_X1 port map( C1 => n2341, C2 => n2409, A => n2340, B => n2339
                           , ZN => OUTALU(13));
   U1622 : AOI222_X1 port map( A1 => n2343, A2 => n2397, B1 => n2364, B2 => 
                           n2461, C1 => n2395, C2 => n2342, ZN => n2363);
   U1623 : AOI22_X1 port map( A1 => n2469, A2 => n2346, B1 => n2345, B2 => 
                           n2344, ZN => n2350);
   U1624 : AOI22_X1 port map( A1 => n2473, A2 => n2348, B1 => n2472, B2 => 
                           n2347, ZN => n2349);
   U1625 : AOI21_X1 port map( B1 => n2350, B2 => n2349, A => n2409, ZN => n2356
                           );
   U1626 : OAI22_X1 port map( A1 => n2633, A2 => DATA2(12), B1 => n2716, B2 => 
                           DATA1(12), ZN => n2632);
   U1627 : INV_X1 port map( A => n2632, ZN => n2567);
   U1628 : OAI211_X1 port map( C1 => n2360, C2 => n2352, A => n2405, B => n2351
                           , ZN => n2354);
   U1629 : OAI211_X1 port map( C1 => n2365, C2 => n2367, A => DATA1(12), B => 
                           DATA2(12), ZN => n2353);
   U1630 : OAI211_X1 port map( C1 => n2567, C2 => n2416, A => n2354, B => n2353
                           , ZN => n2355);
   U1631 : AOI211_X1 port map( C1 => n2422, C2 => dataout_mul_12_port, A => 
                           n2356, B => n2355, ZN => n2362);
   U1632 : OAI211_X1 port map( C1 => n2360, C2 => n2359, A => n2358, B => n2357
                           , ZN => n2361);
   U1633 : OAI211_X1 port map( C1 => n2363, C2 => n2382, A => n2362, B => n2361
                           , ZN => OUTALU(12));
   U1634 : AOI22_X1 port map( A1 => n2397, A2 => n2364, B1 => n2461, B2 => 
                           n2395, ZN => n2383);
   U1635 : AOI221_X1 port map( B1 => n2367, B2 => DATA1(11), C1 => n2393, C2 =>
                           n2366, A => n2365, ZN => n2368);
   U1636 : NAND2_X1 port map( A1 => DATA1(11), A2 => n2717, ZN => n2566);
   U1637 : OAI22_X1 port map( A1 => n2368, A2 => n2717, B1 => n2416, B2 => 
                           n2566, ZN => n2369);
   U1638 : AOI21_X1 port map( B1 => n2422, B2 => dataout_mul_11_port, A => 
                           n2369, ZN => n2381);
   U1639 : INV_X1 port map( A => n2373, ZN => n2371);
   U1640 : XOR2_X1 port map( A => n2371, B => n2370, Z => n2379);
   U1641 : INV_X1 port map( A => n2374, ZN => n2372);
   U1642 : AOI221_X1 port map( B1 => n2374, B2 => n2373, C1 => n2372, C2 => 
                           n2371, A => n2388, ZN => n2378);
   U1643 : NOR3_X1 port map( A1 => n2376, A2 => n2409, A3 => n2375, ZN => n2377
                           );
   U1644 : AOI211_X1 port map( C1 => n2405, C2 => n2379, A => n2378, B => n2377
                           , ZN => n2380);
   U1645 : OAI211_X1 port map( C1 => n2383, C2 => n2382, A => n2381, B => n2380
                           , ZN => OUTALU(11));
   U1646 : AOI22_X1 port map( A1 => n2386, A2 => n2385, B1 => n2481, B2 => 
                           n2384, ZN => n2410);
   U1647 : NAND2_X1 port map( A1 => n2405, A2 => n2387, ZN => n2390);
   U1648 : OR2_X1 port map( A1 => n2389, A2 => n2388, ZN => n2401);
   U1649 : AOI22_X1 port map( A1 => n2404, A2 => n2391, B1 => n2390, B2 => 
                           n2401, ZN => n2403);
   U1650 : OAI21_X1 port map( B1 => n2718, B2 => n2412, A => n2392, ZN => n2394
                           );
   U1651 : AOI22_X1 port map( A1 => DATA1(10), A2 => DATA2(10), B1 => n2718, B2
                           => n2516, ZN => n2625);
   U1652 : AOI22_X1 port map( A1 => DATA1(10), A2 => n2394, B1 => n2393, B2 => 
                           n2625, ZN => n2399);
   U1653 : NAND3_X1 port map( A1 => n2397, A2 => n2396, A3 => n2395, ZN => 
                           n2398);
   U1654 : OAI211_X1 port map( C1 => n2401, C2 => n2400, A => n2399, B => n2398
                           , ZN => n2402);
   U1655 : AOI211_X1 port map( C1 => n2422, C2 => dataout_mul_10_port, A => 
                           n2403, B => n2402, ZN => n2408);
   U1656 : NAND3_X1 port map( A1 => n2406, A2 => n2405, A3 => n2404, ZN => 
                           n2407);
   U1657 : OAI211_X1 port map( C1 => n2410, C2 => n2409, A => n2408, B => n2407
                           , ZN => OUTALU(10));
   U1658 : OAI21_X1 port map( B1 => n2730, B2 => n2412, A => n2411, ZN => n2419
                           );
   U1659 : OAI22_X1 port map( A1 => n2730, A2 => DATA1(0), B1 => n2603, B2 => 
                           DATA2(0), ZN => n2514);
   U1660 : INV_X1 port map( A => n2514, ZN => n2417);
   U1661 : NOR2_X1 port map( A1 => n2414, A2 => n2413, ZN => n2421);
   U1662 : OAI22_X1 port map( A1 => n2417, A2 => n2416, B1 => n2421, B2 => 
                           n2415, ZN => n2418);
   U1663 : AOI21_X1 port map( B1 => DATA1(0), B2 => n2419, A => n2418, ZN => 
                           n2694);
   U1664 : AOI22_X1 port map( A1 => n2422, A2 => dataout_mul_0_port, B1 => 
                           n2421, B2 => n2420, ZN => n2693);
   U1665 : INV_X1 port map( A => n2423, ZN => n2491);
   U1666 : INV_X1 port map( A => n2424, ZN => n2462);
   U1667 : INV_X1 port map( A => n2425, ZN => n2450);
   U1668 : OAI211_X1 port map( C1 => n2428, C2 => n2603, A => n2427, B => n2426
                           , ZN => n2429);
   U1669 : AOI211_X1 port map( C1 => DATA1(4), C2 => n2431, A => n2430, B => 
                           n2429, ZN => n2432);
   U1670 : INV_X1 port map( A => n2432, ZN => n2437);
   U1671 : AOI222_X1 port map( A1 => n2438, A2 => n2437, B1 => n2436, B2 => 
                           n2435, C1 => n2434, C2 => n2433, ZN => n2439);
   U1672 : OAI22_X1 port map( A1 => n2442, A2 => n2441, B1 => n2440, B2 => 
                           n2439, ZN => n2448);
   U1673 : OAI22_X1 port map( A1 => n2446, A2 => n2445, B1 => n2444, B2 => 
                           n2443, ZN => n2447);
   U1674 : AOI211_X1 port map( C1 => n2450, C2 => n2449, A => n2448, B => n2447
                           , ZN => n2453);
   U1675 : OAI22_X1 port map( A1 => n2454, A2 => n2453, B1 => n2452, B2 => 
                           n2451, ZN => n2460);
   U1676 : OAI22_X1 port map( A1 => n2458, A2 => n2457, B1 => n2456, B2 => 
                           n2455, ZN => n2459);
   U1677 : AOI211_X1 port map( C1 => n2462, C2 => n2461, A => n2460, B => n2459
                           , ZN => n2464);
   U1678 : OAI222_X1 port map( A1 => n2468, A2 => n2467, B1 => n2466, B2 => 
                           n2465, C1 => n2464, C2 => n2463, ZN => n2471);
   U1679 : AOI22_X1 port map( A1 => n2472, A2 => n2471, B1 => n2470, B2 => 
                           n2469, ZN => n2478);
   U1680 : AOI22_X1 port map( A1 => n2476, A2 => n2475, B1 => n2474, B2 => 
                           n2473, ZN => n2477);
   U1681 : OAI211_X1 port map( C1 => n2480, C2 => n2479, A => n2478, B => n2477
                           , ZN => n2482);
   U1682 : AOI22_X1 port map( A1 => n2484, A2 => n2483, B1 => n2482, B2 => 
                           n2481, ZN => n2490);
   U1683 : AOI22_X1 port map( A1 => n2488, A2 => n2487, B1 => n2486, B2 => 
                           n2485, ZN => n2489);
   U1684 : OAI211_X1 port map( C1 => n2492, C2 => n2491, A => n2490, B => n2489
                           , ZN => n2495);
   U1685 : AOI222_X1 port map( A1 => n2498, A2 => n2497, B1 => n2496, B2 => 
                           n2495, C1 => n2494, C2 => n2493, ZN => n2499);
   U1686 : INV_X1 port map( A => n2499, ZN => n2502);
   U1687 : AOI22_X1 port map( A1 => n2503, A2 => n2502, B1 => n2501, B2 => 
                           n2500, ZN => n2509);
   U1688 : AOI22_X1 port map( A1 => n2507, A2 => n2506, B1 => n2505, B2 => 
                           n2504, ZN => n2508);
   U1689 : OAI211_X1 port map( C1 => n2511, C2 => n2510, A => n2509, B => n2508
                           , ZN => n2687);
   U1690 : OAI21_X1 port map( B1 => DATA2(26), B2 => n2512, A => n2594, ZN => 
                           n2671);
   U1691 : AOI22_X1 port map( A1 => n2599, A2 => DATA2(31), B1 => n2698, B2 => 
                           DATA1(30), ZN => n2681);
   U1692 : INV_X1 port map( A => n2681, ZN => n2515);
   U1693 : NOR4_X1 port map( A1 => n2671, A2 => n2515, A3 => n2514, A4 => n2513
                           , ZN => n2530_port);
   U1694 : OAI21_X1 port map( B1 => DATA2(10), B2 => n2516, A => n2566, ZN => 
                           n2629);
   U1695 : INV_X1 port map( A => n2629, ZN => n2518_port);
   U1696 : AOI22_X1 port map( A1 => n2714, A2 => DATA1(14), B1 => n2713, B2 => 
                           DATA1(15), ZN => n2641);
   U1697 : AOI21_X1 port map( B1 => n2710, B2 => DATA1(18), A => n2517_port, ZN
                           => n2651);
   U1698 : AOI22_X1 port map( A1 => n2706, A2 => DATA1(22), B1 => n2705, B2 => 
                           DATA1(23), ZN => n2660);
   U1699 : AND4_X1 port map( A1 => n2518_port, A2 => n2641, A3 => n2651, A4 => 
                           n2660, ZN => n2529_port);
   U1700 : NOR4_X1 port map( A1 => n2522_port, A2 => n2521_port, A3 => 
                           n2520_port, A4 => n2519_port, ZN => n2528_port);
   U1701 : NOR4_X1 port map( A1 => n2526_port, A2 => n2525_port, A3 => 
                           n2524_port, A4 => n2523_port, ZN => n2527_port);
   U1702 : NAND4_X1 port map( A1 => n2530_port, A2 => n2529_port, A3 => 
                           n2528_port, A4 => n2527_port, ZN => n2544_port);
   U1703 : OAI22_X1 port map( A1 => n2718, A2 => DATA1(10), B1 => n2717, B2 => 
                           DATA1(11), ZN => n2568);
   U1704 : AOI22_X1 port map( A1 => DATA2(14), A2 => n2532_port, B1 => 
                           DATA2(15), B2 => n2531_port, ZN => n2574);
   U1705 : INV_X1 port map( A => n2574, ZN => n2533_port);
   U1706 : OR4_X1 port map( A1 => n2568, A2 => n2632, A3 => n2533_port, A4 => 
                           n2638, ZN => n2542_port);
   U1707 : AOI22_X1 port map( A1 => DATA2(6), A2 => n2534_port, B1 => DATA2(7),
                           B2 => n2620, ZN => n2560);
   U1708 : INV_X1 port map( A => n2557, ZN => n2624);
   U1709 : NAND4_X1 port map( A1 => n2606, A2 => n2550, A3 => n2560, A4 => 
                           n2624, ZN => n2541_port);
   U1710 : OAI21_X1 port map( B1 => n2702, B2 => DATA1(26), A => n2669, ZN => 
                           n2595);
   U1711 : INV_X1 port map( A => n2595, ZN => n2536_port);
   U1712 : AOI21_X1 port map( B1 => DATA2(30), B2 => n2535_port, A => n2679, ZN
                           => n2601);
   U1713 : AOI21_X1 port map( B1 => DATA1(6), B2 => n2724, A => n2558, ZN => 
                           n2622);
   U1714 : NAND4_X1 port map( A1 => n2536_port, A2 => n2670, A3 => n2601, A4 =>
                           n2622, ZN => n2540_port);
   U1715 : AOI21_X1 port map( B1 => DATA2(18), B2 => n2537_port, A => n2649, ZN
                           => n2538_port);
   U1716 : INV_X1 port map( A => n2538_port, ZN => n2581);
   U1717 : OAI22_X1 port map( A1 => n2705, A2 => DATA1(23), B1 => n2706, B2 => 
                           DATA1(22), ZN => n2589);
   U1718 : OR4_X1 port map( A1 => n2581, A2 => n2648, A3 => n2589, A4 => n2658,
                           ZN => n2539_port);
   U1719 : OR4_X1 port map( A1 => n2542_port, A2 => n2541_port, A3 => 
                           n2540_port, A4 => n2539_port, ZN => n2543_port);
   U1720 : OAI21_X1 port map( B1 => n2544_port, B2 => n2543_port, A => n2695, 
                           ZN => n2546_port);
   U1721 : INV_X1 port map( A => FUNC(0), ZN => n2545_port);
   U1722 : AOI211_X1 port map( C1 => FUNC(2), C2 => n2546_port, A => FUNC(1), B
                           => n2545_port, ZN => n2686);
   U1723 : AOI22_X1 port map( A1 => DATA2(25), A2 => n2668, B1 => DATA2(24), B2
                           => n2661, ZN => n2593);
   U1724 : AOI22_X1 port map( A1 => DATA2(21), A2 => n2652, B1 => DATA2(20), B2
                           => n2653, ZN => n2586);
   U1725 : OAI21_X1 port map( B1 => DATA2(1), B2 => n2604, A => DATA2(0), ZN =>
                           n2547_port);
   U1726 : OAI22_X1 port map( A1 => DATA1(0), A2 => n2547_port, B1 => DATA1(1),
                           B2 => n2729, ZN => n2548_port);
   U1727 : AOI22_X1 port map( A1 => DATA2(2), A2 => n2611, B1 => n2606, B2 => 
                           n2548_port, ZN => n2549);
   U1728 : INV_X1 port map( A => n2549, ZN => n2551);
   U1729 : NOR2_X1 port map( A1 => n2727, A2 => DATA1(3), ZN => n2615);
   U1730 : NAND2_X1 port map( A1 => n2727, A2 => DATA1(3), ZN => n2609);
   U1731 : OAI211_X1 port map( C1 => n2551, C2 => n2615, A => n2609, B => n2550
                           , ZN => n2552);
   U1732 : INV_X1 port map( A => n2552, ZN => n2556);
   U1733 : NAND2_X1 port map( A1 => DATA2(5), A2 => n2553, ZN => n2616);
   U1734 : OAI21_X1 port map( B1 => DATA1(4), B2 => n2726, A => n2616, ZN => 
                           n2555);
   U1735 : NOR2_X1 port map( A1 => n2553, A2 => DATA2(5), ZN => n2619);
   U1736 : INV_X1 port map( A => n2619, ZN => n2554);
   U1737 : OAI211_X1 port map( C1 => n2556, C2 => n2555, A => n2617, B => n2554
                           , ZN => n2559);
   U1738 : AOI211_X1 port map( C1 => n2560, C2 => n2559, A => n2558, B => n2557
                           , ZN => n2561);
   U1739 : AOI21_X1 port map( B1 => DATA2(8), B2 => n2562, A => n2561, ZN => 
                           n2565);
   U1740 : INV_X1 port map( A => n2627, ZN => n2563);
   U1741 : AOI211_X1 port map( C1 => n2565, C2 => n2564, A => n2563, B => n2625
                           , ZN => n2569);
   U1742 : OAI211_X1 port map( C1 => n2569, C2 => n2568, A => n2567, B => n2566
                           , ZN => n2570);
   U1743 : OAI211_X1 port map( C1 => DATA1(12), C2 => n2716, A => n2570, B => 
                           n2634, ZN => n2571);
   U1744 : OAI211_X1 port map( C1 => DATA2(13), C2 => n2602, A => n2635, B => 
                           n2571, ZN => n2573);
   U1745 : AOI211_X1 port map( C1 => n2574, C2 => n2573, A => n2572, B => n2638
                           , ZN => n2575);
   U1746 : AOI21_X1 port map( B1 => DATA2(16), B2 => n2643, A => n2575, ZN => 
                           n2578);
   U1747 : AOI211_X1 port map( C1 => n2578, C2 => n2644, A => n2577, B => n2576
                           , ZN => n2582);
   U1748 : INV_X1 port map( A => n2648, ZN => n2580);
   U1749 : OAI211_X1 port map( C1 => n2582, C2 => n2581, A => n2580, B => n2579
                           , ZN => n2585);
   U1750 : NOR2_X1 port map( A1 => DATA2(21), A2 => n2652, ZN => n2584);
   U1751 : AOI211_X1 port map( C1 => n2586, C2 => n2585, A => n2584, B => n2583
                           , ZN => n2590);
   U1752 : INV_X1 port map( A => n2658, ZN => n2588);
   U1753 : OAI211_X1 port map( C1 => n2590, C2 => n2589, A => n2588, B => n2587
                           , ZN => n2592);
   U1754 : NOR2_X1 port map( A1 => DATA2(25), A2 => n2668, ZN => n2663);
   U1755 : INV_X1 port map( A => n2591, ZN => n2666);
   U1756 : AOI211_X1 port map( C1 => n2593, C2 => n2592, A => n2663, B => n2666
                           , ZN => n2596);
   U1757 : OAI211_X1 port map( C1 => n2596, C2 => n2595, A => n2670, B => n2594
                           , ZN => n2597);
   U1758 : OAI211_X1 port map( C1 => DATA1(28), C2 => n2700, A => n2597, B => 
                           n2677, ZN => n2598);
   U1759 : NAND3_X1 port map( A1 => n2678, A2 => n2674, A3 => n2598, ZN => 
                           n2600);
   U1760 : AOI22_X1 port map( A1 => n2601, A2 => n2600, B1 => DATA2(31), B2 => 
                           n2599, ZN => n2684);
   U1761 : NOR2_X1 port map( A1 => DATA2(13), A2 => n2602, ZN => n2637);
   U1762 : NOR2_X1 port map( A1 => DATA2(0), A2 => n2603, ZN => n2608);
   U1763 : NOR2_X1 port map( A1 => DATA2(1), A2 => n2604, ZN => n2607);
   U1764 : NAND2_X1 port map( A1 => DATA2(1), A2 => n2604, ZN => n2605);
   U1765 : OAI211_X1 port map( C1 => n2608, C2 => n2607, A => n2606, B => n2605
                           , ZN => n2610);
   U1766 : OAI211_X1 port map( C1 => DATA2(2), C2 => n2611, A => n2610, B => 
                           n2609, ZN => n2612);
   U1767 : OAI21_X1 port map( B1 => DATA1(4), B2 => n2726, A => n2612, ZN => 
                           n2614);
   U1768 : OAI22_X1 port map( A1 => n2615, A2 => n2614, B1 => DATA2(4), B2 => 
                           n2613, ZN => n2618);
   U1769 : OAI211_X1 port map( C1 => n2619, C2 => n2618, A => n2617, B => n2616
                           , ZN => n2621);
   U1770 : AOI22_X1 port map( A1 => n2622, A2 => n2621, B1 => DATA2(7), B2 => 
                           n2620, ZN => n2623);
   U1771 : AOI22_X1 port map( A1 => DATA1(8), A2 => n2720, B1 => n2624, B2 => 
                           n2623, ZN => n2628);
   U1772 : AOI211_X1 port map( C1 => n2628, C2 => n2627, A => n2626, B => n2625
                           , ZN => n2630);
   U1773 : OAI22_X1 port map( A1 => DATA1(11), A2 => n2717, B1 => n2630, B2 => 
                           n2629, ZN => n2631);
   U1774 : OAI22_X1 port map( A1 => DATA2(12), A2 => n2633, B1 => n2632, B2 => 
                           n2631, ZN => n2636);
   U1775 : OAI211_X1 port map( C1 => n2637, C2 => n2636, A => n2635, B => n2634
                           , ZN => n2640);
   U1776 : AOI211_X1 port map( C1 => n2641, C2 => n2640, A => n2639, B => n2638
                           , ZN => n2647);
   U1777 : OAI21_X1 port map( B1 => DATA2(16), B2 => n2643, A => n2642, ZN => 
                           n2646);
   U1778 : OAI211_X1 port map( C1 => n2647, C2 => n2646, A => n2645, B => n2644
                           , ZN => n2650);
   U1779 : AOI211_X1 port map( C1 => n2651, C2 => n2650, A => n2649, B => n2648
                           , ZN => n2657);
   U1780 : OAI22_X1 port map( A1 => DATA2(20), A2 => n2653, B1 => DATA2(21), B2
                           => n2652, ZN => n2656);
   U1781 : OAI211_X1 port map( C1 => n2657, C2 => n2656, A => n2655, B => n2654
                           , ZN => n2659);
   U1782 : AOI21_X1 port map( B1 => n2660, B2 => n2659, A => n2658, ZN => n2665
                           );
   U1783 : NOR2_X1 port map( A1 => DATA2(24), A2 => n2661, ZN => n2662);
   U1784 : AOI211_X1 port map( C1 => n2665, C2 => n2664, A => n2663, B => n2662
                           , ZN => n2667);
   U1785 : AOI211_X1 port map( C1 => DATA2(25), C2 => n2668, A => n2667, B => 
                           n2666, ZN => n2672);
   U1786 : OAI211_X1 port map( C1 => n2672, C2 => n2671, A => n2670, B => n2669
                           , ZN => n2673);
   U1787 : OAI211_X1 port map( C1 => DATA2(28), C2 => n2675, A => n2674, B => 
                           n2673, ZN => n2676);
   U1788 : NAND3_X1 port map( A1 => n2678, A2 => n2677, A3 => n2676, ZN => 
                           n2680);
   U1789 : AOI21_X1 port map( B1 => n2681, B2 => n2680, A => n2679, ZN => n2683
                           );
   U1790 : OAI221_X1 port map( B1 => FUNC(3), B2 => n2684, C1 => n2695, C2 => 
                           n2683, A => n2682, ZN => n2685);
   U1791 : AOI22_X1 port map( A1 => n2688, A2 => n2687, B1 => n2686, B2 => 
                           n2685, ZN => n2692);
   U1792 : NAND3_X1 port map( A1 => n2690, A2 => FUNC(3), A3 => n2689, ZN => 
                           n2691);
   U1793 : NAND4_X1 port map( A1 => n2694, A2 => n2693, A3 => n2692, A4 => 
                           n2691, ZN => OUTALU(0));
   U1794 : NAND2_X1 port map( A1 => n2696, A2 => n2695, ZN => n2732);
   U1795 : CLKBUF_X1 port map( A => n2732, Z => n2722);
   U1796 : NAND2_X1 port map( A1 => FUNC(3), A2 => n2696, ZN => n2731);
   U1797 : INV_X1 port map( A => DATA2(31), ZN => n2697);
   U1798 : AOI22_X1 port map( A1 => DATA2(31), A2 => n2722, B1 => n2721, B2 => 
                           n2697, ZN => N2548);
   U1799 : AOI22_X1 port map( A1 => DATA2(30), A2 => n2732, B1 => n2731, B2 => 
                           n2698, ZN => N2547);
   U1800 : AOI22_X1 port map( A1 => DATA2(29), A2 => n2722, B1 => n2721, B2 => 
                           n2699, ZN => N2546);
   U1801 : AOI22_X1 port map( A1 => DATA2(28), A2 => n2732, B1 => n2731, B2 => 
                           n2700, ZN => N2545);
   U1802 : AOI22_X1 port map( A1 => DATA2(27), A2 => n2722, B1 => n2721, B2 => 
                           n2701, ZN => N2544);
   U1803 : AOI22_X1 port map( A1 => DATA2(26), A2 => n2732, B1 => n2731, B2 => 
                           n2702, ZN => N2543);
   U1804 : INV_X1 port map( A => DATA2(25), ZN => n2703);
   U1805 : AOI22_X1 port map( A1 => DATA2(25), A2 => n2722, B1 => n2721, B2 => 
                           n2703, ZN => N2542);
   U1806 : AOI22_X1 port map( A1 => DATA2(24), A2 => n2732, B1 => n2731, B2 => 
                           n2704, ZN => N2541);
   U1807 : AOI22_X1 port map( A1 => DATA2(23), A2 => n2722, B1 => n2721, B2 => 
                           n2705, ZN => N2540);
   U1808 : AOI22_X1 port map( A1 => DATA2(22), A2 => n2732, B1 => n2731, B2 => 
                           n2706, ZN => N2539);
   U1809 : INV_X1 port map( A => DATA2(21), ZN => n2707);
   U1810 : AOI22_X1 port map( A1 => DATA2(21), A2 => n2732, B1 => n2731, B2 => 
                           n2707, ZN => N2538);
   U1811 : AOI22_X1 port map( A1 => DATA2(20), A2 => n2732, B1 => n2731, B2 => 
                           n2708, ZN => N2537);
   U1812 : AOI22_X1 port map( A1 => DATA2(19), A2 => n2722, B1 => n2721, B2 => 
                           n2709, ZN => N2536);
   U1813 : AOI22_X1 port map( A1 => DATA2(18), A2 => n2722, B1 => n2721, B2 => 
                           n2710, ZN => N2535);
   U1814 : INV_X1 port map( A => DATA2(17), ZN => n2711);
   U1815 : AOI22_X1 port map( A1 => DATA2(17), A2 => n2722, B1 => n2721, B2 => 
                           n2711, ZN => N2534);
   U1816 : AOI22_X1 port map( A1 => DATA2(16), A2 => n2722, B1 => n2721, B2 => 
                           n2712, ZN => N2533);
   U1817 : AOI22_X1 port map( A1 => DATA2(15), A2 => n2722, B1 => n2721, B2 => 
                           n2713, ZN => N2532);
   U1818 : AOI22_X1 port map( A1 => DATA2(14), A2 => n2722, B1 => n2721, B2 => 
                           n2714, ZN => N2531);
   U1819 : AOI22_X1 port map( A1 => DATA2(13), A2 => n2722, B1 => n2721, B2 => 
                           n2715, ZN => N2530);
   U1820 : AOI22_X1 port map( A1 => DATA2(12), A2 => n2722, B1 => n2721, B2 => 
                           n2716, ZN => N2529);
   U1821 : AOI22_X1 port map( A1 => DATA2(11), A2 => n2722, B1 => n2721, B2 => 
                           n2717, ZN => N2528);
   U1822 : AOI22_X1 port map( A1 => DATA2(10), A2 => n2722, B1 => n2721, B2 => 
                           n2718, ZN => N2527);
   U1823 : AOI22_X1 port map( A1 => DATA2(9), A2 => n2722, B1 => n2721, B2 => 
                           n2719, ZN => N2526);
   U1824 : AOI22_X1 port map( A1 => DATA2(8), A2 => n2722, B1 => n2721, B2 => 
                           n2720, ZN => N2525);
   U1825 : INV_X1 port map( A => DATA2(7), ZN => n2723);
   U1826 : AOI22_X1 port map( A1 => DATA2(7), A2 => n2732, B1 => n2731, B2 => 
                           n2723, ZN => N2524);
   U1827 : AOI22_X1 port map( A1 => DATA2(6), A2 => n2732, B1 => n2731, B2 => 
                           n2724, ZN => N2523);
   U1828 : AOI22_X1 port map( A1 => DATA2(5), A2 => n2732, B1 => n2731, B2 => 
                           n2725, ZN => N2522);
   U1829 : AOI22_X1 port map( A1 => DATA2(4), A2 => n2732, B1 => n2731, B2 => 
                           n2726, ZN => N2521);
   U1830 : AOI22_X1 port map( A1 => DATA2(3), A2 => n2732, B1 => n2731, B2 => 
                           n2727, ZN => N2520);
   U1831 : AOI22_X1 port map( A1 => DATA2(2), A2 => n2732, B1 => n2731, B2 => 
                           n2728, ZN => N2519);
   U1832 : AOI22_X1 port map( A1 => DATA2(1), A2 => n2732, B1 => n2731, B2 => 
                           n2729, ZN => N2518);
   U1833 : AOI22_X1 port map( A1 => DATA2(0), A2 => n2732, B1 => n2731, B2 => 
                           n2730, ZN => N2517);
   U1834 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           A2 => n2733, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1835 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN
                           => n2735);
   U1836 : NAND2_X1 port map( A1 => data2_mul_3_port, A2 => n2735, ZN => n2770)
                           ;
   U1837 : INV_X1 port map( A => data2_mul_3_port, ZN => n2768);
   U1838 : NAND3_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, 
                           A3 => n2768, ZN => n2767);
   U1839 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2769, B1 => data1_mul_1_port, B2 => n2763, ZN
                           => n2736);
   U1840 : OAI221_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           B2 => n2770, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           C2 => n2767, A => n2736, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1841 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           n2763, B2 => data1_mul_2_port, ZN => n2738);
   U1842 : INV_X1 port map( A => n2770, ZN => n2764);
   U1843 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2764, ZN => n2737);
   U1844 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, 
                           C2 => n2767, A => n2738, B => n2737, ZN => 
                           boothmul_pipelined_i_mux_out_1_4_port);
   U1845 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n2763, B2 => data1_mul_3_port, ZN => n2740);
   U1846 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, ZN => 
                           n2739);
   U1847 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, 
                           C2 => n2767, A => n2740, B => n2739, ZN => 
                           boothmul_pipelined_i_mux_out_1_5_port);
   U1848 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n2763, B2 => data1_mul_4_port, ZN => n2742);
   U1849 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n2741);
   U1850 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, 
                           C2 => n2767, A => n2742, B => n2741, ZN => 
                           boothmul_pipelined_i_mux_out_1_6_port);
   U1851 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n2763, B2 => data1_mul_5_port, ZN => n2744);
   U1852 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n2743);
   U1853 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, 
                           C2 => n2767, A => n2744, B => n2743, ZN => 
                           boothmul_pipelined_i_mux_out_1_7_port);
   U1854 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n2763, B2 => data1_mul_6_port, ZN => n2746);
   U1855 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n2745);
   U1856 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, 
                           C2 => n2767, A => n2746, B => n2745, ZN => 
                           boothmul_pipelined_i_mux_out_1_8_port);
   U1857 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n2763, B2 => data1_mul_7_port, ZN => n2748);
   U1858 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n2747);
   U1859 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, 
                           C2 => n2767, A => n2748, B => n2747, ZN => 
                           boothmul_pipelined_i_mux_out_1_9_port);
   U1860 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n2763, B2 => data1_mul_8_port, ZN => n2750);
   U1861 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n2749);
   U1862 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, 
                           C2 => n2767, A => n2750, B => n2749, ZN => 
                           boothmul_pipelined_i_mux_out_1_10_port);
   U1863 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n2763, B2 => data1_mul_9_port, ZN => n2752);
   U1864 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n2751);
   U1865 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, 
                           C2 => n2767, A => n2752, B => n2751, ZN => 
                           boothmul_pipelined_i_mux_out_1_11_port);
   U1866 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n2763, B2 => data1_mul_10_port, ZN => n2754);
   U1867 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n2753);
   U1868 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, 
                           C2 => n2767, A => n2754, B => n2753, ZN => 
                           boothmul_pipelined_i_mux_out_1_12_port);
   U1869 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n2763, B2 => data1_mul_11_port, ZN => n2756);
   U1870 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n2755);
   U1871 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, 
                           C2 => n2767, A => n2756, B => n2755, ZN => 
                           boothmul_pipelined_i_mux_out_1_13_port);
   U1872 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n2763, B2 => data1_mul_12_port, ZN => n2758);
   U1873 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n2757);
   U1874 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, 
                           C2 => n2767, A => n2758, B => n2757, ZN => 
                           boothmul_pipelined_i_mux_out_1_14_port);
   U1875 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n2763, B2 => data1_mul_13_port, ZN => n2760);
   U1876 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n2759);
   U1877 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, 
                           C2 => n2767, A => n2760, B => n2759, ZN => 
                           boothmul_pipelined_i_mux_out_1_15_port);
   U1878 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n2763, B2 => data1_mul_14_port, ZN => n2762);
   U1879 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n2761);
   U1880 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, 
                           C2 => n2767, A => n2762, B => n2761, ZN => 
                           boothmul_pipelined_i_mux_out_1_16_port);
   U1881 : AOI22_X1 port map( A1 => n2769, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n2763, B2 => data1_mul_15_port, ZN => n2766);
   U1882 : NAND2_X1 port map( A1 => n2764, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n2765);
   U1883 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, 
                           C2 => n2767, A => n2766, B => n2765, ZN => 
                           boothmul_pipelined_i_mux_out_1_17_port);
   U1884 : OAI21_X1 port map( B1 => data2_mul_1_port, B2 => data2_mul_2_port, A
                           => n2768, ZN => n2772);
   U1885 : INV_X1 port map( A => n2769, ZN => n2771);
   U1886 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_119_port, ZN 
                           => n2809);
   U1887 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN 
                           => n2811);
   U1888 : OAI222_X1 port map( A1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           A2 => n2772, B1 => n2771, B2 => n2809, C1 => n2770, 
                           C2 => n2811, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1889 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n2774);
   U1890 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n2774, ZN => n2812);
   U1891 : NAND3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           A3 => n3025, ZN => n2806);
   U1892 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2807, B1 => data1_mul_1_port, B2 => n2802, ZN
                           => n2775);
   U1893 : OAI221_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           B2 => n2812, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           C2 => n2806, A => n2775, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1894 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B2 => 
                           n2807, ZN => n2777);
   U1895 : INV_X1 port map( A => n2812, ZN => n2803);
   U1896 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2803, ZN => n2776);
   U1897 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, A 
                           => n2777, B => n2776, ZN => 
                           boothmul_pipelined_i_mux_out_2_6_port);
   U1898 : AOI22_X1 port map( A1 => data1_mul_3_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n2807, ZN => n2779);
   U1899 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n2803, ZN => n2778);
   U1900 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, A 
                           => n2779, B => n2778, ZN => 
                           boothmul_pipelined_i_mux_out_2_7_port);
   U1901 : AOI22_X1 port map( A1 => data1_mul_4_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n2807, ZN => n2781);
   U1902 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n2803, ZN => n2780);
   U1903 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, A 
                           => n2781, B => n2780, ZN => 
                           boothmul_pipelined_i_mux_out_2_8_port);
   U1904 : AOI22_X1 port map( A1 => data1_mul_5_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n2807, ZN => n2783);
   U1905 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n2803, ZN => n2782);
   U1906 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, A 
                           => n2783, B => n2782, ZN => 
                           boothmul_pipelined_i_mux_out_2_9_port);
   U1907 : AOI22_X1 port map( A1 => data1_mul_6_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n2807, ZN => n2785);
   U1908 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n2803, ZN => n2784);
   U1909 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, A 
                           => n2785, B => n2784, ZN => 
                           boothmul_pipelined_i_mux_out_2_10_port);
   U1910 : AOI22_X1 port map( A1 => data1_mul_7_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n2807, ZN => n2787);
   U1911 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n2803, ZN => n2786);
   U1912 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, A 
                           => n2787, B => n2786, ZN => 
                           boothmul_pipelined_i_mux_out_2_11_port);
   U1913 : AOI22_X1 port map( A1 => data1_mul_8_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n2807, ZN => n2789);
   U1914 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n2803, ZN => n2788);
   U1915 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, A 
                           => n2789, B => n2788, ZN => 
                           boothmul_pipelined_i_mux_out_2_12_port);
   U1916 : AOI22_X1 port map( A1 => data1_mul_9_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n2807, ZN => n2791);
   U1917 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n2803, ZN => n2790);
   U1918 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, A 
                           => n2791, B => n2790, ZN => 
                           boothmul_pipelined_i_mux_out_2_13_port);
   U1919 : AOI22_X1 port map( A1 => data1_mul_10_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n2807, ZN => n2793);
   U1920 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n2803, ZN => n2792);
   U1921 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, A 
                           => n2793, B => n2792, ZN => 
                           boothmul_pipelined_i_mux_out_2_14_port);
   U1922 : AOI22_X1 port map( A1 => data1_mul_11_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n2807, ZN => n2795);
   U1923 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n2803, ZN => n2794);
   U1924 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, A 
                           => n2795, B => n2794, ZN => 
                           boothmul_pipelined_i_mux_out_2_15_port);
   U1925 : AOI22_X1 port map( A1 => data1_mul_12_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n2807, ZN => n2797);
   U1926 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n2803, ZN => n2796);
   U1927 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, A 
                           => n2797, B => n2796, ZN => 
                           boothmul_pipelined_i_mux_out_2_16_port);
   U1928 : AOI22_X1 port map( A1 => data1_mul_13_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n2807, ZN => n2799);
   U1929 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n2803, ZN => n2798);
   U1930 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, A 
                           => n2799, B => n2798, ZN => 
                           boothmul_pipelined_i_mux_out_2_17_port);
   U1931 : AOI22_X1 port map( A1 => data1_mul_14_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n2807, ZN => n2801);
   U1932 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n2803, ZN => n2800);
   U1933 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, A 
                           => n2801, B => n2800, ZN => 
                           boothmul_pipelined_i_mux_out_2_18_port);
   U1934 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n2802, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n2807, ZN => n2805);
   U1935 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n2803, ZN => n2804);
   U1936 : OAI211_X1 port map( C1 => n2806, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, A 
                           => n2805, B => n2804, ZN => 
                           boothmul_pipelined_i_mux_out_2_19_port);
   U1937 : INV_X1 port map( A => n2807, ZN => n2810);
   U1938 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n3025, ZN => n2808);
   U1939 : OAI222_X1 port map( A1 => n2812, A2 => n2811, B1 => n2810, B2 => 
                           n2809, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           C2 => n2808, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1940 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_61_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_153_port, ZN
                           => n2815);
   U1941 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_38_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_176_port, ZN
                           => n2814);
   U1942 : NAND2_X1 port map( A1 => n2815, A2 => n2814, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1943 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_152_port, ZN
                           => n2817);
   U1944 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_37_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n2816);
   U1945 : NAND2_X1 port map( A1 => n2817, A2 => n2816, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1946 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_151_port, ZN
                           => n2819);
   U1947 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_36_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n2818);
   U1948 : NAND2_X1 port map( A1 => n2819, A2 => n2818, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1949 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_150_port, ZN
                           => n2821);
   U1950 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_35_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n2820);
   U1951 : NAND2_X1 port map( A1 => n2821, A2 => n2820, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1952 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_149_port, ZN
                           => n2823);
   U1953 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_34_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n2822);
   U1954 : NAND2_X1 port map( A1 => n2823, A2 => n2822, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1955 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_148_port, ZN
                           => n2825);
   U1956 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_33_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n2824);
   U1957 : NAND2_X1 port map( A1 => n2825, A2 => n2824, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1958 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_147_port, ZN
                           => n2827);
   U1959 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_32_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n2826);
   U1960 : NAND2_X1 port map( A1 => n2827, A2 => n2826, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1961 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_146_port, ZN
                           => n2829);
   U1962 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_31_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n2828);
   U1963 : NAND2_X1 port map( A1 => n2829, A2 => n2828, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U1964 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_145_port, ZN
                           => n2831);
   U1965 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_30_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n2830);
   U1966 : NAND2_X1 port map( A1 => n2831, A2 => n2830, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U1967 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_144_port, ZN
                           => n2833);
   U1968 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_29_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n2832);
   U1969 : NAND2_X1 port map( A1 => n2833, A2 => n2832, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U1970 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_143_port, ZN
                           => n2835);
   U1971 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_28_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n2834);
   U1972 : NAND2_X1 port map( A1 => n2835, A2 => n2834, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U1973 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_142_port, ZN
                           => n2837);
   U1974 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_27_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n2836);
   U1975 : NAND2_X1 port map( A1 => n2837, A2 => n2836, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U1976 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_141_port, ZN
                           => n2839);
   U1977 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_26_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n2838);
   U1978 : NAND2_X1 port map( A1 => n2839, A2 => n2838, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U1979 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_140_port, ZN
                           => n2841);
   U1980 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_25_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n2840);
   U1981 : NAND2_X1 port map( A1 => n2841, A2 => n2840, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U1982 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_139_port, ZN
                           => n2843);
   U1983 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_24_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_162_port, ZN
                           => n2842);
   U1984 : NAND2_X1 port map( A1 => n2843, A2 => n2842, ZN => 
                           boothmul_pipelined_i_mux_out_3_21_port);
   U1985 : AOI22_X1 port map( A1 => n2845, A2 => 
                           boothmul_pipelined_i_muxes_in_3_46_port, B1 => n2844
                           , B2 => boothmul_pipelined_i_muxes_in_3_138_port, ZN
                           => n2849);
   U1986 : AOI22_X1 port map( A1 => n2847, A2 => 
                           boothmul_pipelined_i_muxes_in_3_23_port, B1 => n2846
                           , B2 => boothmul_pipelined_i_muxes_in_3_161_port, ZN
                           => n2848);
   U1987 : NAND2_X1 port map( A1 => n2849, A2 => n2848, ZN => 
                           boothmul_pipelined_i_mux_out_3_22_port);
   U1988 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_65_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_165_port, ZN
                           => n2852);
   U1989 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_40_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_190_port, ZN
                           => n2851);
   U1990 : NAND2_X1 port map( A1 => n2852, A2 => n2851, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U1991 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_164_port, ZN
                           => n2854);
   U1992 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_39_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n2853);
   U1993 : NAND2_X1 port map( A1 => n2854, A2 => n2853, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U1994 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_163_port, ZN
                           => n2856);
   U1995 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_38_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n2855);
   U1996 : NAND2_X1 port map( A1 => n2856, A2 => n2855, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U1997 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_162_port, ZN
                           => n2858);
   U1998 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_37_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n2857);
   U1999 : NAND2_X1 port map( A1 => n2858, A2 => n2857, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2000 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_161_port, ZN
                           => n2860);
   U2001 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_36_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n2859);
   U2002 : NAND2_X1 port map( A1 => n2860, A2 => n2859, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2003 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_160_port, ZN
                           => n2862);
   U2004 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_35_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n2861);
   U2005 : NAND2_X1 port map( A1 => n2862, A2 => n2861, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2006 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_159_port, ZN
                           => n2864);
   U2007 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_34_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n2863);
   U2008 : NAND2_X1 port map( A1 => n2864, A2 => n2863, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2009 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_158_port, ZN
                           => n2866);
   U2010 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_33_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n2865);
   U2011 : NAND2_X1 port map( A1 => n2866, A2 => n2865, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2012 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_157_port, ZN
                           => n2868);
   U2013 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_32_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n2867);
   U2014 : NAND2_X1 port map( A1 => n2868, A2 => n2867, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2015 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_156_port, ZN
                           => n2870);
   U2016 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_31_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n2869);
   U2017 : NAND2_X1 port map( A1 => n2870, A2 => n2869, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2018 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_155_port, ZN
                           => n2872);
   U2019 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_30_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n2871);
   U2020 : NAND2_X1 port map( A1 => n2872, A2 => n2871, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2021 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_154_port, ZN
                           => n2874);
   U2022 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_29_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n2873);
   U2023 : NAND2_X1 port map( A1 => n2874, A2 => n2873, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2024 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_153_port, ZN
                           => n2876);
   U2025 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_28_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n2875);
   U2026 : NAND2_X1 port map( A1 => n2876, A2 => n2875, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2027 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_152_port, ZN
                           => n2878);
   U2028 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_27_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n2877);
   U2029 : NAND2_X1 port map( A1 => n2878, A2 => n2877, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2030 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_151_port, ZN
                           => n2880);
   U2031 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_26_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_176_port, ZN
                           => n2879);
   U2032 : NAND2_X1 port map( A1 => n2880, A2 => n2879, ZN => 
                           boothmul_pipelined_i_mux_out_4_23_port);
   U2033 : AOI22_X1 port map( A1 => n2882, A2 => 
                           boothmul_pipelined_i_muxes_in_4_50_port, B1 => n2881
                           , B2 => boothmul_pipelined_i_muxes_in_4_150_port, ZN
                           => n2886);
   U2034 : AOI22_X1 port map( A1 => n2884, A2 => 
                           boothmul_pipelined_i_muxes_in_4_25_port, B1 => n2883
                           , B2 => boothmul_pipelined_i_muxes_in_4_175_port, ZN
                           => n2885);
   U2035 : NAND2_X1 port map( A1 => n2886, A2 => n2885, ZN => 
                           boothmul_pipelined_i_mux_out_4_24_port);
   U2036 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_69_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_177_port, ZN
                           => n2889);
   U2037 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_42_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_204_port, ZN
                           => n2888);
   U2038 : NAND2_X1 port map( A1 => n2889, A2 => n2888, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2039 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_176_port, ZN
                           => n2891);
   U2040 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_41_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n2890);
   U2041 : NAND2_X1 port map( A1 => n2891, A2 => n2890, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2042 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_175_port, ZN
                           => n2893);
   U2043 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_40_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n2892);
   U2044 : NAND2_X1 port map( A1 => n2893, A2 => n2892, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2045 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_174_port, ZN
                           => n2895);
   U2046 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_39_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n2894);
   U2047 : NAND2_X1 port map( A1 => n2895, A2 => n2894, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2048 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_173_port, ZN
                           => n2897);
   U2049 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_38_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n2896);
   U2050 : NAND2_X1 port map( A1 => n2897, A2 => n2896, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2051 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_172_port, ZN
                           => n2899);
   U2052 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_37_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n2898);
   U2053 : NAND2_X1 port map( A1 => n2899, A2 => n2898, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2054 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_171_port, ZN
                           => n2901);
   U2055 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_36_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n2900);
   U2056 : NAND2_X1 port map( A1 => n2901, A2 => n2900, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2057 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_170_port, ZN
                           => n2903);
   U2058 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_35_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n2902);
   U2059 : NAND2_X1 port map( A1 => n2903, A2 => n2902, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2060 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_169_port, ZN
                           => n2905);
   U2061 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_34_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n2904);
   U2062 : NAND2_X1 port map( A1 => n2905, A2 => n2904, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2063 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_168_port, ZN
                           => n2907);
   U2064 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_33_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n2906);
   U2065 : NAND2_X1 port map( A1 => n2907, A2 => n2906, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2066 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_167_port, ZN
                           => n2909);
   U2067 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_32_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n2908);
   U2068 : NAND2_X1 port map( A1 => n2909, A2 => n2908, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2069 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_166_port, ZN
                           => n2911);
   U2070 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_31_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n2910);
   U2071 : NAND2_X1 port map( A1 => n2911, A2 => n2910, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2072 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_165_port, ZN
                           => n2913);
   U2073 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_30_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n2912);
   U2074 : NAND2_X1 port map( A1 => n2913, A2 => n2912, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2075 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_164_port, ZN
                           => n2915);
   U2076 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_29_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n2914);
   U2077 : NAND2_X1 port map( A1 => n2915, A2 => n2914, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2078 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_163_port, ZN
                           => n2917);
   U2079 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_28_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_190_port, ZN
                           => n2916);
   U2080 : NAND2_X1 port map( A1 => n2917, A2 => n2916, ZN => 
                           boothmul_pipelined_i_mux_out_5_25_port);
   U2081 : AOI22_X1 port map( A1 => n2919, A2 => 
                           boothmul_pipelined_i_muxes_in_5_54_port, B1 => n2918
                           , B2 => boothmul_pipelined_i_muxes_in_5_162_port, ZN
                           => n2923);
   U2082 : AOI22_X1 port map( A1 => n2921, A2 => 
                           boothmul_pipelined_i_muxes_in_5_27_port, B1 => n2920
                           , B2 => boothmul_pipelined_i_muxes_in_5_189_port, ZN
                           => n2922);
   U2083 : NAND2_X1 port map( A1 => n2923, A2 => n2922, ZN => 
                           boothmul_pipelined_i_mux_out_5_26_port);
   U2084 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_73_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_189_port, ZN
                           => n2926);
   U2085 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_44_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_218_port, ZN
                           => n2925);
   U2086 : NAND2_X1 port map( A1 => n2926, A2 => n2925, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2087 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_188_port, ZN
                           => n2928);
   U2088 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_43_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n2927);
   U2089 : NAND2_X1 port map( A1 => n2928, A2 => n2927, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2090 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_187_port, ZN
                           => n2930);
   U2091 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_42_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n2929);
   U2092 : NAND2_X1 port map( A1 => n2930, A2 => n2929, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2093 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_186_port, ZN
                           => n2932);
   U2094 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_41_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n2931);
   U2095 : NAND2_X1 port map( A1 => n2932, A2 => n2931, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2096 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_185_port, ZN
                           => n2934);
   U2097 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_40_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n2933);
   U2098 : NAND2_X1 port map( A1 => n2934, A2 => n2933, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2099 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_184_port, ZN
                           => n2936);
   U2100 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_39_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n2935);
   U2101 : NAND2_X1 port map( A1 => n2936, A2 => n2935, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2102 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_183_port, ZN
                           => n2938);
   U2103 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_38_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n2937);
   U2104 : NAND2_X1 port map( A1 => n2938, A2 => n2937, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2105 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_182_port, ZN
                           => n2940);
   U2106 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_37_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n2939);
   U2107 : NAND2_X1 port map( A1 => n2940, A2 => n2939, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2108 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_181_port, ZN
                           => n2942);
   U2109 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_36_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n2941);
   U2110 : NAND2_X1 port map( A1 => n2942, A2 => n2941, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2111 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_180_port, ZN
                           => n2944);
   U2112 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_35_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n2943);
   U2113 : NAND2_X1 port map( A1 => n2944, A2 => n2943, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2114 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_179_port, ZN
                           => n2946);
   U2115 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_34_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n2945);
   U2116 : NAND2_X1 port map( A1 => n2946, A2 => n2945, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2117 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_178_port, ZN
                           => n2948);
   U2118 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_33_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n2947);
   U2119 : NAND2_X1 port map( A1 => n2948, A2 => n2947, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2120 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_177_port, ZN
                           => n2950);
   U2121 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_32_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n2949);
   U2122 : NAND2_X1 port map( A1 => n2950, A2 => n2949, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2123 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_176_port, ZN
                           => n2952);
   U2124 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_31_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n2951);
   U2125 : NAND2_X1 port map( A1 => n2952, A2 => n2951, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2126 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_175_port, ZN
                           => n2954);
   U2127 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_30_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_204_port, ZN
                           => n2953);
   U2128 : NAND2_X1 port map( A1 => n2954, A2 => n2953, ZN => 
                           boothmul_pipelined_i_mux_out_6_27_port);
   U2129 : AOI22_X1 port map( A1 => n2956, A2 => 
                           boothmul_pipelined_i_muxes_in_6_58_port, B1 => n2955
                           , B2 => boothmul_pipelined_i_muxes_in_6_174_port, ZN
                           => n2960);
   U2130 : AOI22_X1 port map( A1 => n2958, A2 => 
                           boothmul_pipelined_i_muxes_in_6_29_port, B1 => n2957
                           , B2 => boothmul_pipelined_i_muxes_in_6_203_port, ZN
                           => n2959);
   U2131 : NAND2_X1 port map( A1 => n2960, A2 => n2959, ZN => 
                           boothmul_pipelined_i_mux_out_6_28_port);
   U2132 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_46_port
                           , ZN => n2963);
   U2133 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_201_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_77_port
                           , ZN => n2962);
   U2134 : NAND2_X1 port map( A1 => n2963, A2 => n2962, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2135 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_231_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_45_port
                           , ZN => n2965);
   U2136 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_200_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_76_port
                           , ZN => n2964);
   U2137 : NAND2_X1 port map( A1 => n2965, A2 => n2964, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2138 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_230_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_44_port
                           , ZN => n2967);
   U2139 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_199_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_75_port
                           , ZN => n2966);
   U2140 : NAND2_X1 port map( A1 => n2967, A2 => n2966, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2141 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_229_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_43_port
                           , ZN => n2969);
   U2142 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_198_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_74_port
                           , ZN => n2968);
   U2143 : NAND2_X1 port map( A1 => n2969, A2 => n2968, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2144 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_228_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_42_port
                           , ZN => n2971);
   U2145 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_197_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_73_port
                           , ZN => n2970);
   U2146 : NAND2_X1 port map( A1 => n2971, A2 => n2970, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2147 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_227_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_41_port
                           , ZN => n2973);
   U2148 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_196_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_72_port
                           , ZN => n2972);
   U2149 : NAND2_X1 port map( A1 => n2973, A2 => n2972, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2150 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_226_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_40_port
                           , ZN => n2975);
   U2151 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_195_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_71_port
                           , ZN => n2974);
   U2152 : NAND2_X1 port map( A1 => n2975, A2 => n2974, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2153 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_225_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_39_port
                           , ZN => n2977);
   U2154 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_194_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_70_port
                           , ZN => n2976);
   U2155 : NAND2_X1 port map( A1 => n2977, A2 => n2976, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2156 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_224_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_38_port
                           , ZN => n2979);
   U2157 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_193_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_69_port
                           , ZN => n2978);
   U2158 : NAND2_X1 port map( A1 => n2979, A2 => n2978, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2159 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_223_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_37_port
                           , ZN => n2981);
   U2160 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_192_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_68_port
                           , ZN => n2980);
   U2161 : NAND2_X1 port map( A1 => n2981, A2 => n2980, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2162 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_222_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_36_port
                           , ZN => n2983);
   U2163 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_191_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_67_port
                           , ZN => n2982);
   U2164 : NAND2_X1 port map( A1 => n2983, A2 => n2982, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2165 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_221_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_35_port
                           , ZN => n2985);
   U2166 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_190_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_66_port
                           , ZN => n2984);
   U2167 : NAND2_X1 port map( A1 => n2985, A2 => n2984, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2168 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_220_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_34_port
                           , ZN => n2987);
   U2169 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_189_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_65_port
                           , ZN => n2986);
   U2170 : NAND2_X1 port map( A1 => n2987, A2 => n2986, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2171 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_219_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_33_port
                           , ZN => n2989);
   U2172 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_188_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_64_port
                           , ZN => n2988);
   U2173 : NAND2_X1 port map( A1 => n2989, A2 => n2988, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2174 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_32_port
                           , ZN => n2991);
   U2175 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_187_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_63_port
                           , ZN => n2990);
   U2176 : NAND2_X1 port map( A1 => n2991, A2 => n2990, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2177 : AOI22_X1 port map( A1 => n2993, A2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, B1 => 
                           n2992, B2 => boothmul_pipelined_i_muxes_in_7_31_port
                           , ZN => n2997);
   U2178 : AOI22_X1 port map( A1 => n2995, A2 => 
                           boothmul_pipelined_i_muxes_in_7_186_port, B1 => 
                           n2994, B2 => boothmul_pipelined_i_muxes_in_7_62_port
                           , ZN => n2996);
   U2179 : NAND2_X1 port map( A1 => n2997, A2 => n2996, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2180 : OAI222_X1 port map( A1 => n3018, A2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, 
                           B1 => n3013, B2 => n2998, C1 => n3012, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           ZN => boothmul_pipelined_i_sum_out_1_1_port);
   U2181 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN 
                           => n3000);
   U2182 : OAI222_X1 port map( A1 => n3013, A2 => n3000, B1 => n3012, B2 => 
                           n2999, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2183 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN 
                           => n3001);
   U2184 : OAI222_X1 port map( A1 => n3013, A2 => n3001, B1 => n3012, B2 => 
                           n3000, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2185 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN 
                           => n3002);
   U2186 : OAI222_X1 port map( A1 => n3013, A2 => n3002, B1 => n3012, B2 => 
                           n3001, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2187 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN 
                           => n3003);
   U2188 : OAI222_X1 port map( A1 => n3013, A2 => n3003, B1 => n3012, B2 => 
                           n3002, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2189 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN 
                           => n3004);
   U2190 : OAI222_X1 port map( A1 => n3013, A2 => n3004, B1 => n3012, B2 => 
                           n3003, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2191 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN 
                           => n3005);
   U2192 : OAI222_X1 port map( A1 => n3013, A2 => n3005, B1 => n3012, B2 => 
                           n3004, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2193 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN 
                           => n3006);
   U2194 : OAI222_X1 port map( A1 => n3013, A2 => n3006, B1 => n3012, B2 => 
                           n3005, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2195 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN 
                           => n3007);
   U2196 : OAI222_X1 port map( A1 => n3013, A2 => n3007, B1 => n3012, B2 => 
                           n3006, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2197 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN 
                           => n3008);
   U2198 : OAI222_X1 port map( A1 => n3013, A2 => n3008, B1 => n3012, B2 => 
                           n3007, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2199 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN 
                           => n3009);
   U2200 : OAI222_X1 port map( A1 => n3013, A2 => n3009, B1 => n3012, B2 => 
                           n3008, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2201 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN 
                           => n3010);
   U2202 : OAI222_X1 port map( A1 => n3013, A2 => n3010, B1 => n3012, B2 => 
                           n3009, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2203 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN 
                           => n3011);
   U2204 : OAI222_X1 port map( A1 => n3013, A2 => n3011, B1 => n3012, B2 => 
                           n3010, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, 
                           C2 => n3018, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2205 : INV_X1 port map( A => n3012, ZN => n3016);
   U2206 : INV_X1 port map( A => n3013, ZN => n3015);
   U2207 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n3016, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n3015, ZN => n3014);
   U2208 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           B2 => n3018, A => n3014, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2209 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n3016, B1 => n3015, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n3017);
   U2210 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           B2 => n3018, A => n3017, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, 
      n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, 
      n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
      n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, 
      n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, 
      n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, 
      n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
      n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, 
      n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, 
      n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
      n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, 
      n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, 
      n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
      n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, 
      n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, 
      n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, 
      n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, 
      n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, 
      n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, 
      n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
      n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, 
      n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
      n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, 
      n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, 
      n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, 
      n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, 
      n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, 
      n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, 
      n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, 
      n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, 
      n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, 
      n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, 
      n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, 
      n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, 
      n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, 
      n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, 
      n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, 
      n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, 
      n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
      n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, 
      n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, 
      n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, 
      n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, 
      n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, 
      n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, 
      n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, 
      n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
      n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, 
      n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, 
      n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, 
      n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, 
      n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
      n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, 
      n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, 
      n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, 
      n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, 
      n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, 
      n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, 
      n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, 
      n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
      n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, 
      n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, 
      n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, 
      n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
      n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, 
      n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, 
      n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
      n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, 
      n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
      n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, 
      n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
      n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, 
      n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, 
      n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590 : std_logic;

begin
   
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n6517);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n6266);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1527);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1528);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n6246);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n6236);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n6478);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n6727);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n5977);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n6710);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n5953);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n6105);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n5839);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n5827);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n6337);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n6569);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n6067);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n5786);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n6308);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n5773);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n6036);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n6520);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n6192);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n5923);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n6674);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n6661);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n6400);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n6153);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n6397);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n6388);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n6129);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n6374);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n6613);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n6505);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1529);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1530);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n6245);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n6235);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n6477);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n6464);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n6224);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n5963);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n6201);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n6442);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n6098);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n5826);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n6580);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n6330);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n5800);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n6556);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n6043);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n6296);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n5766);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n6027);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n6275);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n6687);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n6412);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n5914);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n5901);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n6152);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n6645);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n6387);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n6128);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n5853);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n6612);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n6353);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1531);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1532);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n6244);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n6486);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n6230);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n5981);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n5976);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n6709);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n6200);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n6701);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n6427);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n5825);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n6579);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n6568);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n5799);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n5785);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n6546);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n6295);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n6527);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n6026);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n5740);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n6504);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n6174);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n6660);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n5900);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n5890);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n6644);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n6635);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n5866);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n5852);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n6365);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n6594);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n6097);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1533);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n6000);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n5991);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n6476);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n6726);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n5975);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n6708);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n5952);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n6441);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n6191);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n6686);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n6578);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n6329);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n6066);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n6555);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n6545);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n6294);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n5765);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n5752);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n5739);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n6503);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1534);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n6170);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n5899);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n5889);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n5878);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n6634);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n6127);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n6623);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n6611);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n5847);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n5838);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n5824);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n6490);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n5990);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n6475);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n6725);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n6223);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n6209);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n6450);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n6700);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n6190);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n6423);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n6673);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n6328);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n6065);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n6051);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n6307);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n6293);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n5764);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n6025);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n6516);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n6265);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1535);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1536);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n5898);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n6151);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n6396);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n6633);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n6126);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n6373);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n6610);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n5846);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n5837);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n6086);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n6577);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n5989);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n6474);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n6227);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n5974);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n6707);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n5951);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n6440);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n6189);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n6685);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n6672);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n6405);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n5798);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n6050);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n6544);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n6536);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n6282);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n6024);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n5738);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n6264);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1537);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1538);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n6243);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n5888);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n6137);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n5871);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n5865);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n6622);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n6364);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n6104);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n5836);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n6085);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n6576);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n6327);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n6741);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n6724);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n6222);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n6208);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n5950);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n6699);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n5935);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n6422);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n5921);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n6404);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n6653);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n6554);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n6306);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n5772);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n6035);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n6280);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n6015);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n6502);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1539);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1540);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n6756);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n6485);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n6395);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n6632);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n6125);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n6113);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n6609);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n6352);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n6343);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n6084);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n5809);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n6326);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n5797);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n6463);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n5973);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n6706);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n6199);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n6439);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n5934);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n6684);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n6671);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n5913);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n6165);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n6150);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n6543);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n6535);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n5763);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n6023);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n6014);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n6263);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1541);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1542);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n5999);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n6234);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n6473);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n6386);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n5864);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n6621);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n6363);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n6351);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n6096);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n5823);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n6077);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n6567);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n5796);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n6314);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n5972);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n6455);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n6198);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n6698);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n5933);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n6179);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n6173);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n5912);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n6164);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n5887);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n6394);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n6292);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n5762);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n5751);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n6274);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n6501);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1543);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1544);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n6755);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n6484);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n6740);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n6723);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n6124);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n6112);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n6608);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n6350);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n5835);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n5822);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n6336);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n6566);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n6064);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n6049);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n6542);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n5962);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n6197);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n6697);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n6689);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n6421);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n6670);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n5911);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n5897);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n6149);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n5877);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n6631);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n6281);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n6021);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n6013);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n6261);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1545);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1546);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n6242);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n6748);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n6472);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n6462);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n5971);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n6372);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n6606);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n6349);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n5834);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n5821);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n6076);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n6564);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n5794);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n6313);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n6042);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n6534);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n5948);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n6437);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n5931);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n6420);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n6172);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n6659);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n6162);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n6148);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n6393);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n6630);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n6123);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n6022);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n6515);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n6262);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1547);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1548);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n6754);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n5988);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n6471);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n6461);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n6221);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n6207);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n6607);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n5845);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n6342);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n6083);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n5808);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n6565);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n5795);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n6048);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n5778);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n6291);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n6526);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n6438);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n5932);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n6683);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n5920);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n6169);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n6163);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n6398);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n6643);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n6385);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n5863);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n6620);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n5747);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n6512);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n6497);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1549);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n6241);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n6747);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n6739);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n6722);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n5970);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n5961);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n5949);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n6360);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n5843);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n6094);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n5818);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n6574);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n6563);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n6060);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n6046);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n6303);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n6288);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n5758);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n6037);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n6028);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n6276);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n6506);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1550);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1551);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n6492);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n6237);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n6743);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n6729);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n5979);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n6375);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n6106);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n6596);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n6100);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n5829);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n6338);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n6570);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n5801);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n5787);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n6310);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n6538);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n5954);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n6702);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n6193);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n6180);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n6413);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n6662);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n6401);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n6154);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n5879);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n6389);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n5867);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n6521);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n5741);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n6267);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1552);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1553);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n6491);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n5992);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n6742);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n6728);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n5978);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n6210);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n6366);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n6595);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n6099);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n5828);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n6581);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n6331);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n6068);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n6052);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n6309);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n6537);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n5767);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n6443);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n5936);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n6688);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n6675);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n5915);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n5902);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n5891);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n6646);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n6636);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n6130);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n5854);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n5774);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n5768);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n5753);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n6277);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n6507);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1554);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1555);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1556);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1557);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1558);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1559);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n6132);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n5855);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n6614);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n6597);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n5841);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n6583);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n5810);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n6333);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n6070);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n6557);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n6547);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n6211);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n6703);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n6445);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n5937);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n6425);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n6676);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n5917);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n6654);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n6155);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n5880);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n5872);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n6432);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n5929);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n6680);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n5918);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n6167);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n6650);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n6145);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n5876);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n6383);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n6120);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n6370);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n6272);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n6498);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1560);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1561);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n6752);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n6482);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n6736);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n6718);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n6219);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n5960);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n5945);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n6102);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n6586);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n5819);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n5806);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n6322);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n6061);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n5783);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n6541);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n6532);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n5759);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n5748);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n6186);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n6681);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n6668);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n5909);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n6161);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n5885);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n6135);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n5870);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n6121);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n6618);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n6361);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n6499);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1562);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1563);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n6489);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n6746);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n6469);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n6719);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n5967);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n6204);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n6448);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n6433);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n5833);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n5820);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n6575);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n6323);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n5793);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n6553);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n6041);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n6289);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n5760);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n5749);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n6513);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n6666);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n6657);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n6158);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n6144);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n6641);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n5869);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n5859);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n6109);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n6602);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n6347);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n6093);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1564);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n5996);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n6481);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n6733);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n6716);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n5965);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n6452);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n5944);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n6431);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n5927);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n6176);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n6334);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n6321);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n5792);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n6045);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n6301);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n6531);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n6033);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n6279);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n6012);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n6259);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1565);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n6658);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n6159);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n5883);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n5874);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n6627);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n6119);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n5851);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n6603);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n6101);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n6585);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n5817);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n6751);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n5985);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n6734);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n6460);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n5966);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n6453);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n6196);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n6695);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n5928);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n6419);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n6171);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n6562);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n6059);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n6552);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n6302);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n5771);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n5757);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n6019);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n6271);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n6496);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1566);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1567);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n5922);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n5919);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n6403);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n6651);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n5886);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n6136);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n6628);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n6122);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n6619);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n6604);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n5844);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1568);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1569);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n5997);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n6233);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n6470);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n6720);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n6220);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n6705);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n6449);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n6434);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n6187);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n6082);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n5807);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n6325);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n6063);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n5784);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n6305);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n6290);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n6034);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n5750);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n6514);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n6500);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n6411);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n5910);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n6652);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n6147);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n6642);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n6629);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n5862);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n6111);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n6362);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n6593);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n6587);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1570);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n5998);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n6483);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n6738);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n6721);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n5969);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n6206);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n5947);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n6436);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n5930);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n6178);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n6340);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n6075);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n6320);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n6058);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n5782);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n6540);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n6287);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n5756);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n6018);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n6511);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n6258);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n6143);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n6391);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n6626);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n5858);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n6369);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n6358);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n6592);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n6092);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n6079);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n6074);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n6319);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n6732);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n6459);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n6217);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n5959);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n5943);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n6430);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n5926);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n6679);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n6665);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n6166);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n5896);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n6047);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n6304);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n6533);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n5761);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n6020);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n6273);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n6260);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1571);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1572);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n6487);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n6232);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n6392);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n6384);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n5861);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n6371);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n6605);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n6103);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n6095);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n6081);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n6335);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n6324);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n6062);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n5980);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n5968);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n6205);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n5946);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n6435);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n6188);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n6682);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n6669);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n6168);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n6399);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n6146);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n6311);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n6039);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n6038);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n6522);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n5742);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n6268);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1573);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1574);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n6753);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n5987);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n6737);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n6160);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n5884);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n5875);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n6382);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n5860);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n6110);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n6359);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n6348);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n5832);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n6080);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n6573);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n5986);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n6735);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n6717);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n6218);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n6454);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n6447);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n6696);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n6185);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n6177);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n6667);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n5908);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n6561);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n5791);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n6551);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n5777);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n6286);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n6032);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n6017);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n6510);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n6256);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1575);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n6488);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n6157);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n6142);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n6640);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n6381);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n6118);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n6617);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n6357);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n6346);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n6091);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n5816);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n5805);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n6745);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n6468);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n6715);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n5964);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n6203);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n5942);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n6429);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n5925);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n6418);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n6664);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n5907);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n6057);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n5781);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n6300);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n6530);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n6525);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n5746);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n6011);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n6257);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1576);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1577);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n6240);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n6637);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n6131);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n6624);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n6367);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n5848);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n5840);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n6087);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n6582);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n6332);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n6069);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n6315);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n6225);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n6711);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n6202);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n6444);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n6690);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n6424);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n6175);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n5916);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n5903);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n5892);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n6647);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n6299);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n6285);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n6031);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n5745);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n6509);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n6495);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1578);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n6247);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n5993);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n6479);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n6465);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n6380);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n6117);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n5850);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n6601);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n6591);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n6584);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n5815);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n5804);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n6318);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n6056);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n5780);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n6216);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n6451);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n5941);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n6694);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n5924);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n6417);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n6410);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n5906);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n6649);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n5882);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n6639);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n6297);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n5769);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n6523);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n5743);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n6269);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1579);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n6239);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n6231);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n6229);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n6714);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n6089);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n5814);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n6072);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n6317);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n5790);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n6550);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n6040);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n6529);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n6030);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n6278);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n5737);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n6416);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n6409);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n6656);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n5894);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n6140);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n6134);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n6625);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n6116);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n6368);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n6600);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n6344);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1580);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1581);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n5995);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n6744);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n6466);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n6457);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n6214);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n5957);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n5940);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n6692);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n6183);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n6339);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n6073);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n6560);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n6055);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n5779);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n6298);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n6284);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n5755);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n6519);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n6010);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n6494);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n6663);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n6402);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n5895);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n6141);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n5873);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n6379);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n5857);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n6108);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n6356);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n6345);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n6090);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n6750);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n5984);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n6467);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n6458);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n6215);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n5958);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n6195);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n6693);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n6184);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n6678);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n6354);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n5842);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n5831);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n6078);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n6572);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n6559);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n5788);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n6044);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n6539);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n5770);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n5754);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n6691);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n6181);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n6415);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n6407);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n5904);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n5893);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n6138);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n6638);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n6377);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n5856);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n6615);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n6270);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n6493);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1582);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1583);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n5994);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n5982);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n6731);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n6456);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n6212);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n6704);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n6194);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n6590);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n6088);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n5813);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n5803);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n6316);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n5789);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n6549);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n5776);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n6283);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n6029);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n6016);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n6182);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n6677);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n6408);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n5905);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n6648);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n6139);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n6390);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n6378);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n6115);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n6616);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n6355);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n6255);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1584);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1585);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n6749);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n5983);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n6228);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n6713);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n6213);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n5956);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n5939);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n6428);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n5868);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n6376);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n6107);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n6598);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n6588);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n5830);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n5811);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n6571);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n6071);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n6053);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n6548);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n6712);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n5955);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n6446);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n5938);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n6426);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n6414);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n6406);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n6655);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n6156);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n5881);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n6133);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n6524);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n5744);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n6009);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n6253);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1586);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1587);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n6248);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n6238);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n6480);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n6730);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n6226);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n5849);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n6599);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n6589);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n6341);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n5812);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n5802);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n6558);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n6054);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n6312);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n5775);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n6528);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n6005);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n6252);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n5733);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n6251);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n6250);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n6004);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n6003);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n6002);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n6001);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n6249);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n6114);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n6518);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n6508);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n6254);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1588);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1589);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n5736);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n5735);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n6008);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n6007);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n5734);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n6006);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1590);
   U3 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n3995, ZN => n3996);
   U4 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n3992, ZN => n3993);
   U5 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n3989, ZN => n3990);
   U6 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4092, ZN => n4093);
   U7 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4057, ZN => n4058);
   U8 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4050, ZN => n4051);
   U9 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4007, ZN => n4008);
   U10 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4026, ZN => n4029);
   U11 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4047, ZN => n4048);
   U12 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4003, ZN => n4004);
   U13 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4044, ZN => n4045);
   U14 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n4041, ZN => n4042);
   U15 : NAND2_X2 port map( A1 => RESET_BAR, A2 => DATAIN(2), ZN => n4175);
   U16 : NAND2_X2 port map( A1 => RESET_BAR, A2 => DATAIN(17), ZN => n4158);
   U17 : NAND2_X2 port map( A1 => RESET_BAR, A2 => DATAIN(6), ZN => n4171);
   U18 : NAND2_X2 port map( A1 => RESET_BAR, A2 => DATAIN(5), ZN => n4172);
   U19 : NAND3_X2 port map( A1 => RESET_BAR, A2 => ENABLE, A3 => RD1, ZN => 
                           n5732);
   U20 : NAND3_X2 port map( A1 => RESET_BAR, A2 => ENABLE, A3 => RD2, ZN => 
                           n4958);
   U21 : INV_X2 port map( A => n4976, ZN => n5717);
   U22 : INV_X2 port map( A => n4975, ZN => n5720);
   U23 : INV_X2 port map( A => n4977, ZN => n5707);
   U24 : INV_X2 port map( A => n4978, ZN => n5718);
   U25 : INV_X2 port map( A => n4974, ZN => n5708);
   U26 : INV_X2 port map( A => n4197, ZN => n4941);
   U27 : INV_X2 port map( A => n4196, ZN => n4933);
   U28 : INV_X2 port map( A => n4979, ZN => n5671);
   U29 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n4002, ZN => n4006);
   U30 : INV_X1 port map( A => ADD_WR(0), ZN => n4002);
   U31 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => n4104, ZN => n4099);
   U32 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n4006, ZN => n4117);
   U33 : CLKBUF_X1 port map( A => n4176, Z => n4033);
   U34 : CLKBUF_X1 port map( A => n4174, Z => n4032);
   U35 : CLKBUF_X1 port map( A => n4097, Z => n4095);
   U36 : CLKBUF_X1 port map( A => n4063, Z => n4061);
   U37 : CLKBUF_X1 port map( A => n4005, Z => n4003);
   U38 : CLKBUF_X1 port map( A => n3987, Z => n3985);
   U39 : CLKBUF_X1 port map( A => n4170, Z => n4030);
   U40 : CLKBUF_X1 port map( A => n4054, Z => n4056);
   U41 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n4106);
   U42 : INV_X1 port map( A => ADD_WR(4), ZN => n3984);
   U43 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n3984, ZN => n4036);
   U44 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => n4036, ZN => n4012);
   U45 : NAND2_X1 port map( A1 => n4106, A2 => n4012, ZN => n3987);
   U46 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n3985, ZN => n3986);
   U47 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(31), ZN => n4107);
   U48 : OAI22_X1 port map( A1 => n6253, A2 => n3986, B1 => n4107, B2 => n3985,
                           ZN => n2166);
   U49 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(30), ZN => n4145);
   U50 : CLKBUF_X1 port map( A => n4145, Z => n4081);
   U51 : OAI22_X1 port map( A1 => n6254, A2 => n3986, B1 => n3985, B2 => n4081,
                           ZN => n2165);
   U52 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(29), ZN => n4146);
   U53 : CLKBUF_X1 port map( A => n4146, Z => n4082);
   U54 : OAI22_X1 port map( A1 => n6493, A2 => n3986, B1 => n3985, B2 => n4082,
                           ZN => n2164);
   U55 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(28), ZN => n4147);
   U56 : CLKBUF_X1 port map( A => n4147, Z => n4083);
   U57 : OAI22_X1 port map( A1 => n6255, A2 => n3986, B1 => n3985, B2 => n4083,
                           ZN => n2163);
   U58 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(27), ZN => n4148);
   U59 : CLKBUF_X1 port map( A => n4148, Z => n4084);
   U60 : OAI22_X1 port map( A1 => n6494, A2 => n3986, B1 => n3985, B2 => n4084,
                           ZN => n2162);
   U61 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(26), ZN => n4149);
   U62 : CLKBUF_X1 port map( A => n4149, Z => n4085);
   U63 : OAI22_X1 port map( A1 => n6495, A2 => n3986, B1 => n3985, B2 => n4085,
                           ZN => n2161);
   U64 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(25), ZN => n4150);
   U65 : CLKBUF_X1 port map( A => n4150, Z => n4086);
   U66 : OAI22_X1 port map( A1 => n6256, A2 => n3986, B1 => n3985, B2 => n4086,
                           ZN => n2160);
   U67 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(24), ZN => n4151);
   U68 : CLKBUF_X1 port map( A => n4151, Z => n4087);
   U69 : OAI22_X1 port map( A1 => n6257, A2 => n3986, B1 => n3985, B2 => n4087,
                           ZN => n2159);
   U70 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(23), ZN => n4152);
   U71 : CLKBUF_X1 port map( A => n4152, Z => n4013);
   U72 : OAI22_X1 port map( A1 => n6258, A2 => n3986, B1 => n3987, B2 => n4013,
                           ZN => n2158);
   U73 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(22), ZN => n4153);
   U74 : CLKBUF_X1 port map( A => n4153, Z => n4014);
   U75 : OAI22_X1 port map( A1 => n6259, A2 => n3986, B1 => n3987, B2 => n4014,
                           ZN => n2157);
   U76 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(21), ZN => n4154);
   U77 : CLKBUF_X1 port map( A => n4154, Z => n4015);
   U78 : OAI22_X1 port map( A1 => n6496, A2 => n3986, B1 => n3987, B2 => n4015,
                           ZN => n2156);
   U79 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(20), ZN => n4155);
   U80 : CLKBUF_X1 port map( A => n4155, Z => n4016);
   U81 : OAI22_X1 port map( A1 => n6497, A2 => n3986, B1 => n3987, B2 => n4016,
                           ZN => n2155);
   U82 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(19), ZN => n4156);
   U83 : CLKBUF_X1 port map( A => n4156, Z => n4017);
   U84 : OAI22_X1 port map( A1 => n6498, A2 => n3986, B1 => n3987, B2 => n4017,
                           ZN => n2154);
   U85 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(18), ZN => n4157);
   U86 : CLKBUF_X1 port map( A => n4157, Z => n4018);
   U87 : OAI22_X1 port map( A1 => n6499, A2 => n3986, B1 => n3987, B2 => n4018,
                           ZN => n2153);
   U88 : OAI22_X1 port map( A1 => n6260, A2 => n3986, B1 => n3987, B2 => n4158,
                           ZN => n2152);
   U89 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(16), ZN => n4159);
   U90 : CLKBUF_X1 port map( A => n4159, Z => n4019);
   U91 : OAI22_X1 port map( A1 => n6500, A2 => n3986, B1 => n3987, B2 => n4019,
                           ZN => n2151);
   U92 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(15), ZN => n4160);
   U93 : CLKBUF_X1 port map( A => n4160, Z => n4020);
   U94 : OAI22_X1 port map( A1 => n6261, A2 => n3986, B1 => n3987, B2 => n4020,
                           ZN => n2150);
   U95 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(14), ZN => n4161);
   U96 : CLKBUF_X1 port map( A => n4161, Z => n4021);
   U97 : OAI22_X1 port map( A1 => n6262, A2 => n3986, B1 => n3987, B2 => n4021,
                           ZN => n2149);
   U98 : CLKBUF_X1 port map( A => n3986, Z => n3988);
   U99 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(13), ZN => n4162);
   U100 : CLKBUF_X1 port map( A => n4162, Z => n4022);
   U101 : OAI22_X1 port map( A1 => n6501, A2 => n3988, B1 => n3987, B2 => n4022
                           , ZN => n2148);
   U102 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(12), ZN => n4163);
   U103 : CLKBUF_X1 port map( A => n4163, Z => n4023);
   U104 : OAI22_X1 port map( A1 => n6263, A2 => n3986, B1 => n3985, B2 => n4023
                           , ZN => n2147);
   U105 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(11), ZN => n4164);
   U106 : CLKBUF_X1 port map( A => n4164, Z => n4024);
   U107 : OAI22_X1 port map( A1 => n6502, A2 => n3986, B1 => n3985, B2 => n4024
                           , ZN => n2146);
   U108 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(10), ZN => n4165);
   U109 : CLKBUF_X1 port map( A => n4165, Z => n4025);
   U110 : OAI22_X1 port map( A1 => n6264, A2 => n3986, B1 => n3985, B2 => n4025
                           , ZN => n2145);
   U111 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(9), ZN => n4167);
   U112 : CLKBUF_X1 port map( A => n4167, Z => n4027);
   U113 : OAI22_X1 port map( A1 => n6265, A2 => n3986, B1 => n3985, B2 => n4027
                           , ZN => n2144);
   U114 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(8), ZN => n4168);
   U115 : CLKBUF_X1 port map( A => n4168, Z => n4028);
   U116 : OAI22_X1 port map( A1 => n6503, A2 => n3986, B1 => n3985, B2 => n4028
                           , ZN => n2143);
   U117 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(7), ZN => n4170);
   U118 : OAI22_X1 port map( A1 => n6504, A2 => n3988, B1 => n3987, B2 => n4030
                           , ZN => n2142);
   U119 : OAI22_X1 port map( A1 => n6505, A2 => n3988, B1 => n3987, B2 => n4171
                           , ZN => n2141);
   U120 : OAI22_X1 port map( A1 => n6266, A2 => n3988, B1 => n3987, B2 => n4172
                           , ZN => n2140);
   U121 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(4), ZN => n4173);
   U122 : CLKBUF_X1 port map( A => n4173, Z => n4031);
   U123 : OAI22_X1 port map( A1 => n6267, A2 => n3988, B1 => n3987, B2 => n4031
                           , ZN => n2139);
   U124 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(3), ZN => n4174);
   U125 : OAI22_X1 port map( A1 => n6506, A2 => n3988, B1 => n3987, B2 => n4032
                           , ZN => n2138);
   U126 : OAI22_X1 port map( A1 => n6268, A2 => n3988, B1 => n3987, B2 => n4175
                           , ZN => n2137);
   U127 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(1), ZN => n4176);
   U128 : OAI22_X1 port map( A1 => n6507, A2 => n3988, B1 => n3987, B2 => n4033
                           , ZN => n2136);
   U129 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(0), ZN => n4178);
   U130 : CLKBUF_X1 port map( A => n4178, Z => n4035);
   U131 : OAI22_X1 port map( A1 => n6269, A2 => n3988, B1 => n3987, B2 => n4035
                           , ZN => n2135);
   U132 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n4002, ZN 
                           => n4112);
   U133 : NAND2_X1 port map( A1 => n4012, A2 => n4112, ZN => n3991);
   U134 : CLKBUF_X1 port map( A => n3991, Z => n3989);
   U135 : OAI22_X1 port map( A1 => n6009, A2 => n3990, B1 => n4107, B2 => n3989
                           , ZN => n2134);
   U136 : OAI22_X1 port map( A1 => n6508, A2 => n3990, B1 => n4081, B2 => n3989
                           , ZN => n2133);
   U137 : OAI22_X1 port map( A1 => n6270, A2 => n3990, B1 => n4082, B2 => n3989
                           , ZN => n2132);
   U138 : OAI22_X1 port map( A1 => n5737, A2 => n3990, B1 => n4083, B2 => n3989
                           , ZN => n2131);
   U139 : OAI22_X1 port map( A1 => n6010, A2 => n3990, B1 => n4084, B2 => n3989
                           , ZN => n2130);
   U140 : OAI22_X1 port map( A1 => n6509, A2 => n3990, B1 => n4085, B2 => n3989
                           , ZN => n2129);
   U141 : OAI22_X1 port map( A1 => n6510, A2 => n3990, B1 => n4086, B2 => n3989
                           , ZN => n2128);
   U142 : OAI22_X1 port map( A1 => n6011, A2 => n3990, B1 => n4087, B2 => n3989
                           , ZN => n2127);
   U143 : OAI22_X1 port map( A1 => n6511, A2 => n3990, B1 => n4013, B2 => n3989
                           , ZN => n2126);
   U144 : OAI22_X1 port map( A1 => n6012, A2 => n3990, B1 => n4014, B2 => n3989
                           , ZN => n2125);
   U145 : OAI22_X1 port map( A1 => n6271, A2 => n3990, B1 => n4015, B2 => n3989
                           , ZN => n2124);
   U146 : OAI22_X1 port map( A1 => n6512, A2 => n3990, B1 => n4016, B2 => n3991
                           , ZN => n2123);
   U147 : OAI22_X1 port map( A1 => n6272, A2 => n3990, B1 => n4017, B2 => n3991
                           , ZN => n2122);
   U148 : OAI22_X1 port map( A1 => n6513, A2 => n3990, B1 => n4018, B2 => n3991
                           , ZN => n2121);
   U149 : OAI22_X1 port map( A1 => n6273, A2 => n3990, B1 => n4158, B2 => n3991
                           , ZN => n2120);
   U150 : OAI22_X1 port map( A1 => n6514, A2 => n3990, B1 => n4019, B2 => n3991
                           , ZN => n2119);
   U151 : OAI22_X1 port map( A1 => n6013, A2 => n3990, B1 => n4020, B2 => n3991
                           , ZN => n2118);
   U152 : OAI22_X1 port map( A1 => n6515, A2 => n3990, B1 => n4021, B2 => n3991
                           , ZN => n2117);
   U153 : OAI22_X1 port map( A1 => n6274, A2 => n3990, B1 => n4022, B2 => n3991
                           , ZN => n2116);
   U154 : OAI22_X1 port map( A1 => n6014, A2 => n3990, B1 => n4023, B2 => n3991
                           , ZN => n2115);
   U155 : OAI22_X1 port map( A1 => n6015, A2 => n3990, B1 => n4024, B2 => n3989
                           , ZN => n2114);
   U156 : OAI22_X1 port map( A1 => n5738, A2 => n3990, B1 => n4025, B2 => n3989
                           , ZN => n2113);
   U157 : OAI22_X1 port map( A1 => n6516, A2 => n3990, B1 => n4027, B2 => n3989
                           , ZN => n2112);
   U158 : OAI22_X1 port map( A1 => n5739, A2 => n3990, B1 => n4028, B2 => n3991
                           , ZN => n2111);
   U159 : OAI22_X1 port map( A1 => n5740, A2 => n3990, B1 => n4030, B2 => n3991
                           , ZN => n2110);
   U160 : OAI22_X1 port map( A1 => n6275, A2 => n3990, B1 => n4171, B2 => n3991
                           , ZN => n2109);
   U161 : OAI22_X1 port map( A1 => n6517, A2 => n3990, B1 => n4172, B2 => n3991
                           , ZN => n2108);
   U162 : OAI22_X1 port map( A1 => n5741, A2 => n3990, B1 => n4031, B2 => n3991
                           , ZN => n2107);
   U163 : OAI22_X1 port map( A1 => n6276, A2 => n3990, B1 => n4032, B2 => n3991
                           , ZN => n2106);
   U164 : OAI22_X1 port map( A1 => n5742, A2 => n3990, B1 => n4175, B2 => n3991
                           , ZN => n2105);
   U165 : OAI22_X1 port map( A1 => n6277, A2 => n3990, B1 => n4033, B2 => n3991
                           , ZN => n2104);
   U166 : OAI22_X1 port map( A1 => n5743, A2 => n3990, B1 => n4035, B2 => n3991
                           , ZN => n2103);
   U167 : NAND2_X1 port map( A1 => n4012, A2 => n4117, ZN => n3994);
   U168 : CLKBUF_X1 port map( A => n3994, Z => n3992);
   U169 : OAI22_X1 port map( A1 => n5744, A2 => n3993, B1 => n4107, B2 => n3992
                           , ZN => n2102);
   U170 : OAI22_X1 port map( A1 => n6518, A2 => n3993, B1 => n4081, B2 => n3992
                           , ZN => n2101);
   U171 : OAI22_X1 port map( A1 => n6016, A2 => n3993, B1 => n4082, B2 => n3992
                           , ZN => n2100);
   U172 : OAI22_X1 port map( A1 => n6278, A2 => n3993, B1 => n4083, B2 => n3992
                           , ZN => n2099);
   U173 : OAI22_X1 port map( A1 => n6519, A2 => n3993, B1 => n4084, B2 => n3992
                           , ZN => n2098);
   U174 : OAI22_X1 port map( A1 => n5745, A2 => n3993, B1 => n4085, B2 => n3992
                           , ZN => n2097);
   U175 : OAI22_X1 port map( A1 => n6017, A2 => n3993, B1 => n4086, B2 => n3992
                           , ZN => n2096);
   U176 : OAI22_X1 port map( A1 => n5746, A2 => n3993, B1 => n4087, B2 => n3992
                           , ZN => n2095);
   U177 : OAI22_X1 port map( A1 => n6018, A2 => n3993, B1 => n4013, B2 => n3992
                           , ZN => n2094);
   U178 : OAI22_X1 port map( A1 => n6279, A2 => n3993, B1 => n4014, B2 => n3992
                           , ZN => n2093);
   U179 : OAI22_X1 port map( A1 => n6019, A2 => n3993, B1 => n4015, B2 => n3992
                           , ZN => n2092);
   U180 : OAI22_X1 port map( A1 => n5747, A2 => n3993, B1 => n4016, B2 => n3994
                           , ZN => n2091);
   U181 : OAI22_X1 port map( A1 => n5748, A2 => n3993, B1 => n4017, B2 => n3994
                           , ZN => n2090);
   U182 : OAI22_X1 port map( A1 => n5749, A2 => n3993, B1 => n4018, B2 => n3994
                           , ZN => n2089);
   U183 : OAI22_X1 port map( A1 => n6020, A2 => n3993, B1 => n4158, B2 => n3994
                           , ZN => n2088);
   U184 : OAI22_X1 port map( A1 => n5750, A2 => n3993, B1 => n4019, B2 => n3994
                           , ZN => n2087);
   U185 : OAI22_X1 port map( A1 => n6021, A2 => n3993, B1 => n4020, B2 => n3994
                           , ZN => n2086);
   U186 : OAI22_X1 port map( A1 => n6022, A2 => n3993, B1 => n4021, B2 => n3994
                           , ZN => n2085);
   U187 : OAI22_X1 port map( A1 => n5751, A2 => n3993, B1 => n4022, B2 => n3994
                           , ZN => n2084);
   U188 : OAI22_X1 port map( A1 => n6023, A2 => n3993, B1 => n4023, B2 => n3994
                           , ZN => n2083);
   U189 : OAI22_X1 port map( A1 => n6280, A2 => n3993, B1 => n4024, B2 => n3992
                           , ZN => n2082);
   U190 : OAI22_X1 port map( A1 => n6024, A2 => n3993, B1 => n4025, B2 => n3992
                           , ZN => n2081);
   U191 : OAI22_X1 port map( A1 => n6025, A2 => n3993, B1 => n4027, B2 => n3992
                           , ZN => n2080);
   U192 : OAI22_X1 port map( A1 => n5752, A2 => n3993, B1 => n4028, B2 => n3994
                           , ZN => n2079);
   U193 : OAI22_X1 port map( A1 => n6026, A2 => n3993, B1 => n4030, B2 => n3994
                           , ZN => n2078);
   U194 : OAI22_X1 port map( A1 => n6027, A2 => n3993, B1 => n4171, B2 => n3994
                           , ZN => n2077);
   U195 : OAI22_X1 port map( A1 => n6520, A2 => n3993, B1 => n4172, B2 => n3994
                           , ZN => n2076);
   U196 : OAI22_X1 port map( A1 => n6521, A2 => n3993, B1 => n4031, B2 => n3994
                           , ZN => n2075);
   U197 : OAI22_X1 port map( A1 => n6028, A2 => n3993, B1 => n4032, B2 => n3994
                           , ZN => n2074);
   U198 : OAI22_X1 port map( A1 => n6522, A2 => n3993, B1 => n4175, B2 => n3994
                           , ZN => n2073);
   U199 : OAI22_X1 port map( A1 => n5753, A2 => n3993, B1 => n4033, B2 => n3994
                           , ZN => n2072);
   U200 : OAI22_X1 port map( A1 => n6523, A2 => n3993, B1 => n4035, B2 => n3994
                           , ZN => n2071);
   U201 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n4010);
   U202 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n4010, ZN => n4122);
   U203 : NAND2_X1 port map( A1 => n4012, A2 => n4122, ZN => n3997);
   U204 : CLKBUF_X1 port map( A => n3997, Z => n3995);
   U205 : OAI22_X1 port map( A1 => n6524, A2 => n3996, B1 => n4107, B2 => n3995
                           , ZN => n2070);
   U206 : OAI22_X1 port map( A1 => n5754, A2 => n3996, B1 => n4081, B2 => n3995
                           , ZN => n2069);
   U207 : OAI22_X1 port map( A1 => n6029, A2 => n3996, B1 => n4082, B2 => n3995
                           , ZN => n2068);
   U208 : OAI22_X1 port map( A1 => n6030, A2 => n3996, B1 => n4083, B2 => n3995
                           , ZN => n2067);
   U209 : OAI22_X1 port map( A1 => n5755, A2 => n3996, B1 => n4084, B2 => n3995
                           , ZN => n2066);
   U210 : OAI22_X1 port map( A1 => n6031, A2 => n3996, B1 => n4085, B2 => n3995
                           , ZN => n2065);
   U211 : OAI22_X1 port map( A1 => n6032, A2 => n3996, B1 => n4086, B2 => n3995
                           , ZN => n2064);
   U212 : OAI22_X1 port map( A1 => n6525, A2 => n3996, B1 => n4087, B2 => n3995
                           , ZN => n2063);
   U213 : OAI22_X1 port map( A1 => n5756, A2 => n3996, B1 => n4013, B2 => n3995
                           , ZN => n2062);
   U214 : OAI22_X1 port map( A1 => n6033, A2 => n3996, B1 => n4014, B2 => n3995
                           , ZN => n2061);
   U215 : OAI22_X1 port map( A1 => n5757, A2 => n3996, B1 => n4015, B2 => n3995
                           , ZN => n2060);
   U216 : OAI22_X1 port map( A1 => n5758, A2 => n3996, B1 => n4016, B2 => n3997
                           , ZN => n2059);
   U217 : OAI22_X1 port map( A1 => n5759, A2 => n3996, B1 => n4017, B2 => n3997
                           , ZN => n2058);
   U218 : OAI22_X1 port map( A1 => n5760, A2 => n3996, B1 => n4018, B2 => n3997
                           , ZN => n2057);
   U219 : OAI22_X1 port map( A1 => n5761, A2 => n3996, B1 => n4158, B2 => n3997
                           , ZN => n2056);
   U220 : OAI22_X1 port map( A1 => n6034, A2 => n3996, B1 => n4019, B2 => n3997
                           , ZN => n2055);
   U221 : OAI22_X1 port map( A1 => n6281, A2 => n3996, B1 => n4020, B2 => n3997
                           , ZN => n2054);
   U222 : OAI22_X1 port map( A1 => n6526, A2 => n3996, B1 => n4021, B2 => n3997
                           , ZN => n2053);
   U223 : OAI22_X1 port map( A1 => n5762, A2 => n3996, B1 => n4022, B2 => n3997
                           , ZN => n2052);
   U224 : OAI22_X1 port map( A1 => n5763, A2 => n3996, B1 => n4023, B2 => n3997
                           , ZN => n2051);
   U225 : OAI22_X1 port map( A1 => n6035, A2 => n3996, B1 => n4024, B2 => n3995
                           , ZN => n2050);
   U226 : OAI22_X1 port map( A1 => n6282, A2 => n3996, B1 => n4025, B2 => n3995
                           , ZN => n2049);
   U227 : OAI22_X1 port map( A1 => n5764, A2 => n3996, B1 => n4027, B2 => n3995
                           , ZN => n2048);
   U228 : OAI22_X1 port map( A1 => n5765, A2 => n3996, B1 => n4028, B2 => n3997
                           , ZN => n2047);
   U229 : OAI22_X1 port map( A1 => n6527, A2 => n3996, B1 => n4030, B2 => n3997
                           , ZN => n2046);
   U230 : OAI22_X1 port map( A1 => n5766, A2 => n3996, B1 => n4171, B2 => n3997
                           , ZN => n2045);
   U231 : OAI22_X1 port map( A1 => n6036, A2 => n3996, B1 => n4172, B2 => n3997
                           , ZN => n2044);
   U232 : OAI22_X1 port map( A1 => n5767, A2 => n3996, B1 => n4031, B2 => n3997
                           , ZN => n2043);
   U233 : OAI22_X1 port map( A1 => n6037, A2 => n3996, B1 => n4032, B2 => n3997
                           , ZN => n2042);
   U234 : OAI22_X1 port map( A1 => n6038, A2 => n3996, B1 => n4175, B2 => n3997
                           , ZN => n2041);
   U235 : OAI22_X1 port map( A1 => n5768, A2 => n3996, B1 => n4033, B2 => n3997
                           , ZN => n2040);
   U236 : OAI22_X1 port map( A1 => n5769, A2 => n3996, B1 => n4035, B2 => n3997
                           , ZN => n2039);
   U237 : INV_X1 port map( A => ADD_WR(2), ZN => n4011);
   U238 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n4011, ZN 
                           => n4127);
   U239 : NAND2_X1 port map( A1 => n4012, A2 => n4127, ZN => n4000);
   U240 : CLKBUF_X1 port map( A => n4000, Z => n3998);
   U241 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n3998, ZN => n3999);
   U242 : OAI22_X1 port map( A1 => n6528, A2 => n3999, B1 => n4107, B2 => n3998
                           , ZN => n2038);
   U243 : OAI22_X1 port map( A1 => n5770, A2 => n3999, B1 => n4081, B2 => n3998
                           , ZN => n2037);
   U244 : OAI22_X1 port map( A1 => n6283, A2 => n3999, B1 => n4082, B2 => n3998
                           , ZN => n2036);
   U245 : OAI22_X1 port map( A1 => n6529, A2 => n3999, B1 => n4083, B2 => n3998
                           , ZN => n2035);
   U246 : OAI22_X1 port map( A1 => n6284, A2 => n3999, B1 => n4084, B2 => n3998
                           , ZN => n2034);
   U247 : OAI22_X1 port map( A1 => n6285, A2 => n3999, B1 => n4085, B2 => n3998
                           , ZN => n2033);
   U248 : OAI22_X1 port map( A1 => n6286, A2 => n3999, B1 => n4086, B2 => n3998
                           , ZN => n2032);
   U249 : OAI22_X1 port map( A1 => n6530, A2 => n3999, B1 => n4087, B2 => n3998
                           , ZN => n2031);
   U250 : OAI22_X1 port map( A1 => n6287, A2 => n3999, B1 => n4013, B2 => n3998
                           , ZN => n2030);
   U251 : OAI22_X1 port map( A1 => n6531, A2 => n3999, B1 => n4014, B2 => n3998
                           , ZN => n2029);
   U252 : OAI22_X1 port map( A1 => n5771, A2 => n3999, B1 => n4015, B2 => n3998
                           , ZN => n2028);
   U253 : OAI22_X1 port map( A1 => n6288, A2 => n3999, B1 => n4016, B2 => n4000
                           , ZN => n2027);
   U254 : OAI22_X1 port map( A1 => n6532, A2 => n3999, B1 => n4017, B2 => n4000
                           , ZN => n2026);
   U255 : OAI22_X1 port map( A1 => n6289, A2 => n3999, B1 => n4018, B2 => n4000
                           , ZN => n2025);
   U256 : OAI22_X1 port map( A1 => n6533, A2 => n3999, B1 => n4158, B2 => n4000
                           , ZN => n2024);
   U257 : CLKBUF_X1 port map( A => n3999, Z => n4001);
   U258 : OAI22_X1 port map( A1 => n6290, A2 => n4001, B1 => n4019, B2 => n4000
                           , ZN => n2023);
   U259 : OAI22_X1 port map( A1 => n6534, A2 => n3999, B1 => n4020, B2 => n4000
                           , ZN => n2022);
   U260 : OAI22_X1 port map( A1 => n6291, A2 => n3999, B1 => n4021, B2 => n4000
                           , ZN => n2021);
   U261 : OAI22_X1 port map( A1 => n6292, A2 => n3999, B1 => n4022, B2 => n4000
                           , ZN => n2020);
   U262 : OAI22_X1 port map( A1 => n6535, A2 => n3999, B1 => n4023, B2 => n4000
                           , ZN => n2019);
   U263 : OAI22_X1 port map( A1 => n5772, A2 => n3999, B1 => n4024, B2 => n3998
                           , ZN => n2018);
   U264 : OAI22_X1 port map( A1 => n6536, A2 => n3999, B1 => n4025, B2 => n3998
                           , ZN => n2017);
   U265 : OAI22_X1 port map( A1 => n6293, A2 => n3999, B1 => n4027, B2 => n3998
                           , ZN => n2016);
   U266 : OAI22_X1 port map( A1 => n6294, A2 => n3999, B1 => n4028, B2 => n4000
                           , ZN => n2015);
   U267 : OAI22_X1 port map( A1 => n6295, A2 => n4001, B1 => n4030, B2 => n4000
                           , ZN => n2014);
   U268 : OAI22_X1 port map( A1 => n6296, A2 => n4001, B1 => n4171, B2 => n4000
                           , ZN => n2013);
   U269 : OAI22_X1 port map( A1 => n5773, A2 => n4001, B1 => n4172, B2 => n4000
                           , ZN => n2012);
   U270 : OAI22_X1 port map( A1 => n6537, A2 => n4001, B1 => n4031, B2 => n4000
                           , ZN => n2011);
   U271 : OAI22_X1 port map( A1 => n6538, A2 => n4001, B1 => n4032, B2 => n4000
                           , ZN => n2010);
   U272 : OAI22_X1 port map( A1 => n6039, A2 => n4001, B1 => n4175, B2 => n4000
                           , ZN => n2009);
   U273 : OAI22_X1 port map( A1 => n5774, A2 => n4001, B1 => n4033, B2 => n4000
                           , ZN => n2008);
   U274 : OAI22_X1 port map( A1 => n6297, A2 => n4001, B1 => n4035, B2 => n4000
                           , ZN => n2007);
   U275 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n4002, A3 => n4011, ZN => 
                           n4132);
   U276 : NAND2_X1 port map( A1 => n4012, A2 => n4132, ZN => n4005);
   U277 : OAI22_X1 port map( A1 => n5775, A2 => n4004, B1 => n4107, B2 => n4003
                           , ZN => n2006);
   U278 : OAI22_X1 port map( A1 => n6539, A2 => n4004, B1 => n4081, B2 => n4003
                           , ZN => n2005);
   U279 : OAI22_X1 port map( A1 => n5776, A2 => n4004, B1 => n4082, B2 => n4003
                           , ZN => n2004);
   U280 : OAI22_X1 port map( A1 => n6040, A2 => n4004, B1 => n4083, B2 => n4003
                           , ZN => n2003);
   U281 : OAI22_X1 port map( A1 => n6298, A2 => n4004, B1 => n4084, B2 => n4003
                           , ZN => n2002);
   U282 : OAI22_X1 port map( A1 => n6299, A2 => n4004, B1 => n4085, B2 => n4003
                           , ZN => n2001);
   U283 : OAI22_X1 port map( A1 => n5777, A2 => n4004, B1 => n4086, B2 => n4003
                           , ZN => n2000);
   U284 : OAI22_X1 port map( A1 => n6300, A2 => n4004, B1 => n4087, B2 => n4003
                           , ZN => n1999);
   U285 : OAI22_X1 port map( A1 => n6540, A2 => n4004, B1 => n4013, B2 => n4003
                           , ZN => n1998);
   U286 : OAI22_X1 port map( A1 => n6301, A2 => n4004, B1 => n4014, B2 => n4003
                           , ZN => n1997);
   U287 : OAI22_X1 port map( A1 => n6302, A2 => n4004, B1 => n4015, B2 => n4003
                           , ZN => n1996);
   U288 : OAI22_X1 port map( A1 => n6303, A2 => n4004, B1 => n4016, B2 => n4005
                           , ZN => n1995);
   U289 : OAI22_X1 port map( A1 => n6541, A2 => n4004, B1 => n4017, B2 => n4005
                           , ZN => n1994);
   U290 : OAI22_X1 port map( A1 => n6041, A2 => n4004, B1 => n4018, B2 => n4005
                           , ZN => n1993);
   U291 : OAI22_X1 port map( A1 => n6304, A2 => n4004, B1 => n4158, B2 => n4005
                           , ZN => n1992);
   U292 : OAI22_X1 port map( A1 => n6305, A2 => n4004, B1 => n4019, B2 => n4005
                           , ZN => n1991);
   U293 : OAI22_X1 port map( A1 => n6042, A2 => n4004, B1 => n4020, B2 => n4005
                           , ZN => n1990);
   U294 : OAI22_X1 port map( A1 => n5778, A2 => n4004, B1 => n4021, B2 => n4005
                           , ZN => n1989);
   U295 : OAI22_X1 port map( A1 => n6542, A2 => n4004, B1 => n4022, B2 => n4005
                           , ZN => n1988);
   U296 : OAI22_X1 port map( A1 => n6543, A2 => n4004, B1 => n4023, B2 => n4005
                           , ZN => n1987);
   U297 : OAI22_X1 port map( A1 => n6306, A2 => n4004, B1 => n4024, B2 => n4003
                           , ZN => n1986);
   U298 : OAI22_X1 port map( A1 => n6544, A2 => n4004, B1 => n4025, B2 => n4003
                           , ZN => n1985);
   U299 : OAI22_X1 port map( A1 => n6307, A2 => n4004, B1 => n4027, B2 => n4003
                           , ZN => n1984);
   U300 : OAI22_X1 port map( A1 => n6545, A2 => n4004, B1 => n4028, B2 => n4005
                           , ZN => n1983);
   U301 : OAI22_X1 port map( A1 => n6546, A2 => n4004, B1 => n4030, B2 => n4005
                           , ZN => n1982);
   U302 : OAI22_X1 port map( A1 => n6043, A2 => n4004, B1 => n4171, B2 => n4005
                           , ZN => n1981);
   U303 : OAI22_X1 port map( A1 => n6308, A2 => n4004, B1 => n4172, B2 => n4005
                           , ZN => n1980);
   U304 : OAI22_X1 port map( A1 => n6309, A2 => n4004, B1 => n4031, B2 => n4005
                           , ZN => n1979);
   U305 : OAI22_X1 port map( A1 => n6310, A2 => n4004, B1 => n4032, B2 => n4005
                           , ZN => n1978);
   U306 : OAI22_X1 port map( A1 => n6311, A2 => n4004, B1 => n4175, B2 => n4005
                           , ZN => n1977);
   U307 : OAI22_X1 port map( A1 => n6547, A2 => n4004, B1 => n4033, B2 => n4005
                           , ZN => n1976);
   U308 : OAI22_X1 port map( A1 => n6548, A2 => n4004, B1 => n4035, B2 => n4005
                           , ZN => n1975);
   U309 : NOR2_X1 port map( A1 => n4011, A2 => n4006, ZN => n4137);
   U310 : NAND2_X1 port map( A1 => n4012, A2 => n4137, ZN => n4009);
   U311 : CLKBUF_X1 port map( A => n4009, Z => n4007);
   U312 : OAI22_X1 port map( A1 => n6312, A2 => n4008, B1 => n4107, B2 => n4007
                           , ZN => n1974);
   U313 : OAI22_X1 port map( A1 => n6044, A2 => n4008, B1 => n4081, B2 => n4007
                           , ZN => n1973);
   U314 : OAI22_X1 port map( A1 => n6549, A2 => n4008, B1 => n4082, B2 => n4007
                           , ZN => n1972);
   U315 : OAI22_X1 port map( A1 => n6550, A2 => n4008, B1 => n4083, B2 => n4007
                           , ZN => n1971);
   U316 : OAI22_X1 port map( A1 => n5779, A2 => n4008, B1 => n4084, B2 => n4007
                           , ZN => n1970);
   U317 : OAI22_X1 port map( A1 => n5780, A2 => n4008, B1 => n4085, B2 => n4007
                           , ZN => n1969);
   U318 : OAI22_X1 port map( A1 => n6551, A2 => n4008, B1 => n4086, B2 => n4007
                           , ZN => n1968);
   U319 : OAI22_X1 port map( A1 => n5781, A2 => n4008, B1 => n4087, B2 => n4007
                           , ZN => n1967);
   U320 : OAI22_X1 port map( A1 => n5782, A2 => n4008, B1 => n4013, B2 => n4007
                           , ZN => n1966);
   U321 : OAI22_X1 port map( A1 => n6045, A2 => n4008, B1 => n4014, B2 => n4007
                           , ZN => n1965);
   U322 : OAI22_X1 port map( A1 => n6552, A2 => n4008, B1 => n4015, B2 => n4007
                           , ZN => n1964);
   U323 : OAI22_X1 port map( A1 => n6046, A2 => n4008, B1 => n4016, B2 => n4009
                           , ZN => n1963);
   U324 : OAI22_X1 port map( A1 => n5783, A2 => n4008, B1 => n4017, B2 => n4009
                           , ZN => n1962);
   U325 : OAI22_X1 port map( A1 => n6553, A2 => n4008, B1 => n4018, B2 => n4009
                           , ZN => n1961);
   U326 : OAI22_X1 port map( A1 => n6047, A2 => n4008, B1 => n4158, B2 => n4009
                           , ZN => n1960);
   U327 : OAI22_X1 port map( A1 => n5784, A2 => n4008, B1 => n4019, B2 => n4009
                           , ZN => n1959);
   U328 : OAI22_X1 port map( A1 => n6313, A2 => n4008, B1 => n4020, B2 => n4009
                           , ZN => n1958);
   U329 : OAI22_X1 port map( A1 => n6048, A2 => n4008, B1 => n4021, B2 => n4009
                           , ZN => n1957);
   U330 : OAI22_X1 port map( A1 => n6049, A2 => n4008, B1 => n4022, B2 => n4009
                           , ZN => n1956);
   U331 : OAI22_X1 port map( A1 => n6314, A2 => n4008, B1 => n4023, B2 => n4009
                           , ZN => n1955);
   U332 : OAI22_X1 port map( A1 => n6554, A2 => n4008, B1 => n4024, B2 => n4007
                           , ZN => n1954);
   U333 : OAI22_X1 port map( A1 => n6050, A2 => n4008, B1 => n4025, B2 => n4007
                           , ZN => n1953);
   U334 : OAI22_X1 port map( A1 => n6051, A2 => n4008, B1 => n4027, B2 => n4007
                           , ZN => n1952);
   U335 : OAI22_X1 port map( A1 => n6555, A2 => n4008, B1 => n4028, B2 => n4009
                           , ZN => n1951);
   U336 : OAI22_X1 port map( A1 => n5785, A2 => n4008, B1 => n4030, B2 => n4009
                           , ZN => n1950);
   U337 : OAI22_X1 port map( A1 => n6556, A2 => n4008, B1 => n4171, B2 => n4009
                           , ZN => n1949);
   U338 : OAI22_X1 port map( A1 => n5786, A2 => n4008, B1 => n4172, B2 => n4009
                           , ZN => n1948);
   U339 : OAI22_X1 port map( A1 => n6052, A2 => n4008, B1 => n4031, B2 => n4009
                           , ZN => n1947);
   U340 : OAI22_X1 port map( A1 => n5787, A2 => n4008, B1 => n4032, B2 => n4009
                           , ZN => n1946);
   U341 : OAI22_X1 port map( A1 => n6315, A2 => n4008, B1 => n4175, B2 => n4009
                           , ZN => n1945);
   U342 : OAI22_X1 port map( A1 => n6557, A2 => n4008, B1 => n4033, B2 => n4009
                           , ZN => n1944);
   U343 : OAI22_X1 port map( A1 => n6053, A2 => n4008, B1 => n4035, B2 => n4009
                           , ZN => n1943);
   U344 : NOR2_X1 port map( A1 => n4011, A2 => n4010, ZN => n4143);
   U345 : NAND2_X1 port map( A1 => n4012, A2 => n4143, ZN => n4034);
   U346 : CLKBUF_X1 port map( A => n4034, Z => n4026);
   U347 : OAI22_X1 port map( A1 => n6054, A2 => n4029, B1 => n4107, B2 => n4026
                           , ZN => n1942);
   U348 : OAI22_X1 port map( A1 => n5788, A2 => n4029, B1 => n4081, B2 => n4026
                           , ZN => n1941);
   U349 : OAI22_X1 port map( A1 => n5789, A2 => n4029, B1 => n4082, B2 => n4026
                           , ZN => n1940);
   U350 : OAI22_X1 port map( A1 => n5790, A2 => n4029, B1 => n4083, B2 => n4026
                           , ZN => n1939);
   U351 : OAI22_X1 port map( A1 => n6055, A2 => n4029, B1 => n4084, B2 => n4026
                           , ZN => n1938);
   U352 : OAI22_X1 port map( A1 => n6056, A2 => n4029, B1 => n4085, B2 => n4026
                           , ZN => n1937);
   U353 : OAI22_X1 port map( A1 => n5791, A2 => n4029, B1 => n4086, B2 => n4026
                           , ZN => n1936);
   U354 : OAI22_X1 port map( A1 => n6057, A2 => n4029, B1 => n4087, B2 => n4026
                           , ZN => n1935);
   U355 : OAI22_X1 port map( A1 => n6058, A2 => n4029, B1 => n4013, B2 => n4026
                           , ZN => n1934);
   U356 : OAI22_X1 port map( A1 => n5792, A2 => n4029, B1 => n4014, B2 => n4026
                           , ZN => n1933);
   U357 : OAI22_X1 port map( A1 => n6059, A2 => n4029, B1 => n4015, B2 => n4026
                           , ZN => n1932);
   U358 : OAI22_X1 port map( A1 => n6060, A2 => n4029, B1 => n4016, B2 => n4034
                           , ZN => n1931);
   U359 : OAI22_X1 port map( A1 => n6061, A2 => n4029, B1 => n4017, B2 => n4034
                           , ZN => n1930);
   U360 : OAI22_X1 port map( A1 => n5793, A2 => n4029, B1 => n4018, B2 => n4034
                           , ZN => n1929);
   U361 : OAI22_X1 port map( A1 => n6062, A2 => n4029, B1 => n4158, B2 => n4034
                           , ZN => n1928);
   U362 : OAI22_X1 port map( A1 => n6063, A2 => n4029, B1 => n4019, B2 => n4034
                           , ZN => n1927);
   U363 : OAI22_X1 port map( A1 => n5794, A2 => n4029, B1 => n4020, B2 => n4034
                           , ZN => n1926);
   U364 : OAI22_X1 port map( A1 => n5795, A2 => n4029, B1 => n4021, B2 => n4034
                           , ZN => n1925);
   U365 : OAI22_X1 port map( A1 => n6064, A2 => n4029, B1 => n4022, B2 => n4034
                           , ZN => n1924);
   U366 : OAI22_X1 port map( A1 => n5796, A2 => n4029, B1 => n4023, B2 => n4034
                           , ZN => n1923);
   U367 : OAI22_X1 port map( A1 => n5797, A2 => n4029, B1 => n4024, B2 => n4026
                           , ZN => n1922);
   U368 : OAI22_X1 port map( A1 => n5798, A2 => n4029, B1 => n4025, B2 => n4026
                           , ZN => n1921);
   U369 : OAI22_X1 port map( A1 => n6065, A2 => n4029, B1 => n4027, B2 => n4026
                           , ZN => n1920);
   U370 : OAI22_X1 port map( A1 => n6066, A2 => n4029, B1 => n4028, B2 => n4034
                           , ZN => n1919);
   U371 : OAI22_X1 port map( A1 => n5799, A2 => n4029, B1 => n4030, B2 => n4034
                           , ZN => n1918);
   U372 : OAI22_X1 port map( A1 => n5800, A2 => n4029, B1 => n4171, B2 => n4034
                           , ZN => n1917);
   U373 : OAI22_X1 port map( A1 => n6067, A2 => n4029, B1 => n4172, B2 => n4034
                           , ZN => n1916);
   U374 : OAI22_X1 port map( A1 => n6068, A2 => n4029, B1 => n4031, B2 => n4034
                           , ZN => n1915);
   U375 : OAI22_X1 port map( A1 => n5801, A2 => n4029, B1 => n4032, B2 => n4034
                           , ZN => n1914);
   U376 : OAI22_X1 port map( A1 => n6069, A2 => n4029, B1 => n4175, B2 => n4034
                           , ZN => n1913);
   U377 : OAI22_X1 port map( A1 => n6070, A2 => n4029, B1 => n4033, B2 => n4034
                           , ZN => n1912);
   U378 : OAI22_X1 port map( A1 => n6071, A2 => n4029, B1 => n4035, B2 => n4034
                           , ZN => n1911);
   U379 : INV_X1 port map( A => ADD_WR(3), ZN => n4105);
   U380 : NOR2_X1 port map( A1 => n4105, A2 => n4036, ZN => n4060);
   U381 : NAND2_X1 port map( A1 => n4106, A2 => n4060, ZN => n4039);
   U382 : CLKBUF_X1 port map( A => n4039, Z => n4037);
   U383 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4037, ZN => n4038);
   U384 : OAI22_X1 port map( A1 => n6558, A2 => n4038, B1 => n4107, B2 => n4037
                           , ZN => n1910);
   U385 : OAI22_X1 port map( A1 => n6559, A2 => n4038, B1 => n4145, B2 => n4037
                           , ZN => n1909);
   U386 : OAI22_X1 port map( A1 => n6316, A2 => n4038, B1 => n4146, B2 => n4037
                           , ZN => n1908);
   U387 : OAI22_X1 port map( A1 => n6317, A2 => n4038, B1 => n4147, B2 => n4037
                           , ZN => n1907);
   U388 : OAI22_X1 port map( A1 => n6560, A2 => n4038, B1 => n4148, B2 => n4037
                           , ZN => n1906);
   U389 : OAI22_X1 port map( A1 => n6318, A2 => n4038, B1 => n4149, B2 => n4037
                           , ZN => n1905);
   U390 : OAI22_X1 port map( A1 => n6561, A2 => n4038, B1 => n4150, B2 => n4037
                           , ZN => n1904);
   U391 : OAI22_X1 port map( A1 => n6319, A2 => n4038, B1 => n4151, B2 => n4037
                           , ZN => n1903);
   U392 : OAI22_X1 port map( A1 => n6320, A2 => n4038, B1 => n4152, B2 => n4037
                           , ZN => n1902);
   U393 : OAI22_X1 port map( A1 => n6321, A2 => n4038, B1 => n4153, B2 => n4037
                           , ZN => n1901);
   U394 : OAI22_X1 port map( A1 => n6562, A2 => n4038, B1 => n4154, B2 => n4037
                           , ZN => n1900);
   U395 : OAI22_X1 port map( A1 => n6563, A2 => n4038, B1 => n4155, B2 => n4039
                           , ZN => n1899);
   U396 : OAI22_X1 port map( A1 => n6322, A2 => n4038, B1 => n4156, B2 => n4039
                           , ZN => n1898);
   U397 : OAI22_X1 port map( A1 => n6323, A2 => n4038, B1 => n4157, B2 => n4039
                           , ZN => n1897);
   U398 : OAI22_X1 port map( A1 => n6324, A2 => n4038, B1 => n4158, B2 => n4039
                           , ZN => n1896);
   U399 : OAI22_X1 port map( A1 => n6325, A2 => n4038, B1 => n4159, B2 => n4039
                           , ZN => n1895);
   U400 : OAI22_X1 port map( A1 => n6564, A2 => n4038, B1 => n4160, B2 => n4039
                           , ZN => n1894);
   U401 : CLKBUF_X1 port map( A => n4038, Z => n4040);
   U402 : OAI22_X1 port map( A1 => n6565, A2 => n4040, B1 => n4161, B2 => n4039
                           , ZN => n1893);
   U403 : OAI22_X1 port map( A1 => n6566, A2 => n4038, B1 => n4162, B2 => n4039
                           , ZN => n1892);
   U404 : OAI22_X1 port map( A1 => n6567, A2 => n4038, B1 => n4163, B2 => n4039
                           , ZN => n1891);
   U405 : OAI22_X1 port map( A1 => n6326, A2 => n4038, B1 => n4164, B2 => n4037
                           , ZN => n1890);
   U406 : OAI22_X1 port map( A1 => n6327, A2 => n4038, B1 => n4165, B2 => n4037
                           , ZN => n1889);
   U407 : OAI22_X1 port map( A1 => n6328, A2 => n4038, B1 => n4167, B2 => n4037
                           , ZN => n1888);
   U408 : OAI22_X1 port map( A1 => n6329, A2 => n4038, B1 => n4168, B2 => n4039
                           , ZN => n1887);
   U409 : OAI22_X1 port map( A1 => n6568, A2 => n4040, B1 => n4170, B2 => n4039
                           , ZN => n1886);
   U410 : OAI22_X1 port map( A1 => n6330, A2 => n4040, B1 => n4171, B2 => n4039
                           , ZN => n1885);
   U411 : OAI22_X1 port map( A1 => n6569, A2 => n4040, B1 => n4172, B2 => n4039
                           , ZN => n1884);
   U412 : OAI22_X1 port map( A1 => n6331, A2 => n4040, B1 => n4173, B2 => n4039
                           , ZN => n1883);
   U413 : OAI22_X1 port map( A1 => n6570, A2 => n4040, B1 => n4174, B2 => n4039
                           , ZN => n1882);
   U414 : OAI22_X1 port map( A1 => n6332, A2 => n4040, B1 => n4175, B2 => n4039
                           , ZN => n1881);
   U415 : OAI22_X1 port map( A1 => n6333, A2 => n4040, B1 => n4176, B2 => n4039
                           , ZN => n1880);
   U416 : OAI22_X1 port map( A1 => n6571, A2 => n4040, B1 => n4178, B2 => n4039
                           , ZN => n1879);
   U417 : NAND2_X1 port map( A1 => n4112, A2 => n4060, ZN => n4043);
   U418 : CLKBUF_X1 port map( A => n4043, Z => n4041);
   U419 : OAI22_X1 port map( A1 => n5802, A2 => n4042, B1 => n4107, B2 => n4041
                           , ZN => n1878);
   U420 : OAI22_X1 port map( A1 => n6572, A2 => n4042, B1 => n4145, B2 => n4041
                           , ZN => n1877);
   U421 : OAI22_X1 port map( A1 => n5803, A2 => n4042, B1 => n4146, B2 => n4041
                           , ZN => n1876);
   U422 : OAI22_X1 port map( A1 => n6072, A2 => n4042, B1 => n4147, B2 => n4041
                           , ZN => n1875);
   U423 : OAI22_X1 port map( A1 => n6073, A2 => n4042, B1 => n4148, B2 => n4041
                           , ZN => n1874);
   U424 : OAI22_X1 port map( A1 => n5804, A2 => n4042, B1 => n4149, B2 => n4041
                           , ZN => n1873);
   U425 : OAI22_X1 port map( A1 => n5805, A2 => n4042, B1 => n4150, B2 => n4041
                           , ZN => n1872);
   U426 : OAI22_X1 port map( A1 => n6074, A2 => n4042, B1 => n4151, B2 => n4041
                           , ZN => n1871);
   U427 : OAI22_X1 port map( A1 => n6075, A2 => n4042, B1 => n4152, B2 => n4041
                           , ZN => n1870);
   U428 : OAI22_X1 port map( A1 => n6334, A2 => n4042, B1 => n4153, B2 => n4041
                           , ZN => n1869);
   U429 : OAI22_X1 port map( A1 => n6573, A2 => n4042, B1 => n4154, B2 => n4041
                           , ZN => n1868);
   U430 : OAI22_X1 port map( A1 => n6574, A2 => n4042, B1 => n4155, B2 => n4043
                           , ZN => n1867);
   U431 : OAI22_X1 port map( A1 => n5806, A2 => n4042, B1 => n4156, B2 => n4043
                           , ZN => n1866);
   U432 : OAI22_X1 port map( A1 => n6575, A2 => n4042, B1 => n4157, B2 => n4043
                           , ZN => n1865);
   U433 : OAI22_X1 port map( A1 => n6335, A2 => n4042, B1 => n4158, B2 => n4043
                           , ZN => n1864);
   U434 : OAI22_X1 port map( A1 => n5807, A2 => n4042, B1 => n4159, B2 => n4043
                           , ZN => n1863);
   U435 : OAI22_X1 port map( A1 => n6076, A2 => n4042, B1 => n4160, B2 => n4043
                           , ZN => n1862);
   U436 : OAI22_X1 port map( A1 => n5808, A2 => n4042, B1 => n4161, B2 => n4043
                           , ZN => n1861);
   U437 : OAI22_X1 port map( A1 => n6336, A2 => n4042, B1 => n4162, B2 => n4043
                           , ZN => n1860);
   U438 : OAI22_X1 port map( A1 => n6077, A2 => n4042, B1 => n4163, B2 => n4043
                           , ZN => n1859);
   U439 : OAI22_X1 port map( A1 => n5809, A2 => n4042, B1 => n4164, B2 => n4041
                           , ZN => n1858);
   U440 : OAI22_X1 port map( A1 => n6576, A2 => n4042, B1 => n4165, B2 => n4041
                           , ZN => n1857);
   U441 : OAI22_X1 port map( A1 => n6577, A2 => n4042, B1 => n4167, B2 => n4041
                           , ZN => n1856);
   U442 : OAI22_X1 port map( A1 => n6578, A2 => n4042, B1 => n4168, B2 => n4043
                           , ZN => n1855);
   U443 : OAI22_X1 port map( A1 => n6579, A2 => n4042, B1 => n4170, B2 => n4043
                           , ZN => n1854);
   U444 : OAI22_X1 port map( A1 => n6580, A2 => n4042, B1 => n4171, B2 => n4043
                           , ZN => n1853);
   U445 : OAI22_X1 port map( A1 => n6337, A2 => n4042, B1 => n4172, B2 => n4043
                           , ZN => n1852);
   U446 : OAI22_X1 port map( A1 => n6581, A2 => n4042, B1 => n4173, B2 => n4043
                           , ZN => n1851);
   U447 : OAI22_X1 port map( A1 => n6338, A2 => n4042, B1 => n4174, B2 => n4043
                           , ZN => n1850);
   U448 : OAI22_X1 port map( A1 => n6582, A2 => n4042, B1 => n4175, B2 => n4043
                           , ZN => n1849);
   U449 : OAI22_X1 port map( A1 => n5810, A2 => n4042, B1 => n4176, B2 => n4043
                           , ZN => n1848);
   U450 : OAI22_X1 port map( A1 => n5811, A2 => n4042, B1 => n4178, B2 => n4043
                           , ZN => n1847);
   U451 : NAND2_X1 port map( A1 => n4117, A2 => n4060, ZN => n4046);
   U452 : CLKBUF_X1 port map( A => n4046, Z => n4044);
   U453 : OAI22_X1 port map( A1 => n5812, A2 => n4045, B1 => n4107, B2 => n4044
                           , ZN => n1846);
   U454 : OAI22_X1 port map( A1 => n6078, A2 => n4045, B1 => n4145, B2 => n4044
                           , ZN => n1845);
   U455 : OAI22_X1 port map( A1 => n5813, A2 => n4045, B1 => n4146, B2 => n4044
                           , ZN => n1844);
   U456 : OAI22_X1 port map( A1 => n5814, A2 => n4045, B1 => n4147, B2 => n4044
                           , ZN => n1843);
   U457 : OAI22_X1 port map( A1 => n6339, A2 => n4045, B1 => n4148, B2 => n4044
                           , ZN => n1842);
   U458 : OAI22_X1 port map( A1 => n5815, A2 => n4045, B1 => n4149, B2 => n4044
                           , ZN => n1841);
   U459 : OAI22_X1 port map( A1 => n5816, A2 => n4045, B1 => n4150, B2 => n4044
                           , ZN => n1840);
   U460 : OAI22_X1 port map( A1 => n6079, A2 => n4045, B1 => n4151, B2 => n4044
                           , ZN => n1839);
   U461 : OAI22_X1 port map( A1 => n6340, A2 => n4045, B1 => n4152, B2 => n4044
                           , ZN => n1838);
   U462 : OAI22_X1 port map( A1 => n5817, A2 => n4045, B1 => n4153, B2 => n4044
                           , ZN => n1837);
   U463 : OAI22_X1 port map( A1 => n6080, A2 => n4045, B1 => n4154, B2 => n4044
                           , ZN => n1836);
   U464 : OAI22_X1 port map( A1 => n5818, A2 => n4045, B1 => n4155, B2 => n4046
                           , ZN => n1835);
   U465 : OAI22_X1 port map( A1 => n5819, A2 => n4045, B1 => n4156, B2 => n4046
                           , ZN => n1834);
   U466 : OAI22_X1 port map( A1 => n5820, A2 => n4045, B1 => n4157, B2 => n4046
                           , ZN => n1833);
   U467 : OAI22_X1 port map( A1 => n6081, A2 => n4045, B1 => n4158, B2 => n4046
                           , ZN => n1832);
   U468 : OAI22_X1 port map( A1 => n6082, A2 => n4045, B1 => n4159, B2 => n4046
                           , ZN => n1831);
   U469 : OAI22_X1 port map( A1 => n5821, A2 => n4045, B1 => n4160, B2 => n4046
                           , ZN => n1830);
   U470 : OAI22_X1 port map( A1 => n6083, A2 => n4045, B1 => n4161, B2 => n4046
                           , ZN => n1829);
   U471 : OAI22_X1 port map( A1 => n5822, A2 => n4045, B1 => n4162, B2 => n4046
                           , ZN => n1828);
   U472 : OAI22_X1 port map( A1 => n5823, A2 => n4045, B1 => n4163, B2 => n4046
                           , ZN => n1827);
   U473 : OAI22_X1 port map( A1 => n6084, A2 => n4045, B1 => n4164, B2 => n4044
                           , ZN => n1826);
   U474 : OAI22_X1 port map( A1 => n6085, A2 => n4045, B1 => n4165, B2 => n4044
                           , ZN => n1825);
   U475 : OAI22_X1 port map( A1 => n6086, A2 => n4045, B1 => n4167, B2 => n4044
                           , ZN => n1824);
   U476 : OAI22_X1 port map( A1 => n5824, A2 => n4045, B1 => n4168, B2 => n4046
                           , ZN => n1823);
   U477 : OAI22_X1 port map( A1 => n5825, A2 => n4045, B1 => n4170, B2 => n4046
                           , ZN => n1822);
   U478 : OAI22_X1 port map( A1 => n5826, A2 => n4045, B1 => n4171, B2 => n4046
                           , ZN => n1821);
   U479 : OAI22_X1 port map( A1 => n5827, A2 => n4045, B1 => n4172, B2 => n4046
                           , ZN => n1820);
   U480 : OAI22_X1 port map( A1 => n5828, A2 => n4045, B1 => n4173, B2 => n4046
                           , ZN => n1819);
   U481 : OAI22_X1 port map( A1 => n5829, A2 => n4045, B1 => n4174, B2 => n4046
                           , ZN => n1818);
   U482 : OAI22_X1 port map( A1 => n6087, A2 => n4045, B1 => n4175, B2 => n4046
                           , ZN => n1817);
   U483 : OAI22_X1 port map( A1 => n6583, A2 => n4045, B1 => n4176, B2 => n4046
                           , ZN => n1816);
   U484 : OAI22_X1 port map( A1 => n5830, A2 => n4045, B1 => n4178, B2 => n4046
                           , ZN => n1815);
   U485 : NAND2_X1 port map( A1 => n4122, A2 => n4060, ZN => n4049);
   U486 : CLKBUF_X1 port map( A => n4049, Z => n4047);
   U487 : OAI22_X1 port map( A1 => n6341, A2 => n4048, B1 => n4107, B2 => n4047
                           , ZN => n1814);
   U488 : OAI22_X1 port map( A1 => n5831, A2 => n4048, B1 => n4145, B2 => n4047
                           , ZN => n1813);
   U489 : OAI22_X1 port map( A1 => n6088, A2 => n4048, B1 => n4146, B2 => n4047
                           , ZN => n1812);
   U490 : OAI22_X1 port map( A1 => n6089, A2 => n4048, B1 => n4147, B2 => n4047
                           , ZN => n1811);
   U491 : OAI22_X1 port map( A1 => n6090, A2 => n4048, B1 => n4148, B2 => n4047
                           , ZN => n1810);
   U492 : OAI22_X1 port map( A1 => n6584, A2 => n4048, B1 => n4149, B2 => n4047
                           , ZN => n1809);
   U493 : OAI22_X1 port map( A1 => n6091, A2 => n4048, B1 => n4150, B2 => n4047
                           , ZN => n1808);
   U494 : OAI22_X1 port map( A1 => n6092, A2 => n4048, B1 => n4151, B2 => n4047
                           , ZN => n1807);
   U495 : OAI22_X1 port map( A1 => n6093, A2 => n4048, B1 => n4152, B2 => n4047
                           , ZN => n1806);
   U496 : OAI22_X1 port map( A1 => n6585, A2 => n4048, B1 => n4153, B2 => n4047
                           , ZN => n1805);
   U497 : OAI22_X1 port map( A1 => n5832, A2 => n4048, B1 => n4154, B2 => n4047
                           , ZN => n1804);
   U498 : OAI22_X1 port map( A1 => n6094, A2 => n4048, B1 => n4155, B2 => n4049
                           , ZN => n1803);
   U499 : OAI22_X1 port map( A1 => n6586, A2 => n4048, B1 => n4156, B2 => n4049
                           , ZN => n1802);
   U500 : OAI22_X1 port map( A1 => n5833, A2 => n4048, B1 => n4157, B2 => n4049
                           , ZN => n1801);
   U501 : OAI22_X1 port map( A1 => n6095, A2 => n4048, B1 => n4158, B2 => n4049
                           , ZN => n1800);
   U502 : OAI22_X1 port map( A1 => n6587, A2 => n4048, B1 => n4159, B2 => n4049
                           , ZN => n1799);
   U503 : OAI22_X1 port map( A1 => n5834, A2 => n4048, B1 => n4160, B2 => n4049
                           , ZN => n1798);
   U504 : OAI22_X1 port map( A1 => n6342, A2 => n4048, B1 => n4161, B2 => n4049
                           , ZN => n1797);
   U505 : OAI22_X1 port map( A1 => n5835, A2 => n4048, B1 => n4162, B2 => n4049
                           , ZN => n1796);
   U506 : OAI22_X1 port map( A1 => n6096, A2 => n4048, B1 => n4163, B2 => n4049
                           , ZN => n1795);
   U507 : OAI22_X1 port map( A1 => n6343, A2 => n4048, B1 => n4164, B2 => n4047
                           , ZN => n1794);
   U508 : OAI22_X1 port map( A1 => n5836, A2 => n4048, B1 => n4165, B2 => n4047
                           , ZN => n1793);
   U509 : OAI22_X1 port map( A1 => n5837, A2 => n4048, B1 => n4167, B2 => n4047
                           , ZN => n1792);
   U510 : OAI22_X1 port map( A1 => n5838, A2 => n4048, B1 => n4168, B2 => n4049
                           , ZN => n1791);
   U511 : OAI22_X1 port map( A1 => n6097, A2 => n4048, B1 => n4170, B2 => n4049
                           , ZN => n1790);
   U512 : OAI22_X1 port map( A1 => n6098, A2 => n4048, B1 => n4171, B2 => n4049
                           , ZN => n1789);
   U513 : OAI22_X1 port map( A1 => n5839, A2 => n4048, B1 => n4172, B2 => n4049
                           , ZN => n1788);
   U514 : OAI22_X1 port map( A1 => n6099, A2 => n4048, B1 => n4173, B2 => n4049
                           , ZN => n1787);
   U515 : OAI22_X1 port map( A1 => n6100, A2 => n4048, B1 => n4174, B2 => n4049
                           , ZN => n1786);
   U516 : OAI22_X1 port map( A1 => n5840, A2 => n4048, B1 => n4175, B2 => n4049
                           , ZN => n1785);
   U517 : OAI22_X1 port map( A1 => n5841, A2 => n4048, B1 => n4176, B2 => n4049
                           , ZN => n1784);
   U518 : OAI22_X1 port map( A1 => n6588, A2 => n4048, B1 => n4178, B2 => n4049
                           , ZN => n1783);
   U519 : NAND2_X1 port map( A1 => n4127, A2 => n4060, ZN => n4052);
   U520 : CLKBUF_X1 port map( A => n4052, Z => n4050);
   U521 : OAI22_X1 port map( A1 => n6589, A2 => n4051, B1 => n4107, B2 => n4050
                           , ZN => n1782);
   U522 : OAI22_X1 port map( A1 => n5842, A2 => n4051, B1 => n4145, B2 => n4050
                           , ZN => n1781);
   U523 : OAI22_X1 port map( A1 => n6590, A2 => n4051, B1 => n4146, B2 => n4050
                           , ZN => n1780);
   U524 : OAI22_X1 port map( A1 => n6344, A2 => n4051, B1 => n4147, B2 => n4050
                           , ZN => n1779);
   U525 : OAI22_X1 port map( A1 => n6345, A2 => n4051, B1 => n4148, B2 => n4050
                           , ZN => n1778);
   U526 : OAI22_X1 port map( A1 => n6591, A2 => n4051, B1 => n4149, B2 => n4050
                           , ZN => n1777);
   U527 : OAI22_X1 port map( A1 => n6346, A2 => n4051, B1 => n4150, B2 => n4050
                           , ZN => n1776);
   U528 : OAI22_X1 port map( A1 => n6592, A2 => n4051, B1 => n4151, B2 => n4050
                           , ZN => n1775);
   U529 : OAI22_X1 port map( A1 => n6347, A2 => n4051, B1 => n4152, B2 => n4050
                           , ZN => n1774);
   U530 : OAI22_X1 port map( A1 => n6101, A2 => n4051, B1 => n4153, B2 => n4050
                           , ZN => n1773);
   U531 : OAI22_X1 port map( A1 => n6348, A2 => n4051, B1 => n4154, B2 => n4050
                           , ZN => n1772);
   U532 : OAI22_X1 port map( A1 => n5843, A2 => n4051, B1 => n4155, B2 => n4052
                           , ZN => n1771);
   U533 : OAI22_X1 port map( A1 => n6102, A2 => n4051, B1 => n4156, B2 => n4052
                           , ZN => n1770);
   U534 : OAI22_X1 port map( A1 => n5844, A2 => n4051, B1 => n4157, B2 => n4052
                           , ZN => n1769);
   U535 : OAI22_X1 port map( A1 => n6103, A2 => n4051, B1 => n4158, B2 => n4052
                           , ZN => n1768);
   U536 : OAI22_X1 port map( A1 => n6593, A2 => n4051, B1 => n4159, B2 => n4052
                           , ZN => n1767);
   U537 : OAI22_X1 port map( A1 => n6349, A2 => n4051, B1 => n4160, B2 => n4052
                           , ZN => n1766);
   U538 : OAI22_X1 port map( A1 => n5845, A2 => n4051, B1 => n4161, B2 => n4052
                           , ZN => n1765);
   U539 : OAI22_X1 port map( A1 => n6350, A2 => n4051, B1 => n4162, B2 => n4052
                           , ZN => n1764);
   U540 : OAI22_X1 port map( A1 => n6351, A2 => n4051, B1 => n4163, B2 => n4052
                           , ZN => n1763);
   U541 : OAI22_X1 port map( A1 => n6352, A2 => n4051, B1 => n4164, B2 => n4050
                           , ZN => n1762);
   U542 : OAI22_X1 port map( A1 => n6104, A2 => n4051, B1 => n4165, B2 => n4050
                           , ZN => n1761);
   U543 : OAI22_X1 port map( A1 => n5846, A2 => n4051, B1 => n4167, B2 => n4050
                           , ZN => n1760);
   U544 : OAI22_X1 port map( A1 => n5847, A2 => n4051, B1 => n4168, B2 => n4052
                           , ZN => n1759);
   U545 : OAI22_X1 port map( A1 => n6594, A2 => n4051, B1 => n4170, B2 => n4052
                           , ZN => n1758);
   U546 : OAI22_X1 port map( A1 => n6353, A2 => n4051, B1 => n4171, B2 => n4052
                           , ZN => n1757);
   U547 : OAI22_X1 port map( A1 => n6105, A2 => n4051, B1 => n4172, B2 => n4052
                           , ZN => n1756);
   U548 : OAI22_X1 port map( A1 => n6595, A2 => n4051, B1 => n4173, B2 => n4052
                           , ZN => n1755);
   U549 : OAI22_X1 port map( A1 => n6596, A2 => n4051, B1 => n4174, B2 => n4052
                           , ZN => n1754);
   U550 : OAI22_X1 port map( A1 => n5848, A2 => n4051, B1 => n4175, B2 => n4052
                           , ZN => n1753);
   U551 : OAI22_X1 port map( A1 => n6597, A2 => n4051, B1 => n4176, B2 => n4052
                           , ZN => n1752);
   U552 : OAI22_X1 port map( A1 => n6598, A2 => n4051, B1 => n4178, B2 => n4052
                           , ZN => n1751);
   U553 : NAND2_X1 port map( A1 => n4132, A2 => n4060, ZN => n4055);
   U554 : CLKBUF_X1 port map( A => n4055, Z => n4053);
   U555 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4053, ZN => n4054);
   U556 : OAI22_X1 port map( A1 => n6599, A2 => n4054, B1 => n4107, B2 => n4053
                           , ZN => n1750);
   U557 : OAI22_X1 port map( A1 => n6354, A2 => n4054, B1 => n4081, B2 => n4053
                           , ZN => n1749);
   U558 : OAI22_X1 port map( A1 => n6355, A2 => n4054, B1 => n4082, B2 => n4053
                           , ZN => n1748);
   U559 : OAI22_X1 port map( A1 => n6600, A2 => n4054, B1 => n4083, B2 => n4053
                           , ZN => n1747);
   U560 : OAI22_X1 port map( A1 => n6356, A2 => n4054, B1 => n4084, B2 => n4053
                           , ZN => n1746);
   U561 : OAI22_X1 port map( A1 => n6601, A2 => n4054, B1 => n4085, B2 => n4053
                           , ZN => n1745);
   U562 : OAI22_X1 port map( A1 => n6357, A2 => n4054, B1 => n4086, B2 => n4053
                           , ZN => n1744);
   U563 : OAI22_X1 port map( A1 => n6358, A2 => n4054, B1 => n4087, B2 => n4053
                           , ZN => n1743);
   U564 : OAI22_X1 port map( A1 => n6602, A2 => n4054, B1 => n4152, B2 => n4053
                           , ZN => n1742);
   U565 : OAI22_X1 port map( A1 => n6603, A2 => n4054, B1 => n4153, B2 => n4053
                           , ZN => n1741);
   U566 : OAI22_X1 port map( A1 => n6359, A2 => n4054, B1 => n4154, B2 => n4053
                           , ZN => n1740);
   U567 : OAI22_X1 port map( A1 => n6360, A2 => n4054, B1 => n4155, B2 => n4055
                           , ZN => n1739);
   U568 : OAI22_X1 port map( A1 => n6361, A2 => n4054, B1 => n4156, B2 => n4055
                           , ZN => n1738);
   U569 : OAI22_X1 port map( A1 => n6604, A2 => n4054, B1 => n4157, B2 => n4055
                           , ZN => n1737);
   U570 : OAI22_X1 port map( A1 => n6605, A2 => n4054, B1 => n4158, B2 => n4055
                           , ZN => n1736);
   U571 : OAI22_X1 port map( A1 => n6362, A2 => n4054, B1 => n4159, B2 => n4055
                           , ZN => n1735);
   U572 : OAI22_X1 port map( A1 => n6606, A2 => n4054, B1 => n4160, B2 => n4055
                           , ZN => n1734);
   U573 : OAI22_X1 port map( A1 => n6607, A2 => n4054, B1 => n4161, B2 => n4055
                           , ZN => n1733);
   U574 : OAI22_X1 port map( A1 => n6608, A2 => n4056, B1 => n4162, B2 => n4055
                           , ZN => n1732);
   U575 : OAI22_X1 port map( A1 => n6363, A2 => n4054, B1 => n4163, B2 => n4055
                           , ZN => n1731);
   U576 : OAI22_X1 port map( A1 => n6609, A2 => n4054, B1 => n4164, B2 => n4053
                           , ZN => n1730);
   U577 : OAI22_X1 port map( A1 => n6364, A2 => n4054, B1 => n4165, B2 => n4053
                           , ZN => n1729);
   U578 : OAI22_X1 port map( A1 => n6610, A2 => n4054, B1 => n4167, B2 => n4053
                           , ZN => n1728);
   U579 : OAI22_X1 port map( A1 => n6611, A2 => n4054, B1 => n4168, B2 => n4055
                           , ZN => n1727);
   U580 : OAI22_X1 port map( A1 => n6365, A2 => n4056, B1 => n4170, B2 => n4055
                           , ZN => n1726);
   U581 : OAI22_X1 port map( A1 => n6612, A2 => n4056, B1 => n4171, B2 => n4055
                           , ZN => n1725);
   U582 : OAI22_X1 port map( A1 => n6613, A2 => n4056, B1 => n4172, B2 => n4055
                           , ZN => n1724);
   U583 : OAI22_X1 port map( A1 => n6366, A2 => n4056, B1 => n4173, B2 => n4055
                           , ZN => n1723);
   U584 : OAI22_X1 port map( A1 => n6106, A2 => n4056, B1 => n4174, B2 => n4055
                           , ZN => n1722);
   U585 : OAI22_X1 port map( A1 => n6367, A2 => n4056, B1 => n4175, B2 => n4055
                           , ZN => n1721);
   U586 : OAI22_X1 port map( A1 => n6614, A2 => n4056, B1 => n4176, B2 => n4055
                           , ZN => n1720);
   U587 : OAI22_X1 port map( A1 => n6107, A2 => n4056, B1 => n4178, B2 => n4055
                           , ZN => n1719);
   U588 : NAND2_X1 port map( A1 => n4137, A2 => n4060, ZN => n4059);
   U589 : CLKBUF_X1 port map( A => n4059, Z => n4057);
   U590 : OAI22_X1 port map( A1 => n5849, A2 => n4058, B1 => n4107, B2 => n4057
                           , ZN => n1718);
   U591 : OAI22_X1 port map( A1 => n6615, A2 => n4058, B1 => n4145, B2 => n4057
                           , ZN => n1717);
   U592 : OAI22_X1 port map( A1 => n6616, A2 => n4058, B1 => n4146, B2 => n4057
                           , ZN => n1716);
   U593 : OAI22_X1 port map( A1 => n6368, A2 => n4058, B1 => n4147, B2 => n4057
                           , ZN => n1715);
   U594 : OAI22_X1 port map( A1 => n6108, A2 => n4058, B1 => n4148, B2 => n4057
                           , ZN => n1714);
   U595 : OAI22_X1 port map( A1 => n5850, A2 => n4058, B1 => n4149, B2 => n4057
                           , ZN => n1713);
   U596 : OAI22_X1 port map( A1 => n6617, A2 => n4058, B1 => n4150, B2 => n4057
                           , ZN => n1712);
   U597 : OAI22_X1 port map( A1 => n6369, A2 => n4058, B1 => n4151, B2 => n4057
                           , ZN => n1711);
   U598 : OAI22_X1 port map( A1 => n6109, A2 => n4058, B1 => n4152, B2 => n4057
                           , ZN => n1710);
   U599 : OAI22_X1 port map( A1 => n5851, A2 => n4058, B1 => n4153, B2 => n4057
                           , ZN => n1709);
   U600 : OAI22_X1 port map( A1 => n6110, A2 => n4058, B1 => n4154, B2 => n4057
                           , ZN => n1708);
   U601 : OAI22_X1 port map( A1 => n6370, A2 => n4058, B1 => n4155, B2 => n4059
                           , ZN => n1707);
   U602 : OAI22_X1 port map( A1 => n6618, A2 => n4058, B1 => n4156, B2 => n4059
                           , ZN => n1706);
   U603 : OAI22_X1 port map( A1 => n6619, A2 => n4058, B1 => n4157, B2 => n4059
                           , ZN => n1705);
   U604 : OAI22_X1 port map( A1 => n6371, A2 => n4058, B1 => n4158, B2 => n4059
                           , ZN => n1704);
   U605 : OAI22_X1 port map( A1 => n6111, A2 => n4058, B1 => n4159, B2 => n4059
                           , ZN => n1703);
   U606 : OAI22_X1 port map( A1 => n6372, A2 => n4058, B1 => n4160, B2 => n4059
                           , ZN => n1702);
   U607 : OAI22_X1 port map( A1 => n6620, A2 => n4058, B1 => n4161, B2 => n4059
                           , ZN => n1701);
   U608 : OAI22_X1 port map( A1 => n6112, A2 => n4058, B1 => n4162, B2 => n4059
                           , ZN => n1700);
   U609 : OAI22_X1 port map( A1 => n6621, A2 => n4058, B1 => n4163, B2 => n4059
                           , ZN => n1699);
   U610 : OAI22_X1 port map( A1 => n6113, A2 => n4058, B1 => n4164, B2 => n4057
                           , ZN => n1698);
   U611 : OAI22_X1 port map( A1 => n6622, A2 => n4058, B1 => n4165, B2 => n4057
                           , ZN => n1697);
   U612 : OAI22_X1 port map( A1 => n6373, A2 => n4058, B1 => n4167, B2 => n4057
                           , ZN => n1696);
   U613 : OAI22_X1 port map( A1 => n6623, A2 => n4058, B1 => n4168, B2 => n4059
                           , ZN => n1695);
   U614 : OAI22_X1 port map( A1 => n5852, A2 => n4058, B1 => n4170, B2 => n4059
                           , ZN => n1694);
   U615 : OAI22_X1 port map( A1 => n5853, A2 => n4058, B1 => n4171, B2 => n4059
                           , ZN => n1693);
   U616 : OAI22_X1 port map( A1 => n6374, A2 => n4058, B1 => n4172, B2 => n4059
                           , ZN => n1692);
   U617 : OAI22_X1 port map( A1 => n5854, A2 => n4058, B1 => n4173, B2 => n4059
                           , ZN => n1691);
   U618 : OAI22_X1 port map( A1 => n6375, A2 => n4058, B1 => n4174, B2 => n4059
                           , ZN => n1690);
   U619 : OAI22_X1 port map( A1 => n6624, A2 => n4058, B1 => n4175, B2 => n4059
                           , ZN => n1689);
   U620 : OAI22_X1 port map( A1 => n5855, A2 => n4058, B1 => n4176, B2 => n4059
                           , ZN => n1688);
   U621 : OAI22_X1 port map( A1 => n6376, A2 => n4058, B1 => n4178, B2 => n4059
                           , ZN => n1687);
   U622 : NAND2_X1 port map( A1 => n4143, A2 => n4060, ZN => n4063);
   U623 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4061, ZN => n4062);
   U624 : OAI22_X1 port map( A1 => n6114, A2 => n4062, B1 => n4107, B2 => n4061
                           , ZN => n1686);
   U625 : OAI22_X1 port map( A1 => n5856, A2 => n4062, B1 => n4145, B2 => n4061
                           , ZN => n1685);
   U626 : OAI22_X1 port map( A1 => n6115, A2 => n4062, B1 => n4146, B2 => n4061
                           , ZN => n1684);
   U627 : OAI22_X1 port map( A1 => n6116, A2 => n4062, B1 => n4147, B2 => n4061
                           , ZN => n1683);
   U628 : OAI22_X1 port map( A1 => n5857, A2 => n4062, B1 => n4148, B2 => n4061
                           , ZN => n1682);
   U629 : OAI22_X1 port map( A1 => n6117, A2 => n4062, B1 => n4149, B2 => n4061
                           , ZN => n1681);
   U630 : OAI22_X1 port map( A1 => n6118, A2 => n4062, B1 => n4150, B2 => n4061
                           , ZN => n1680);
   U631 : OAI22_X1 port map( A1 => n5858, A2 => n4062, B1 => n4151, B2 => n4061
                           , ZN => n1679);
   U632 : OAI22_X1 port map( A1 => n5859, A2 => n4062, B1 => n4152, B2 => n4061
                           , ZN => n1678);
   U633 : OAI22_X1 port map( A1 => n6119, A2 => n4062, B1 => n4153, B2 => n4061
                           , ZN => n1677);
   U634 : OAI22_X1 port map( A1 => n5860, A2 => n4062, B1 => n4154, B2 => n4061
                           , ZN => n1676);
   U635 : OAI22_X1 port map( A1 => n6120, A2 => n4062, B1 => n4155, B2 => n4063
                           , ZN => n1675);
   U636 : OAI22_X1 port map( A1 => n6121, A2 => n4062, B1 => n4156, B2 => n4063
                           , ZN => n1674);
   U637 : OAI22_X1 port map( A1 => n6122, A2 => n4062, B1 => n4157, B2 => n4063
                           , ZN => n1673);
   U638 : OAI22_X1 port map( A1 => n5861, A2 => n4062, B1 => n4158, B2 => n4063
                           , ZN => n1672);
   U639 : OAI22_X1 port map( A1 => n5862, A2 => n4062, B1 => n4159, B2 => n4063
                           , ZN => n1671);
   U640 : OAI22_X1 port map( A1 => n6123, A2 => n4062, B1 => n4160, B2 => n4063
                           , ZN => n1670);
   U641 : OAI22_X1 port map( A1 => n5863, A2 => n4062, B1 => n4161, B2 => n4063
                           , ZN => n1669);
   U642 : CLKBUF_X1 port map( A => n4062, Z => n4064);
   U643 : OAI22_X1 port map( A1 => n6124, A2 => n4064, B1 => n4162, B2 => n4063
                           , ZN => n1668);
   U644 : OAI22_X1 port map( A1 => n5864, A2 => n4062, B1 => n4163, B2 => n4063
                           , ZN => n1667);
   U645 : OAI22_X1 port map( A1 => n6125, A2 => n4062, B1 => n4164, B2 => n4061
                           , ZN => n1666);
   U646 : OAI22_X1 port map( A1 => n5865, A2 => n4062, B1 => n4165, B2 => n4061
                           , ZN => n1665);
   U647 : OAI22_X1 port map( A1 => n6126, A2 => n4062, B1 => n4167, B2 => n4061
                           , ZN => n1664);
   U648 : OAI22_X1 port map( A1 => n6127, A2 => n4062, B1 => n4168, B2 => n4063
                           , ZN => n1663);
   U649 : OAI22_X1 port map( A1 => n5866, A2 => n4064, B1 => n4170, B2 => n4063
                           , ZN => n1662);
   U650 : OAI22_X1 port map( A1 => n6128, A2 => n4064, B1 => n4171, B2 => n4063
                           , ZN => n1661);
   U651 : OAI22_X1 port map( A1 => n6129, A2 => n4064, B1 => n4172, B2 => n4063
                           , ZN => n1660);
   U652 : OAI22_X1 port map( A1 => n6130, A2 => n4064, B1 => n4173, B2 => n4063
                           , ZN => n1659);
   U653 : OAI22_X1 port map( A1 => n5867, A2 => n4064, B1 => n4174, B2 => n4063
                           , ZN => n1658);
   U654 : OAI22_X1 port map( A1 => n6131, A2 => n4064, B1 => n4175, B2 => n4063
                           , ZN => n1657);
   U655 : OAI22_X1 port map( A1 => n6132, A2 => n4064, B1 => n4176, B2 => n4063
                           , ZN => n1656);
   U656 : OAI22_X1 port map( A1 => n5868, A2 => n4064, B1 => n4178, B2 => n4063
                           , ZN => n1655);
   U657 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(4), ZN => 
                           n4104);
   U658 : NAND2_X1 port map( A1 => n4106, A2 => n4099, ZN => n4067);
   U659 : CLKBUF_X1 port map( A => n4067, Z => n4065);
   U660 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4065, ZN => n4066);
   U661 : OAI22_X1 port map( A1 => n6249, A2 => n4066, B1 => n4107, B2 => n4065
                           , ZN => n1654);
   U662 : OAI22_X1 port map( A1 => n6377, A2 => n4066, B1 => n4145, B2 => n4065
                           , ZN => n1653);
   U663 : OAI22_X1 port map( A1 => n6378, A2 => n4066, B1 => n4146, B2 => n4065
                           , ZN => n1652);
   U664 : OAI22_X1 port map( A1 => n6625, A2 => n4066, B1 => n4147, B2 => n4065
                           , ZN => n1651);
   U665 : OAI22_X1 port map( A1 => n6379, A2 => n4066, B1 => n4148, B2 => n4065
                           , ZN => n1650);
   U666 : OAI22_X1 port map( A1 => n6380, A2 => n4066, B1 => n4149, B2 => n4065
                           , ZN => n1649);
   U667 : OAI22_X1 port map( A1 => n6381, A2 => n4066, B1 => n4150, B2 => n4065
                           , ZN => n1648);
   U668 : OAI22_X1 port map( A1 => n6626, A2 => n4066, B1 => n4151, B2 => n4065
                           , ZN => n1647);
   U669 : OAI22_X1 port map( A1 => n5869, A2 => n4066, B1 => n4152, B2 => n4065
                           , ZN => n1646);
   U670 : OAI22_X1 port map( A1 => n6627, A2 => n4066, B1 => n4153, B2 => n4065
                           , ZN => n1645);
   U671 : OAI22_X1 port map( A1 => n6382, A2 => n4066, B1 => n4154, B2 => n4065
                           , ZN => n1644);
   U672 : OAI22_X1 port map( A1 => n6383, A2 => n4066, B1 => n4155, B2 => n4067
                           , ZN => n1643);
   U673 : OAI22_X1 port map( A1 => n5870, A2 => n4066, B1 => n4156, B2 => n4067
                           , ZN => n1642);
   U674 : OAI22_X1 port map( A1 => n6628, A2 => n4066, B1 => n4157, B2 => n4067
                           , ZN => n1641);
   U675 : OAI22_X1 port map( A1 => n6384, A2 => n4066, B1 => n4158, B2 => n4067
                           , ZN => n1640);
   U676 : OAI22_X1 port map( A1 => n6629, A2 => n4066, B1 => n4159, B2 => n4067
                           , ZN => n1639);
   U677 : OAI22_X1 port map( A1 => n6630, A2 => n4066, B1 => n4160, B2 => n4067
                           , ZN => n1638);
   U678 : CLKBUF_X1 port map( A => n4066, Z => n4068);
   U679 : OAI22_X1 port map( A1 => n6385, A2 => n4068, B1 => n4161, B2 => n4067
                           , ZN => n1637);
   U680 : OAI22_X1 port map( A1 => n6631, A2 => n4066, B1 => n4162, B2 => n4067
                           , ZN => n1636);
   U681 : OAI22_X1 port map( A1 => n6386, A2 => n4066, B1 => n4163, B2 => n4067
                           , ZN => n1635);
   U682 : OAI22_X1 port map( A1 => n6632, A2 => n4066, B1 => n4164, B2 => n4065
                           , ZN => n1634);
   U683 : OAI22_X1 port map( A1 => n5871, A2 => n4066, B1 => n4165, B2 => n4065
                           , ZN => n1633);
   U684 : OAI22_X1 port map( A1 => n6633, A2 => n4066, B1 => n4167, B2 => n4065
                           , ZN => n1632);
   U685 : OAI22_X1 port map( A1 => n6634, A2 => n4066, B1 => n4168, B2 => n4067
                           , ZN => n1631);
   U686 : OAI22_X1 port map( A1 => n6635, A2 => n4068, B1 => n4170, B2 => n4067
                           , ZN => n1630);
   U687 : OAI22_X1 port map( A1 => n6387, A2 => n4068, B1 => n4171, B2 => n4067
                           , ZN => n1629);
   U688 : OAI22_X1 port map( A1 => n6388, A2 => n4068, B1 => n4172, B2 => n4067
                           , ZN => n1628);
   U689 : OAI22_X1 port map( A1 => n6636, A2 => n4068, B1 => n4173, B2 => n4067
                           , ZN => n1627);
   U690 : OAI22_X1 port map( A1 => n6389, A2 => n4068, B1 => n4174, B2 => n4067
                           , ZN => n1626);
   U691 : OAI22_X1 port map( A1 => n6637, A2 => n4068, B1 => n4175, B2 => n4067
                           , ZN => n1625);
   U692 : OAI22_X1 port map( A1 => n5872, A2 => n4068, B1 => n4176, B2 => n4067
                           , ZN => n1624);
   U693 : OAI22_X1 port map( A1 => n6133, A2 => n4068, B1 => n4178, B2 => n4067
                           , ZN => n1623);
   U694 : NAND2_X1 port map( A1 => n4112, A2 => n4099, ZN => n4071);
   U695 : CLKBUF_X1 port map( A => n4071, Z => n4069);
   U696 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4069, ZN => n4070);
   U697 : OAI22_X1 port map( A1 => n6001, A2 => n4070, B1 => n4107, B2 => n4069
                           , ZN => n1622);
   U698 : OAI22_X1 port map( A1 => n6638, A2 => n4070, B1 => n4145, B2 => n4069
                           , ZN => n1621);
   U699 : OAI22_X1 port map( A1 => n6390, A2 => n4070, B1 => n4146, B2 => n4069
                           , ZN => n1620);
   U700 : OAI22_X1 port map( A1 => n6134, A2 => n4070, B1 => n4147, B2 => n4069
                           , ZN => n1619);
   U701 : OAI22_X1 port map( A1 => n5873, A2 => n4070, B1 => n4148, B2 => n4069
                           , ZN => n1618);
   U702 : OAI22_X1 port map( A1 => n6639, A2 => n4070, B1 => n4149, B2 => n4069
                           , ZN => n1617);
   U703 : OAI22_X1 port map( A1 => n6640, A2 => n4070, B1 => n4150, B2 => n4069
                           , ZN => n1616);
   U704 : OAI22_X1 port map( A1 => n6391, A2 => n4070, B1 => n4151, B2 => n4069
                           , ZN => n1615);
   U705 : OAI22_X1 port map( A1 => n6641, A2 => n4070, B1 => n4152, B2 => n4069
                           , ZN => n1614);
   U706 : OAI22_X1 port map( A1 => n5874, A2 => n4070, B1 => n4153, B2 => n4069
                           , ZN => n1613);
   U707 : OAI22_X1 port map( A1 => n5875, A2 => n4070, B1 => n4154, B2 => n4069
                           , ZN => n1612);
   U708 : OAI22_X1 port map( A1 => n5876, A2 => n4070, B1 => n4155, B2 => n4071
                           , ZN => n1611);
   U709 : OAI22_X1 port map( A1 => n6135, A2 => n4070, B1 => n4156, B2 => n4071
                           , ZN => n1610);
   U710 : OAI22_X1 port map( A1 => n6136, A2 => n4070, B1 => n4157, B2 => n4071
                           , ZN => n1609);
   U711 : OAI22_X1 port map( A1 => n6392, A2 => n4070, B1 => n4158, B2 => n4071
                           , ZN => n1608);
   U712 : OAI22_X1 port map( A1 => n6642, A2 => n4070, B1 => n4159, B2 => n4071
                           , ZN => n1607);
   U713 : OAI22_X1 port map( A1 => n6393, A2 => n4070, B1 => n4160, B2 => n4071
                           , ZN => n1606);
   U714 : CLKBUF_X1 port map( A => n4070, Z => n4072);
   U715 : OAI22_X1 port map( A1 => n6643, A2 => n4072, B1 => n4161, B2 => n4071
                           , ZN => n1605);
   U716 : OAI22_X1 port map( A1 => n5877, A2 => n4070, B1 => n4162, B2 => n4071
                           , ZN => n1604);
   U717 : OAI22_X1 port map( A1 => n6394, A2 => n4070, B1 => n4163, B2 => n4071
                           , ZN => n1603);
   U718 : OAI22_X1 port map( A1 => n6395, A2 => n4070, B1 => n4164, B2 => n4069
                           , ZN => n1602);
   U719 : OAI22_X1 port map( A1 => n6137, A2 => n4070, B1 => n4165, B2 => n4069
                           , ZN => n1601);
   U720 : OAI22_X1 port map( A1 => n6396, A2 => n4070, B1 => n4167, B2 => n4069
                           , ZN => n1600);
   U721 : OAI22_X1 port map( A1 => n5878, A2 => n4070, B1 => n4168, B2 => n4071
                           , ZN => n1599);
   U722 : OAI22_X1 port map( A1 => n6644, A2 => n4072, B1 => n4170, B2 => n4071
                           , ZN => n1598);
   U723 : OAI22_X1 port map( A1 => n6645, A2 => n4072, B1 => n4171, B2 => n4071
                           , ZN => n1597);
   U724 : OAI22_X1 port map( A1 => n6397, A2 => n4072, B1 => n4172, B2 => n4071
                           , ZN => n1596);
   U725 : OAI22_X1 port map( A1 => n6646, A2 => n4072, B1 => n4173, B2 => n4071
                           , ZN => n1595);
   U726 : OAI22_X1 port map( A1 => n5879, A2 => n4072, B1 => n4174, B2 => n4071
                           , ZN => n1594);
   U727 : OAI22_X1 port map( A1 => n6647, A2 => n4072, B1 => n4175, B2 => n4071
                           , ZN => n1593);
   U728 : OAI22_X1 port map( A1 => n5880, A2 => n4072, B1 => n4176, B2 => n4071
                           , ZN => n1592);
   U729 : OAI22_X1 port map( A1 => n5881, A2 => n4072, B1 => n4178, B2 => n4071
                           , ZN => n1591);
   U730 : NAND2_X1 port map( A1 => n4117, A2 => n4099, ZN => n4075);
   U731 : CLKBUF_X1 port map( A => n4075, Z => n4073);
   U732 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4073, ZN => n4074);
   U733 : OAI22_X1 port map( A1 => n6002, A2 => n4074, B1 => n4107, B2 => n4073
                           , ZN => n1590);
   U734 : OAI22_X1 port map( A1 => n6138, A2 => n4074, B1 => n4145, B2 => n4073
                           , ZN => n1589);
   U735 : OAI22_X1 port map( A1 => n6139, A2 => n4074, B1 => n4146, B2 => n4073
                           , ZN => n1588);
   U736 : OAI22_X1 port map( A1 => n6140, A2 => n4074, B1 => n4147, B2 => n4073
                           , ZN => n1587);
   U737 : OAI22_X1 port map( A1 => n6141, A2 => n4074, B1 => n4148, B2 => n4073
                           , ZN => n1586);
   U738 : OAI22_X1 port map( A1 => n5882, A2 => n4074, B1 => n4149, B2 => n4073
                           , ZN => n1585);
   U739 : OAI22_X1 port map( A1 => n6142, A2 => n4074, B1 => n4150, B2 => n4073
                           , ZN => n1584);
   U740 : OAI22_X1 port map( A1 => n6143, A2 => n4074, B1 => n4151, B2 => n4073
                           , ZN => n1583);
   U741 : OAI22_X1 port map( A1 => n6144, A2 => n4074, B1 => n4152, B2 => n4073
                           , ZN => n1582);
   U742 : OAI22_X1 port map( A1 => n5883, A2 => n4074, B1 => n4153, B2 => n4073
                           , ZN => n1581);
   U743 : OAI22_X1 port map( A1 => n5884, A2 => n4074, B1 => n4154, B2 => n4073
                           , ZN => n1580);
   U744 : OAI22_X1 port map( A1 => n6145, A2 => n4074, B1 => n4155, B2 => n4075
                           , ZN => n1579);
   U745 : OAI22_X1 port map( A1 => n5885, A2 => n4074, B1 => n4156, B2 => n4075
                           , ZN => n1578);
   U746 : OAI22_X1 port map( A1 => n5886, A2 => n4074, B1 => n4157, B2 => n4075
                           , ZN => n1577);
   U747 : OAI22_X1 port map( A1 => n6146, A2 => n4074, B1 => n4158, B2 => n4075
                           , ZN => n1576);
   U748 : OAI22_X1 port map( A1 => n6147, A2 => n4074, B1 => n4159, B2 => n4075
                           , ZN => n1575);
   U749 : OAI22_X1 port map( A1 => n6148, A2 => n4074, B1 => n4160, B2 => n4075
                           , ZN => n1574);
   U750 : CLKBUF_X1 port map( A => n4074, Z => n4076);
   U751 : OAI22_X1 port map( A1 => n6398, A2 => n4076, B1 => n4161, B2 => n4075
                           , ZN => n1573);
   U752 : OAI22_X1 port map( A1 => n6149, A2 => n4074, B1 => n4162, B2 => n4075
                           , ZN => n1572);
   U753 : OAI22_X1 port map( A1 => n5887, A2 => n4074, B1 => n4163, B2 => n4075
                           , ZN => n1571);
   U754 : OAI22_X1 port map( A1 => n6150, A2 => n4074, B1 => n4164, B2 => n4073
                           , ZN => n1570);
   U755 : OAI22_X1 port map( A1 => n5888, A2 => n4074, B1 => n4165, B2 => n4073
                           , ZN => n1569);
   U756 : OAI22_X1 port map( A1 => n6151, A2 => n4074, B1 => n4167, B2 => n4073
                           , ZN => n1568);
   U757 : OAI22_X1 port map( A1 => n5889, A2 => n4074, B1 => n4168, B2 => n4075
                           , ZN => n1567);
   U758 : OAI22_X1 port map( A1 => n5890, A2 => n4076, B1 => n4170, B2 => n4075
                           , ZN => n1566);
   U759 : OAI22_X1 port map( A1 => n6152, A2 => n4076, B1 => n4171, B2 => n4075
                           , ZN => n1565);
   U760 : OAI22_X1 port map( A1 => n6153, A2 => n4076, B1 => n4172, B2 => n4075
                           , ZN => n1564);
   U761 : OAI22_X1 port map( A1 => n5891, A2 => n4076, B1 => n4173, B2 => n4075
                           , ZN => n1563);
   U762 : OAI22_X1 port map( A1 => n6154, A2 => n4076, B1 => n4174, B2 => n4075
                           , ZN => n1562);
   U763 : OAI22_X1 port map( A1 => n5892, A2 => n4076, B1 => n4175, B2 => n4075
                           , ZN => n1561);
   U764 : OAI22_X1 port map( A1 => n6155, A2 => n4076, B1 => n4176, B2 => n4075
                           , ZN => n1560);
   U765 : OAI22_X1 port map( A1 => n6156, A2 => n4076, B1 => n4178, B2 => n4075
                           , ZN => n1559);
   U766 : NAND2_X1 port map( A1 => n4122, A2 => n4099, ZN => n4079);
   U767 : CLKBUF_X1 port map( A => n4079, Z => n4077);
   U768 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4077, ZN => n4078);
   U769 : OAI22_X1 port map( A1 => n6003, A2 => n4078, B1 => n4107, B2 => n4077
                           , ZN => n1558);
   U770 : OAI22_X1 port map( A1 => n5893, A2 => n4078, B1 => n4145, B2 => n4077
                           , ZN => n1557);
   U771 : OAI22_X1 port map( A1 => n6648, A2 => n4078, B1 => n4146, B2 => n4077
                           , ZN => n1556);
   U772 : OAI22_X1 port map( A1 => n5894, A2 => n4078, B1 => n4147, B2 => n4077
                           , ZN => n1555);
   U773 : OAI22_X1 port map( A1 => n5895, A2 => n4078, B1 => n4148, B2 => n4077
                           , ZN => n1554);
   U774 : OAI22_X1 port map( A1 => n6649, A2 => n4078, B1 => n4149, B2 => n4077
                           , ZN => n1553);
   U775 : OAI22_X1 port map( A1 => n6157, A2 => n4078, B1 => n4150, B2 => n4077
                           , ZN => n1552);
   U776 : OAI22_X1 port map( A1 => n5896, A2 => n4078, B1 => n4151, B2 => n4077
                           , ZN => n1551);
   U777 : OAI22_X1 port map( A1 => n6158, A2 => n4078, B1 => n4152, B2 => n4077
                           , ZN => n1550);
   U778 : OAI22_X1 port map( A1 => n6159, A2 => n4078, B1 => n4153, B2 => n4077
                           , ZN => n1549);
   U779 : OAI22_X1 port map( A1 => n6160, A2 => n4078, B1 => n4154, B2 => n4077
                           , ZN => n1548);
   U780 : OAI22_X1 port map( A1 => n6650, A2 => n4078, B1 => n4155, B2 => n4079
                           , ZN => n1547);
   U781 : OAI22_X1 port map( A1 => n6161, A2 => n4078, B1 => n4156, B2 => n4079
                           , ZN => n1546);
   U782 : OAI22_X1 port map( A1 => n6651, A2 => n4078, B1 => n4157, B2 => n4079
                           , ZN => n1545);
   U783 : OAI22_X1 port map( A1 => n6399, A2 => n4078, B1 => n4158, B2 => n4079
                           , ZN => n1544);
   U784 : OAI22_X1 port map( A1 => n6652, A2 => n4078, B1 => n4159, B2 => n4079
                           , ZN => n1543);
   U785 : OAI22_X1 port map( A1 => n6162, A2 => n4078, B1 => n4160, B2 => n4079
                           , ZN => n1542);
   U786 : CLKBUF_X1 port map( A => n4078, Z => n4080);
   U787 : OAI22_X1 port map( A1 => n6163, A2 => n4080, B1 => n4161, B2 => n4079
                           , ZN => n1541);
   U788 : OAI22_X1 port map( A1 => n5897, A2 => n4078, B1 => n4162, B2 => n4079
                           , ZN => n1540);
   U789 : OAI22_X1 port map( A1 => n6164, A2 => n4078, B1 => n4163, B2 => n4079
                           , ZN => n1539);
   U790 : OAI22_X1 port map( A1 => n6165, A2 => n4078, B1 => n4164, B2 => n4077
                           , ZN => n1538);
   U791 : OAI22_X1 port map( A1 => n6653, A2 => n4078, B1 => n4165, B2 => n4077
                           , ZN => n1537);
   U792 : OAI22_X1 port map( A1 => n5898, A2 => n4078, B1 => n4167, B2 => n4077
                           , ZN => n1536);
   U793 : OAI22_X1 port map( A1 => n5899, A2 => n4078, B1 => n4168, B2 => n4079
                           , ZN => n1535);
   U794 : OAI22_X1 port map( A1 => n5900, A2 => n4080, B1 => n4170, B2 => n4079
                           , ZN => n1534);
   U795 : OAI22_X1 port map( A1 => n5901, A2 => n4080, B1 => n4171, B2 => n4079
                           , ZN => n1533);
   U796 : OAI22_X1 port map( A1 => n6400, A2 => n4080, B1 => n4172, B2 => n4079
                           , ZN => n1532);
   U797 : OAI22_X1 port map( A1 => n5902, A2 => n4080, B1 => n4173, B2 => n4079
                           , ZN => n1531);
   U798 : OAI22_X1 port map( A1 => n6401, A2 => n4080, B1 => n4174, B2 => n4079
                           , ZN => n1530);
   U799 : OAI22_X1 port map( A1 => n5903, A2 => n4080, B1 => n4175, B2 => n4079
                           , ZN => n1529);
   U800 : OAI22_X1 port map( A1 => n6654, A2 => n4080, B1 => n4176, B2 => n4079
                           , ZN => n1528);
   U801 : OAI22_X1 port map( A1 => n6655, A2 => n4080, B1 => n4178, B2 => n4079
                           , ZN => n1527);
   U802 : NAND2_X1 port map( A1 => n4127, A2 => n4099, ZN => n4090);
   U803 : CLKBUF_X1 port map( A => n4090, Z => n4088);
   U804 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4088, ZN => n4089);
   U805 : OAI22_X1 port map( A1 => n6004, A2 => n4089, B1 => n4107, B2 => n4088
                           , ZN => n1526);
   U806 : OAI22_X1 port map( A1 => n5904, A2 => n4089, B1 => n4081, B2 => n4088
                           , ZN => n1525);
   U807 : OAI22_X1 port map( A1 => n5905, A2 => n4089, B1 => n4082, B2 => n4088
                           , ZN => n1524);
   U808 : OAI22_X1 port map( A1 => n6656, A2 => n4089, B1 => n4083, B2 => n4088
                           , ZN => n1523);
   U809 : OAI22_X1 port map( A1 => n6402, A2 => n4089, B1 => n4084, B2 => n4088
                           , ZN => n1522);
   U810 : OAI22_X1 port map( A1 => n5906, A2 => n4089, B1 => n4085, B2 => n4088
                           , ZN => n1521);
   U811 : OAI22_X1 port map( A1 => n5907, A2 => n4089, B1 => n4086, B2 => n4088
                           , ZN => n1520);
   U812 : OAI22_X1 port map( A1 => n6166, A2 => n4089, B1 => n4087, B2 => n4088
                           , ZN => n1519);
   U813 : OAI22_X1 port map( A1 => n6657, A2 => n4089, B1 => n4152, B2 => n4088
                           , ZN => n1518);
   U814 : OAI22_X1 port map( A1 => n6658, A2 => n4089, B1 => n4153, B2 => n4088
                           , ZN => n1517);
   U815 : OAI22_X1 port map( A1 => n5908, A2 => n4089, B1 => n4154, B2 => n4088
                           , ZN => n1516);
   U816 : OAI22_X1 port map( A1 => n6167, A2 => n4089, B1 => n4155, B2 => n4090
                           , ZN => n1515);
   U817 : OAI22_X1 port map( A1 => n5909, A2 => n4089, B1 => n4156, B2 => n4090
                           , ZN => n1514);
   U818 : OAI22_X1 port map( A1 => n6403, A2 => n4089, B1 => n4157, B2 => n4090
                           , ZN => n1513);
   U819 : OAI22_X1 port map( A1 => n6168, A2 => n4089, B1 => n4158, B2 => n4090
                           , ZN => n1512);
   U820 : OAI22_X1 port map( A1 => n5910, A2 => n4089, B1 => n4159, B2 => n4090
                           , ZN => n1511);
   U821 : OAI22_X1 port map( A1 => n6659, A2 => n4089, B1 => n4160, B2 => n4090
                           , ZN => n1510);
   U822 : CLKBUF_X1 port map( A => n4089, Z => n4091);
   U823 : OAI22_X1 port map( A1 => n6169, A2 => n4091, B1 => n4161, B2 => n4090
                           , ZN => n1509);
   U824 : OAI22_X1 port map( A1 => n5911, A2 => n4089, B1 => n4162, B2 => n4090
                           , ZN => n1508);
   U825 : OAI22_X1 port map( A1 => n5912, A2 => n4089, B1 => n4163, B2 => n4090
                           , ZN => n1507);
   U826 : OAI22_X1 port map( A1 => n5913, A2 => n4089, B1 => n4164, B2 => n4088
                           , ZN => n1506);
   U827 : OAI22_X1 port map( A1 => n6404, A2 => n4089, B1 => n4165, B2 => n4088
                           , ZN => n1505);
   U828 : OAI22_X1 port map( A1 => n6405, A2 => n4089, B1 => n4167, B2 => n4088
                           , ZN => n1504);
   U829 : OAI22_X1 port map( A1 => n6170, A2 => n4089, B1 => n4168, B2 => n4090
                           , ZN => n1503);
   U830 : OAI22_X1 port map( A1 => n6660, A2 => n4091, B1 => n4170, B2 => n4090
                           , ZN => n1502);
   U831 : OAI22_X1 port map( A1 => n5914, A2 => n4091, B1 => n4171, B2 => n4090
                           , ZN => n1501);
   U832 : OAI22_X1 port map( A1 => n6661, A2 => n4091, B1 => n4172, B2 => n4090
                           , ZN => n1500);
   U833 : OAI22_X1 port map( A1 => n5915, A2 => n4091, B1 => n4173, B2 => n4090
                           , ZN => n1499);
   U834 : OAI22_X1 port map( A1 => n6662, A2 => n4091, B1 => n4174, B2 => n4090
                           , ZN => n1498);
   U835 : OAI22_X1 port map( A1 => n5916, A2 => n4091, B1 => n4175, B2 => n4090
                           , ZN => n1497);
   U836 : OAI22_X1 port map( A1 => n5917, A2 => n4091, B1 => n4176, B2 => n4090
                           , ZN => n1496);
   U837 : OAI22_X1 port map( A1 => n6406, A2 => n4091, B1 => n4178, B2 => n4090
                           , ZN => n1495);
   U838 : NAND2_X1 port map( A1 => n4132, A2 => n4099, ZN => n4094);
   U839 : CLKBUF_X1 port map( A => n4094, Z => n4092);
   U840 : OAI22_X1 port map( A1 => n6250, A2 => n4093, B1 => n4107, B2 => n4092
                           , ZN => n1494);
   U841 : OAI22_X1 port map( A1 => n6407, A2 => n4093, B1 => n4145, B2 => n4092
                           , ZN => n1493);
   U842 : OAI22_X1 port map( A1 => n6408, A2 => n4093, B1 => n4146, B2 => n4092
                           , ZN => n1492);
   U843 : OAI22_X1 port map( A1 => n6409, A2 => n4093, B1 => n4147, B2 => n4092
                           , ZN => n1491);
   U844 : OAI22_X1 port map( A1 => n6663, A2 => n4093, B1 => n4148, B2 => n4092
                           , ZN => n1490);
   U845 : OAI22_X1 port map( A1 => n6410, A2 => n4093, B1 => n4149, B2 => n4092
                           , ZN => n1489);
   U846 : OAI22_X1 port map( A1 => n6664, A2 => n4093, B1 => n4150, B2 => n4092
                           , ZN => n1488);
   U847 : OAI22_X1 port map( A1 => n6665, A2 => n4093, B1 => n4151, B2 => n4092
                           , ZN => n1487);
   U848 : OAI22_X1 port map( A1 => n6666, A2 => n4093, B1 => n4152, B2 => n4092
                           , ZN => n1486);
   U849 : OAI22_X1 port map( A1 => n6171, A2 => n4093, B1 => n4153, B2 => n4092
                           , ZN => n1485);
   U850 : OAI22_X1 port map( A1 => n6667, A2 => n4093, B1 => n4154, B2 => n4092
                           , ZN => n1484);
   U851 : OAI22_X1 port map( A1 => n5918, A2 => n4093, B1 => n4155, B2 => n4094
                           , ZN => n1483);
   U852 : OAI22_X1 port map( A1 => n6668, A2 => n4093, B1 => n4156, B2 => n4094
                           , ZN => n1482);
   U853 : OAI22_X1 port map( A1 => n5919, A2 => n4093, B1 => n4157, B2 => n4094
                           , ZN => n1481);
   U854 : OAI22_X1 port map( A1 => n6669, A2 => n4093, B1 => n4158, B2 => n4094
                           , ZN => n1480);
   U855 : OAI22_X1 port map( A1 => n6411, A2 => n4093, B1 => n4159, B2 => n4094
                           , ZN => n1479);
   U856 : OAI22_X1 port map( A1 => n6172, A2 => n4093, B1 => n4160, B2 => n4094
                           , ZN => n1478);
   U857 : OAI22_X1 port map( A1 => n5920, A2 => n4093, B1 => n4161, B2 => n4094
                           , ZN => n1477);
   U858 : OAI22_X1 port map( A1 => n6670, A2 => n4093, B1 => n4162, B2 => n4094
                           , ZN => n1476);
   U859 : OAI22_X1 port map( A1 => n6173, A2 => n4093, B1 => n4163, B2 => n4094
                           , ZN => n1475);
   U860 : OAI22_X1 port map( A1 => n6671, A2 => n4093, B1 => n4164, B2 => n4092
                           , ZN => n1474);
   U861 : OAI22_X1 port map( A1 => n5921, A2 => n4093, B1 => n4165, B2 => n4092
                           , ZN => n1473);
   U862 : OAI22_X1 port map( A1 => n6672, A2 => n4093, B1 => n4167, B2 => n4092
                           , ZN => n1472);
   U863 : OAI22_X1 port map( A1 => n6673, A2 => n4093, B1 => n4168, B2 => n4094
                           , ZN => n1471);
   U864 : OAI22_X1 port map( A1 => n6174, A2 => n4093, B1 => n4170, B2 => n4094
                           , ZN => n1470);
   U865 : OAI22_X1 port map( A1 => n6412, A2 => n4093, B1 => n4171, B2 => n4094
                           , ZN => n1469);
   U866 : OAI22_X1 port map( A1 => n6674, A2 => n4093, B1 => n4172, B2 => n4094
                           , ZN => n1468);
   U867 : OAI22_X1 port map( A1 => n6675, A2 => n4093, B1 => n4173, B2 => n4094
                           , ZN => n1467);
   U868 : OAI22_X1 port map( A1 => n6413, A2 => n4093, B1 => n4174, B2 => n4094
                           , ZN => n1466);
   U869 : OAI22_X1 port map( A1 => n6175, A2 => n4093, B1 => n4175, B2 => n4094
                           , ZN => n1465);
   U870 : OAI22_X1 port map( A1 => n6676, A2 => n4093, B1 => n4176, B2 => n4094
                           , ZN => n1464);
   U871 : OAI22_X1 port map( A1 => n6414, A2 => n4093, B1 => n4178, B2 => n4094
                           , ZN => n1463);
   U872 : NAND2_X1 port map( A1 => n4137, A2 => n4099, ZN => n4097);
   U873 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4095, ZN => n4096);
   U874 : OAI22_X1 port map( A1 => n6251, A2 => n4096, B1 => n4107, B2 => n4095
                           , ZN => n1462);
   U875 : OAI22_X1 port map( A1 => n6415, A2 => n4096, B1 => n4145, B2 => n4095
                           , ZN => n1461);
   U876 : OAI22_X1 port map( A1 => n6677, A2 => n4096, B1 => n4146, B2 => n4095
                           , ZN => n1460);
   U877 : OAI22_X1 port map( A1 => n6416, A2 => n4096, B1 => n4147, B2 => n4095
                           , ZN => n1459);
   U878 : OAI22_X1 port map( A1 => n6678, A2 => n4096, B1 => n4148, B2 => n4095
                           , ZN => n1458);
   U879 : OAI22_X1 port map( A1 => n6417, A2 => n4096, B1 => n4149, B2 => n4095
                           , ZN => n1457);
   U880 : OAI22_X1 port map( A1 => n6418, A2 => n4096, B1 => n4150, B2 => n4095
                           , ZN => n1456);
   U881 : OAI22_X1 port map( A1 => n6679, A2 => n4096, B1 => n4151, B2 => n4095
                           , ZN => n1455);
   U882 : OAI22_X1 port map( A1 => n6176, A2 => n4096, B1 => n4152, B2 => n4095
                           , ZN => n1454);
   U883 : OAI22_X1 port map( A1 => n6419, A2 => n4096, B1 => n4153, B2 => n4095
                           , ZN => n1453);
   U884 : OAI22_X1 port map( A1 => n6177, A2 => n4096, B1 => n4154, B2 => n4095
                           , ZN => n1452);
   U885 : OAI22_X1 port map( A1 => n6680, A2 => n4096, B1 => n4155, B2 => n4097
                           , ZN => n1451);
   U886 : OAI22_X1 port map( A1 => n6681, A2 => n4096, B1 => n4156, B2 => n4097
                           , ZN => n1450);
   U887 : OAI22_X1 port map( A1 => n5922, A2 => n4096, B1 => n4157, B2 => n4097
                           , ZN => n1449);
   U888 : OAI22_X1 port map( A1 => n6682, A2 => n4096, B1 => n4158, B2 => n4097
                           , ZN => n1448);
   U889 : OAI22_X1 port map( A1 => n6178, A2 => n4096, B1 => n4159, B2 => n4097
                           , ZN => n1447);
   U890 : OAI22_X1 port map( A1 => n6420, A2 => n4096, B1 => n4160, B2 => n4097
                           , ZN => n1446);
   U891 : CLKBUF_X1 port map( A => n4096, Z => n4098);
   U892 : OAI22_X1 port map( A1 => n6683, A2 => n4098, B1 => n4161, B2 => n4097
                           , ZN => n1445);
   U893 : OAI22_X1 port map( A1 => n6421, A2 => n4096, B1 => n4162, B2 => n4097
                           , ZN => n1444);
   U894 : OAI22_X1 port map( A1 => n6179, A2 => n4096, B1 => n4163, B2 => n4097
                           , ZN => n1443);
   U895 : OAI22_X1 port map( A1 => n6684, A2 => n4096, B1 => n4164, B2 => n4095
                           , ZN => n1442);
   U896 : OAI22_X1 port map( A1 => n6422, A2 => n4096, B1 => n4165, B2 => n4095
                           , ZN => n1441);
   U897 : OAI22_X1 port map( A1 => n6685, A2 => n4096, B1 => n4167, B2 => n4095
                           , ZN => n1440);
   U898 : OAI22_X1 port map( A1 => n6423, A2 => n4096, B1 => n4168, B2 => n4097
                           , ZN => n1439);
   U899 : OAI22_X1 port map( A1 => n6686, A2 => n4098, B1 => n4170, B2 => n4097
                           , ZN => n1438);
   U900 : OAI22_X1 port map( A1 => n6687, A2 => n4098, B1 => n4171, B2 => n4097
                           , ZN => n1437);
   U901 : OAI22_X1 port map( A1 => n5923, A2 => n4098, B1 => n4172, B2 => n4097
                           , ZN => n1436);
   U902 : OAI22_X1 port map( A1 => n6688, A2 => n4098, B1 => n4173, B2 => n4097
                           , ZN => n1435);
   U903 : OAI22_X1 port map( A1 => n6180, A2 => n4098, B1 => n4174, B2 => n4097
                           , ZN => n1434);
   U904 : OAI22_X1 port map( A1 => n6424, A2 => n4098, B1 => n4175, B2 => n4097
                           , ZN => n1433);
   U905 : OAI22_X1 port map( A1 => n6425, A2 => n4098, B1 => n4176, B2 => n4097
                           , ZN => n1432);
   U906 : OAI22_X1 port map( A1 => n6426, A2 => n4098, B1 => n4178, B2 => n4097
                           , ZN => n1431);
   U907 : NAND2_X1 port map( A1 => n4143, A2 => n4099, ZN => n4102);
   U908 : CLKBUF_X1 port map( A => n4102, Z => n4100);
   U909 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4100, ZN => n4101);
   U910 : OAI22_X1 port map( A1 => n5733, A2 => n4101, B1 => n4107, B2 => n4100
                           , ZN => n1430);
   U911 : OAI22_X1 port map( A1 => n6181, A2 => n4101, B1 => n4145, B2 => n4100
                           , ZN => n1429);
   U912 : OAI22_X1 port map( A1 => n6182, A2 => n4101, B1 => n4146, B2 => n4100
                           , ZN => n1428);
   U913 : OAI22_X1 port map( A1 => n6183, A2 => n4101, B1 => n4147, B2 => n4100
                           , ZN => n1427);
   U914 : OAI22_X1 port map( A1 => n6184, A2 => n4101, B1 => n4148, B2 => n4100
                           , ZN => n1426);
   U915 : OAI22_X1 port map( A1 => n5924, A2 => n4101, B1 => n4149, B2 => n4100
                           , ZN => n1425);
   U916 : OAI22_X1 port map( A1 => n5925, A2 => n4101, B1 => n4150, B2 => n4100
                           , ZN => n1424);
   U917 : OAI22_X1 port map( A1 => n5926, A2 => n4101, B1 => n4151, B2 => n4100
                           , ZN => n1423);
   U918 : OAI22_X1 port map( A1 => n5927, A2 => n4101, B1 => n4152, B2 => n4100
                           , ZN => n1422);
   U919 : OAI22_X1 port map( A1 => n5928, A2 => n4101, B1 => n4153, B2 => n4100
                           , ZN => n1421);
   U920 : OAI22_X1 port map( A1 => n6185, A2 => n4101, B1 => n4154, B2 => n4100
                           , ZN => n1420);
   U921 : OAI22_X1 port map( A1 => n5929, A2 => n4101, B1 => n4155, B2 => n4102
                           , ZN => n1419);
   U922 : OAI22_X1 port map( A1 => n6186, A2 => n4101, B1 => n4156, B2 => n4102
                           , ZN => n1418);
   U923 : OAI22_X1 port map( A1 => n6187, A2 => n4101, B1 => n4157, B2 => n4102
                           , ZN => n1417);
   U924 : OAI22_X1 port map( A1 => n6188, A2 => n4101, B1 => n4158, B2 => n4102
                           , ZN => n1416);
   U925 : OAI22_X1 port map( A1 => n5930, A2 => n4101, B1 => n4159, B2 => n4102
                           , ZN => n1415);
   U926 : OAI22_X1 port map( A1 => n5931, A2 => n4101, B1 => n4160, B2 => n4102
                           , ZN => n1414);
   U927 : CLKBUF_X1 port map( A => n4101, Z => n4103);
   U928 : OAI22_X1 port map( A1 => n5932, A2 => n4103, B1 => n4161, B2 => n4102
                           , ZN => n1413);
   U929 : OAI22_X1 port map( A1 => n6689, A2 => n4101, B1 => n4162, B2 => n4102
                           , ZN => n1412);
   U930 : OAI22_X1 port map( A1 => n5933, A2 => n4101, B1 => n4163, B2 => n4102
                           , ZN => n1411);
   U931 : OAI22_X1 port map( A1 => n5934, A2 => n4101, B1 => n4164, B2 => n4100
                           , ZN => n1410);
   U932 : OAI22_X1 port map( A1 => n5935, A2 => n4101, B1 => n4165, B2 => n4100
                           , ZN => n1409);
   U933 : OAI22_X1 port map( A1 => n6189, A2 => n4101, B1 => n4167, B2 => n4100
                           , ZN => n1408);
   U934 : OAI22_X1 port map( A1 => n6190, A2 => n4101, B1 => n4168, B2 => n4102
                           , ZN => n1407);
   U935 : OAI22_X1 port map( A1 => n6191, A2 => n4103, B1 => n4170, B2 => n4102
                           , ZN => n1406);
   U936 : OAI22_X1 port map( A1 => n6427, A2 => n4103, B1 => n4171, B2 => n4102
                           , ZN => n1405);
   U937 : OAI22_X1 port map( A1 => n6192, A2 => n4103, B1 => n4172, B2 => n4102
                           , ZN => n1404);
   U938 : OAI22_X1 port map( A1 => n5936, A2 => n4103, B1 => n4173, B2 => n4102
                           , ZN => n1403);
   U939 : OAI22_X1 port map( A1 => n6193, A2 => n4103, B1 => n4174, B2 => n4102
                           , ZN => n1402);
   U940 : OAI22_X1 port map( A1 => n6690, A2 => n4103, B1 => n4175, B2 => n4102
                           , ZN => n1401);
   U941 : OAI22_X1 port map( A1 => n5937, A2 => n4103, B1 => n4176, B2 => n4102
                           , ZN => n1400);
   U942 : OAI22_X1 port map( A1 => n5938, A2 => n4103, B1 => n4178, B2 => n4102
                           , ZN => n1399);
   U943 : NOR2_X1 port map( A1 => n4105, A2 => n4104, ZN => n4142);
   U944 : NAND2_X1 port map( A1 => n4106, A2 => n4142, ZN => n4110);
   U945 : CLKBUF_X1 port map( A => n4110, Z => n4108);
   U946 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4108, ZN => n4109);
   U947 : CLKBUF_X1 port map( A => n4107, Z => n4144);
   U948 : OAI22_X1 port map( A1 => n6252, A2 => n4109, B1 => n4144, B2 => n4108
                           , ZN => n1398);
   U949 : OAI22_X1 port map( A1 => n6691, A2 => n4109, B1 => n4145, B2 => n4108
                           , ZN => n1397);
   U950 : OAI22_X1 port map( A1 => n6428, A2 => n4109, B1 => n4146, B2 => n4108
                           , ZN => n1396);
   U951 : OAI22_X1 port map( A1 => n6692, A2 => n4109, B1 => n4147, B2 => n4108
                           , ZN => n1395);
   U952 : OAI22_X1 port map( A1 => n6693, A2 => n4109, B1 => n4148, B2 => n4108
                           , ZN => n1394);
   U953 : OAI22_X1 port map( A1 => n6694, A2 => n4109, B1 => n4149, B2 => n4108
                           , ZN => n1393);
   U954 : OAI22_X1 port map( A1 => n6429, A2 => n4109, B1 => n4150, B2 => n4108
                           , ZN => n1392);
   U955 : OAI22_X1 port map( A1 => n6430, A2 => n4109, B1 => n4151, B2 => n4108
                           , ZN => n1391);
   U956 : OAI22_X1 port map( A1 => n6431, A2 => n4109, B1 => n4152, B2 => n4108
                           , ZN => n1390);
   U957 : OAI22_X1 port map( A1 => n6695, A2 => n4109, B1 => n4153, B2 => n4108
                           , ZN => n1389);
   U958 : OAI22_X1 port map( A1 => n6696, A2 => n4109, B1 => n4154, B2 => n4108
                           , ZN => n1388);
   U959 : OAI22_X1 port map( A1 => n6432, A2 => n4109, B1 => n4155, B2 => n4110
                           , ZN => n1387);
   U960 : OAI22_X1 port map( A1 => n6433, A2 => n4109, B1 => n4156, B2 => n4110
                           , ZN => n1386);
   U961 : OAI22_X1 port map( A1 => n6434, A2 => n4109, B1 => n4157, B2 => n4110
                           , ZN => n1385);
   U962 : OAI22_X1 port map( A1 => n6435, A2 => n4109, B1 => n4158, B2 => n4110
                           , ZN => n1384);
   U963 : OAI22_X1 port map( A1 => n6436, A2 => n4109, B1 => n4159, B2 => n4110
                           , ZN => n1383);
   U964 : OAI22_X1 port map( A1 => n6437, A2 => n4109, B1 => n4160, B2 => n4110
                           , ZN => n1382);
   U965 : CLKBUF_X1 port map( A => n4109, Z => n4111);
   U966 : OAI22_X1 port map( A1 => n6438, A2 => n4111, B1 => n4161, B2 => n4110
                           , ZN => n1381);
   U967 : OAI22_X1 port map( A1 => n6697, A2 => n4109, B1 => n4162, B2 => n4110
                           , ZN => n1380);
   U968 : OAI22_X1 port map( A1 => n6698, A2 => n4109, B1 => n4163, B2 => n4110
                           , ZN => n1379);
   U969 : OAI22_X1 port map( A1 => n6439, A2 => n4109, B1 => n4164, B2 => n4108
                           , ZN => n1378);
   U970 : OAI22_X1 port map( A1 => n6699, A2 => n4109, B1 => n4165, B2 => n4108
                           , ZN => n1377);
   U971 : OAI22_X1 port map( A1 => n6440, A2 => n4109, B1 => n4167, B2 => n4108
                           , ZN => n1376);
   U972 : OAI22_X1 port map( A1 => n6700, A2 => n4109, B1 => n4168, B2 => n4110
                           , ZN => n1375);
   U973 : OAI22_X1 port map( A1 => n6441, A2 => n4111, B1 => n4170, B2 => n4110
                           , ZN => n1374);
   U974 : OAI22_X1 port map( A1 => n6701, A2 => n4111, B1 => n4171, B2 => n4110
                           , ZN => n1373);
   U975 : OAI22_X1 port map( A1 => n6442, A2 => n4111, B1 => n4172, B2 => n4110
                           , ZN => n1372);
   U976 : OAI22_X1 port map( A1 => n6443, A2 => n4111, B1 => n4173, B2 => n4110
                           , ZN => n1371);
   U977 : OAI22_X1 port map( A1 => n6702, A2 => n4111, B1 => n4174, B2 => n4110
                           , ZN => n1370);
   U978 : OAI22_X1 port map( A1 => n6444, A2 => n4111, B1 => n4175, B2 => n4110
                           , ZN => n1369);
   U979 : OAI22_X1 port map( A1 => n6445, A2 => n4111, B1 => n4176, B2 => n4110
                           , ZN => n1368);
   U980 : OAI22_X1 port map( A1 => n6446, A2 => n4111, B1 => n4178, B2 => n4110
                           , ZN => n1367);
   U981 : NAND2_X1 port map( A1 => n4112, A2 => n4142, ZN => n4115);
   U982 : CLKBUF_X1 port map( A => n4115, Z => n4113);
   U983 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4113, ZN => n4114);
   U984 : OAI22_X1 port map( A1 => n6005, A2 => n4114, B1 => n4144, B2 => n4113
                           , ZN => n1366);
   U985 : OAI22_X1 port map( A1 => n6194, A2 => n4114, B1 => n4145, B2 => n4113
                           , ZN => n1365);
   U986 : OAI22_X1 port map( A1 => n5939, A2 => n4114, B1 => n4146, B2 => n4113
                           , ZN => n1364);
   U987 : OAI22_X1 port map( A1 => n5940, A2 => n4114, B1 => n4147, B2 => n4113
                           , ZN => n1363);
   U988 : OAI22_X1 port map( A1 => n6195, A2 => n4114, B1 => n4148, B2 => n4113
                           , ZN => n1362);
   U989 : OAI22_X1 port map( A1 => n5941, A2 => n4114, B1 => n4149, B2 => n4113
                           , ZN => n1361);
   U990 : OAI22_X1 port map( A1 => n5942, A2 => n4114, B1 => n4150, B2 => n4113
                           , ZN => n1360);
   U991 : OAI22_X1 port map( A1 => n5943, A2 => n4114, B1 => n4151, B2 => n4113
                           , ZN => n1359);
   U992 : OAI22_X1 port map( A1 => n5944, A2 => n4114, B1 => n4152, B2 => n4113
                           , ZN => n1358);
   U993 : OAI22_X1 port map( A1 => n6196, A2 => n4114, B1 => n4153, B2 => n4113
                           , ZN => n1357);
   U994 : OAI22_X1 port map( A1 => n6447, A2 => n4114, B1 => n4154, B2 => n4113
                           , ZN => n1356);
   U995 : OAI22_X1 port map( A1 => n5945, A2 => n4114, B1 => n4155, B2 => n4115
                           , ZN => n1355);
   U996 : OAI22_X1 port map( A1 => n6448, A2 => n4114, B1 => n4156, B2 => n4115
                           , ZN => n1354);
   U997 : OAI22_X1 port map( A1 => n6449, A2 => n4114, B1 => n4157, B2 => n4115
                           , ZN => n1353);
   U998 : OAI22_X1 port map( A1 => n5946, A2 => n4114, B1 => n4158, B2 => n4115
                           , ZN => n1352);
   U999 : OAI22_X1 port map( A1 => n5947, A2 => n4114, B1 => n4159, B2 => n4115
                           , ZN => n1351);
   U1000 : OAI22_X1 port map( A1 => n5948, A2 => n4114, B1 => n4160, B2 => 
                           n4115, ZN => n1350);
   U1001 : CLKBUF_X1 port map( A => n4114, Z => n4116);
   U1002 : OAI22_X1 port map( A1 => n5949, A2 => n4116, B1 => n4161, B2 => 
                           n4115, ZN => n1349);
   U1003 : OAI22_X1 port map( A1 => n6197, A2 => n4114, B1 => n4162, B2 => 
                           n4115, ZN => n1348);
   U1004 : OAI22_X1 port map( A1 => n6198, A2 => n4114, B1 => n4163, B2 => 
                           n4115, ZN => n1347);
   U1005 : OAI22_X1 port map( A1 => n6199, A2 => n4114, B1 => n4164, B2 => 
                           n4113, ZN => n1346);
   U1006 : OAI22_X1 port map( A1 => n5950, A2 => n4114, B1 => n4165, B2 => 
                           n4113, ZN => n1345);
   U1007 : OAI22_X1 port map( A1 => n5951, A2 => n4114, B1 => n4167, B2 => 
                           n4113, ZN => n1344);
   U1008 : OAI22_X1 port map( A1 => n6450, A2 => n4114, B1 => n4168, B2 => 
                           n4115, ZN => n1343);
   U1009 : OAI22_X1 port map( A1 => n5952, A2 => n4116, B1 => n4170, B2 => 
                           n4115, ZN => n1342);
   U1010 : OAI22_X1 port map( A1 => n6200, A2 => n4116, B1 => n4171, B2 => 
                           n4115, ZN => n1341);
   U1011 : OAI22_X1 port map( A1 => n6201, A2 => n4116, B1 => n4172, B2 => 
                           n4115, ZN => n1340);
   U1012 : OAI22_X1 port map( A1 => n5953, A2 => n4116, B1 => n4173, B2 => 
                           n4115, ZN => n1339);
   U1013 : OAI22_X1 port map( A1 => n5954, A2 => n4116, B1 => n4174, B2 => 
                           n4115, ZN => n1338);
   U1014 : OAI22_X1 port map( A1 => n6202, A2 => n4116, B1 => n4175, B2 => 
                           n4115, ZN => n1337);
   U1015 : OAI22_X1 port map( A1 => n6703, A2 => n4116, B1 => n4176, B2 => 
                           n4115, ZN => n1336);
   U1016 : OAI22_X1 port map( A1 => n5955, A2 => n4116, B1 => n4178, B2 => 
                           n4115, ZN => n1335);
   U1017 : NAND2_X1 port map( A1 => n4117, A2 => n4142, ZN => n4120);
   U1018 : CLKBUF_X1 port map( A => n4120, Z => n4118);
   U1019 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4118, ZN => n4119);
   U1020 : OAI22_X1 port map( A1 => n6006, A2 => n4119, B1 => n4144, B2 => 
                           n4118, ZN => n1334);
   U1021 : OAI22_X1 port map( A1 => n6704, A2 => n4119, B1 => n4145, B2 => 
                           n4118, ZN => n1333);
   U1022 : OAI22_X1 port map( A1 => n5956, A2 => n4119, B1 => n4146, B2 => 
                           n4118, ZN => n1332);
   U1023 : OAI22_X1 port map( A1 => n5957, A2 => n4119, B1 => n4147, B2 => 
                           n4118, ZN => n1331);
   U1024 : OAI22_X1 port map( A1 => n5958, A2 => n4119, B1 => n4148, B2 => 
                           n4118, ZN => n1330);
   U1025 : OAI22_X1 port map( A1 => n6451, A2 => n4119, B1 => n4149, B2 => 
                           n4118, ZN => n1329);
   U1026 : OAI22_X1 port map( A1 => n6203, A2 => n4119, B1 => n4150, B2 => 
                           n4118, ZN => n1328);
   U1027 : OAI22_X1 port map( A1 => n5959, A2 => n4119, B1 => n4151, B2 => 
                           n4118, ZN => n1327);
   U1028 : OAI22_X1 port map( A1 => n6452, A2 => n4119, B1 => n4152, B2 => 
                           n4118, ZN => n1326);
   U1029 : OAI22_X1 port map( A1 => n6453, A2 => n4119, B1 => n4153, B2 => 
                           n4118, ZN => n1325);
   U1030 : OAI22_X1 port map( A1 => n6454, A2 => n4119, B1 => n4154, B2 => 
                           n4118, ZN => n1324);
   U1031 : OAI22_X1 port map( A1 => n5960, A2 => n4119, B1 => n4155, B2 => 
                           n4120, ZN => n1323);
   U1032 : OAI22_X1 port map( A1 => n6204, A2 => n4119, B1 => n4156, B2 => 
                           n4120, ZN => n1322);
   U1033 : OAI22_X1 port map( A1 => n6705, A2 => n4119, B1 => n4157, B2 => 
                           n4120, ZN => n1321);
   U1034 : OAI22_X1 port map( A1 => n6205, A2 => n4119, B1 => n4158, B2 => 
                           n4120, ZN => n1320);
   U1035 : OAI22_X1 port map( A1 => n6206, A2 => n4119, B1 => n4159, B2 => 
                           n4120, ZN => n1319);
   U1036 : OAI22_X1 port map( A1 => n6207, A2 => n4119, B1 => n4160, B2 => 
                           n4120, ZN => n1318);
   U1037 : CLKBUF_X1 port map( A => n4119, Z => n4121);
   U1038 : OAI22_X1 port map( A1 => n5961, A2 => n4121, B1 => n4161, B2 => 
                           n4120, ZN => n1317);
   U1039 : OAI22_X1 port map( A1 => n5962, A2 => n4119, B1 => n4162, B2 => 
                           n4120, ZN => n1316);
   U1040 : OAI22_X1 port map( A1 => n6455, A2 => n4119, B1 => n4163, B2 => 
                           n4120, ZN => n1315);
   U1041 : OAI22_X1 port map( A1 => n6706, A2 => n4119, B1 => n4164, B2 => 
                           n4118, ZN => n1314);
   U1042 : OAI22_X1 port map( A1 => n6208, A2 => n4119, B1 => n4165, B2 => 
                           n4118, ZN => n1313);
   U1043 : OAI22_X1 port map( A1 => n6707, A2 => n4119, B1 => n4167, B2 => 
                           n4118, ZN => n1312);
   U1044 : OAI22_X1 port map( A1 => n6209, A2 => n4119, B1 => n4168, B2 => 
                           n4120, ZN => n1311);
   U1045 : OAI22_X1 port map( A1 => n6708, A2 => n4121, B1 => n4170, B2 => 
                           n4120, ZN => n1310);
   U1046 : OAI22_X1 port map( A1 => n6709, A2 => n4121, B1 => n4171, B2 => 
                           n4120, ZN => n1309);
   U1047 : OAI22_X1 port map( A1 => n5963, A2 => n4121, B1 => n4172, B2 => 
                           n4120, ZN => n1308);
   U1048 : OAI22_X1 port map( A1 => n6710, A2 => n4121, B1 => n4173, B2 => 
                           n4120, ZN => n1307);
   U1049 : OAI22_X1 port map( A1 => n6210, A2 => n4121, B1 => n4174, B2 => 
                           n4120, ZN => n1306);
   U1050 : OAI22_X1 port map( A1 => n6711, A2 => n4121, B1 => n4175, B2 => 
                           n4120, ZN => n1305);
   U1051 : OAI22_X1 port map( A1 => n6211, A2 => n4121, B1 => n4176, B2 => 
                           n4120, ZN => n1304);
   U1052 : OAI22_X1 port map( A1 => n6712, A2 => n4121, B1 => n4178, B2 => 
                           n4120, ZN => n1303);
   U1053 : NAND2_X1 port map( A1 => n4122, A2 => n4142, ZN => n4125);
   U1054 : CLKBUF_X1 port map( A => n4125, Z => n4123);
   U1055 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4123, ZN => n4124);
   U1056 : OAI22_X1 port map( A1 => n5734, A2 => n4124, B1 => n4144, B2 => 
                           n4123, ZN => n1302);
   U1057 : OAI22_X1 port map( A1 => n6212, A2 => n4124, B1 => n4145, B2 => 
                           n4123, ZN => n1301);
   U1058 : OAI22_X1 port map( A1 => n6213, A2 => n4124, B1 => n4146, B2 => 
                           n4123, ZN => n1300);
   U1059 : OAI22_X1 port map( A1 => n6214, A2 => n4124, B1 => n4147, B2 => 
                           n4123, ZN => n1299);
   U1060 : OAI22_X1 port map( A1 => n6215, A2 => n4124, B1 => n4148, B2 => 
                           n4123, ZN => n1298);
   U1061 : OAI22_X1 port map( A1 => n6216, A2 => n4124, B1 => n4149, B2 => 
                           n4123, ZN => n1297);
   U1062 : OAI22_X1 port map( A1 => n5964, A2 => n4124, B1 => n4150, B2 => 
                           n4123, ZN => n1296);
   U1063 : OAI22_X1 port map( A1 => n6217, A2 => n4124, B1 => n4151, B2 => 
                           n4123, ZN => n1295);
   U1064 : OAI22_X1 port map( A1 => n5965, A2 => n4124, B1 => n4152, B2 => 
                           n4123, ZN => n1294);
   U1065 : OAI22_X1 port map( A1 => n5966, A2 => n4124, B1 => n4153, B2 => 
                           n4123, ZN => n1293);
   U1066 : OAI22_X1 port map( A1 => n6218, A2 => n4124, B1 => n4154, B2 => 
                           n4123, ZN => n1292);
   U1067 : OAI22_X1 port map( A1 => n6219, A2 => n4124, B1 => n4155, B2 => 
                           n4125, ZN => n1291);
   U1068 : OAI22_X1 port map( A1 => n5967, A2 => n4124, B1 => n4156, B2 => 
                           n4125, ZN => n1290);
   U1069 : OAI22_X1 port map( A1 => n6220, A2 => n4124, B1 => n4157, B2 => 
                           n4125, ZN => n1289);
   U1070 : OAI22_X1 port map( A1 => n5968, A2 => n4124, B1 => n4158, B2 => 
                           n4125, ZN => n1288);
   U1071 : OAI22_X1 port map( A1 => n5969, A2 => n4124, B1 => n4159, B2 => 
                           n4125, ZN => n1287);
   U1072 : OAI22_X1 port map( A1 => n6221, A2 => n4124, B1 => n4160, B2 => 
                           n4125, ZN => n1286);
   U1073 : CLKBUF_X1 port map( A => n4124, Z => n4126);
   U1074 : OAI22_X1 port map( A1 => n5970, A2 => n4126, B1 => n4161, B2 => 
                           n4125, ZN => n1285);
   U1075 : OAI22_X1 port map( A1 => n5971, A2 => n4124, B1 => n4162, B2 => 
                           n4125, ZN => n1284);
   U1076 : OAI22_X1 port map( A1 => n5972, A2 => n4124, B1 => n4163, B2 => 
                           n4125, ZN => n1283);
   U1077 : OAI22_X1 port map( A1 => n5973, A2 => n4124, B1 => n4164, B2 => 
                           n4123, ZN => n1282);
   U1078 : OAI22_X1 port map( A1 => n6222, A2 => n4124, B1 => n4165, B2 => 
                           n4123, ZN => n1281);
   U1079 : OAI22_X1 port map( A1 => n5974, A2 => n4124, B1 => n4167, B2 => 
                           n4123, ZN => n1280);
   U1080 : OAI22_X1 port map( A1 => n6223, A2 => n4124, B1 => n4168, B2 => 
                           n4125, ZN => n1279);
   U1081 : OAI22_X1 port map( A1 => n5975, A2 => n4126, B1 => n4170, B2 => 
                           n4125, ZN => n1278);
   U1082 : OAI22_X1 port map( A1 => n5976, A2 => n4126, B1 => n4171, B2 => 
                           n4125, ZN => n1277);
   U1083 : OAI22_X1 port map( A1 => n6224, A2 => n4126, B1 => n4172, B2 => 
                           n4125, ZN => n1276);
   U1084 : OAI22_X1 port map( A1 => n5977, A2 => n4126, B1 => n4173, B2 => 
                           n4125, ZN => n1275);
   U1085 : OAI22_X1 port map( A1 => n5978, A2 => n4126, B1 => n4174, B2 => 
                           n4125, ZN => n1274);
   U1086 : OAI22_X1 port map( A1 => n6225, A2 => n4126, B1 => n4175, B2 => 
                           n4125, ZN => n1273);
   U1087 : OAI22_X1 port map( A1 => n5979, A2 => n4126, B1 => n4176, B2 => 
                           n4125, ZN => n1272);
   U1088 : OAI22_X1 port map( A1 => n6226, A2 => n4126, B1 => n4178, B2 => 
                           n4125, ZN => n1271);
   U1089 : NAND2_X1 port map( A1 => n4127, A2 => n4142, ZN => n4130);
   U1090 : CLKBUF_X1 port map( A => n4130, Z => n4128);
   U1091 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4128, ZN => n4129);
   U1092 : OAI22_X1 port map( A1 => n6007, A2 => n4129, B1 => n4144, B2 => 
                           n4128, ZN => n1270);
   U1093 : OAI22_X1 port map( A1 => n6456, A2 => n4129, B1 => n4145, B2 => 
                           n4128, ZN => n1269);
   U1094 : OAI22_X1 port map( A1 => n6713, A2 => n4129, B1 => n4146, B2 => 
                           n4128, ZN => n1268);
   U1095 : OAI22_X1 port map( A1 => n6457, A2 => n4129, B1 => n4147, B2 => 
                           n4128, ZN => n1267);
   U1096 : OAI22_X1 port map( A1 => n6458, A2 => n4129, B1 => n4148, B2 => 
                           n4128, ZN => n1266);
   U1097 : OAI22_X1 port map( A1 => n6714, A2 => n4129, B1 => n4149, B2 => 
                           n4128, ZN => n1265);
   U1098 : OAI22_X1 port map( A1 => n6715, A2 => n4129, B1 => n4150, B2 => 
                           n4128, ZN => n1264);
   U1099 : OAI22_X1 port map( A1 => n6459, A2 => n4129, B1 => n4151, B2 => 
                           n4128, ZN => n1263);
   U1100 : OAI22_X1 port map( A1 => n6716, A2 => n4129, B1 => n4152, B2 => 
                           n4128, ZN => n1262);
   U1101 : OAI22_X1 port map( A1 => n6460, A2 => n4129, B1 => n4153, B2 => 
                           n4128, ZN => n1261);
   U1102 : OAI22_X1 port map( A1 => n6717, A2 => n4129, B1 => n4154, B2 => 
                           n4128, ZN => n1260);
   U1103 : OAI22_X1 port map( A1 => n6718, A2 => n4129, B1 => n4155, B2 => 
                           n4130, ZN => n1259);
   U1104 : OAI22_X1 port map( A1 => n6719, A2 => n4129, B1 => n4156, B2 => 
                           n4130, ZN => n1258);
   U1105 : OAI22_X1 port map( A1 => n6720, A2 => n4129, B1 => n4157, B2 => 
                           n4130, ZN => n1257);
   U1106 : OAI22_X1 port map( A1 => n5980, A2 => n4129, B1 => n4158, B2 => 
                           n4130, ZN => n1256);
   U1107 : OAI22_X1 port map( A1 => n6721, A2 => n4129, B1 => n4159, B2 => 
                           n4130, ZN => n1255);
   U1108 : OAI22_X1 port map( A1 => n6461, A2 => n4129, B1 => n4160, B2 => 
                           n4130, ZN => n1254);
   U1109 : CLKBUF_X1 port map( A => n4129, Z => n4131);
   U1110 : OAI22_X1 port map( A1 => n6722, A2 => n4131, B1 => n4161, B2 => 
                           n4130, ZN => n1253);
   U1111 : OAI22_X1 port map( A1 => n6462, A2 => n4129, B1 => n4162, B2 => 
                           n4130, ZN => n1252);
   U1112 : OAI22_X1 port map( A1 => n6723, A2 => n4129, B1 => n4163, B2 => 
                           n4130, ZN => n1251);
   U1113 : OAI22_X1 port map( A1 => n6463, A2 => n4129, B1 => n4164, B2 => 
                           n4128, ZN => n1250);
   U1114 : OAI22_X1 port map( A1 => n6724, A2 => n4129, B1 => n4165, B2 => 
                           n4128, ZN => n1249);
   U1115 : OAI22_X1 port map( A1 => n6227, A2 => n4129, B1 => n4167, B2 => 
                           n4128, ZN => n1248);
   U1116 : OAI22_X1 port map( A1 => n6725, A2 => n4129, B1 => n4168, B2 => 
                           n4130, ZN => n1247);
   U1117 : OAI22_X1 port map( A1 => n6726, A2 => n4131, B1 => n4170, B2 => 
                           n4130, ZN => n1246);
   U1118 : OAI22_X1 port map( A1 => n5981, A2 => n4131, B1 => n4171, B2 => 
                           n4130, ZN => n1245);
   U1119 : OAI22_X1 port map( A1 => n6464, A2 => n4131, B1 => n4172, B2 => 
                           n4130, ZN => n1244);
   U1120 : OAI22_X1 port map( A1 => n6727, A2 => n4131, B1 => n4173, B2 => 
                           n4130, ZN => n1243);
   U1121 : OAI22_X1 port map( A1 => n6728, A2 => n4131, B1 => n4174, B2 => 
                           n4130, ZN => n1242);
   U1122 : OAI22_X1 port map( A1 => n6465, A2 => n4131, B1 => n4175, B2 => 
                           n4130, ZN => n1241);
   U1123 : OAI22_X1 port map( A1 => n6729, A2 => n4131, B1 => n4176, B2 => 
                           n4130, ZN => n1240);
   U1124 : OAI22_X1 port map( A1 => n6730, A2 => n4131, B1 => n4178, B2 => 
                           n4130, ZN => n1239);
   U1125 : NAND2_X1 port map( A1 => n4132, A2 => n4142, ZN => n4135);
   U1126 : CLKBUF_X1 port map( A => n4135, Z => n4133);
   U1127 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4133, ZN => n4134);
   U1128 : OAI22_X1 port map( A1 => n6008, A2 => n4134, B1 => n4144, B2 => 
                           n4133, ZN => n1238);
   U1129 : OAI22_X1 port map( A1 => n6731, A2 => n4134, B1 => n4145, B2 => 
                           n4133, ZN => n1237);
   U1130 : OAI22_X1 port map( A1 => n6228, A2 => n4134, B1 => n4146, B2 => 
                           n4133, ZN => n1236);
   U1131 : OAI22_X1 port map( A1 => n6466, A2 => n4134, B1 => n4147, B2 => 
                           n4133, ZN => n1235);
   U1132 : OAI22_X1 port map( A1 => n6467, A2 => n4134, B1 => n4148, B2 => 
                           n4133, ZN => n1234);
   U1133 : OAI22_X1 port map( A1 => n6229, A2 => n4134, B1 => n4149, B2 => 
                           n4133, ZN => n1233);
   U1134 : OAI22_X1 port map( A1 => n6468, A2 => n4134, B1 => n4150, B2 => 
                           n4133, ZN => n1232);
   U1135 : OAI22_X1 port map( A1 => n6732, A2 => n4134, B1 => n4151, B2 => 
                           n4133, ZN => n1231);
   U1136 : OAI22_X1 port map( A1 => n6733, A2 => n4134, B1 => n4152, B2 => 
                           n4133, ZN => n1230);
   U1137 : OAI22_X1 port map( A1 => n6734, A2 => n4134, B1 => n4153, B2 => 
                           n4133, ZN => n1229);
   U1138 : OAI22_X1 port map( A1 => n6735, A2 => n4134, B1 => n4154, B2 => 
                           n4133, ZN => n1228);
   U1139 : OAI22_X1 port map( A1 => n6736, A2 => n4134, B1 => n4155, B2 => 
                           n4135, ZN => n1227);
   U1140 : OAI22_X1 port map( A1 => n6469, A2 => n4134, B1 => n4156, B2 => 
                           n4135, ZN => n1226);
   U1141 : OAI22_X1 port map( A1 => n6470, A2 => n4134, B1 => n4157, B2 => 
                           n4135, ZN => n1225);
   U1142 : OAI22_X1 port map( A1 => n6737, A2 => n4134, B1 => n4158, B2 => 
                           n4135, ZN => n1224);
   U1143 : OAI22_X1 port map( A1 => n6738, A2 => n4134, B1 => n4159, B2 => 
                           n4135, ZN => n1223);
   U1144 : OAI22_X1 port map( A1 => n6471, A2 => n4134, B1 => n4160, B2 => 
                           n4135, ZN => n1222);
   U1145 : CLKBUF_X1 port map( A => n4134, Z => n4136);
   U1146 : OAI22_X1 port map( A1 => n6739, A2 => n4136, B1 => n4161, B2 => 
                           n4135, ZN => n1221);
   U1147 : OAI22_X1 port map( A1 => n6472, A2 => n4134, B1 => n4162, B2 => 
                           n4135, ZN => n1220);
   U1148 : OAI22_X1 port map( A1 => n6740, A2 => n4134, B1 => n4163, B2 => 
                           n4135, ZN => n1219);
   U1149 : OAI22_X1 port map( A1 => n6473, A2 => n4134, B1 => n4164, B2 => 
                           n4133, ZN => n1218);
   U1150 : OAI22_X1 port map( A1 => n6741, A2 => n4134, B1 => n4165, B2 => 
                           n4133, ZN => n1217);
   U1151 : OAI22_X1 port map( A1 => n6474, A2 => n4134, B1 => n4167, B2 => 
                           n4133, ZN => n1216);
   U1152 : OAI22_X1 port map( A1 => n6475, A2 => n4134, B1 => n4168, B2 => 
                           n4135, ZN => n1215);
   U1153 : OAI22_X1 port map( A1 => n6476, A2 => n4136, B1 => n4170, B2 => 
                           n4135, ZN => n1214);
   U1154 : OAI22_X1 port map( A1 => n6230, A2 => n4136, B1 => n4171, B2 => 
                           n4135, ZN => n1213);
   U1155 : OAI22_X1 port map( A1 => n6477, A2 => n4136, B1 => n4172, B2 => 
                           n4135, ZN => n1212);
   U1156 : OAI22_X1 port map( A1 => n6478, A2 => n4136, B1 => n4173, B2 => 
                           n4135, ZN => n1211);
   U1157 : OAI22_X1 port map( A1 => n6742, A2 => n4136, B1 => n4174, B2 => 
                           n4135, ZN => n1210);
   U1158 : OAI22_X1 port map( A1 => n6479, A2 => n4136, B1 => n4175, B2 => 
                           n4135, ZN => n1209);
   U1159 : OAI22_X1 port map( A1 => n6743, A2 => n4136, B1 => n4176, B2 => 
                           n4135, ZN => n1208);
   U1160 : OAI22_X1 port map( A1 => n6480, A2 => n4136, B1 => n4178, B2 => 
                           n4135, ZN => n1207);
   U1161 : NAND2_X1 port map( A1 => n4137, A2 => n4142, ZN => n4140);
   U1162 : CLKBUF_X1 port map( A => n4140, Z => n4138);
   U1163 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4138, ZN => n4139);
   U1164 : OAI22_X1 port map( A1 => n5735, A2 => n4139, B1 => n4144, B2 => 
                           n4138, ZN => n1206);
   U1165 : OAI22_X1 port map( A1 => n5982, A2 => n4139, B1 => n4145, B2 => 
                           n4138, ZN => n1205);
   U1166 : OAI22_X1 port map( A1 => n5983, A2 => n4139, B1 => n4146, B2 => 
                           n4138, ZN => n1204);
   U1167 : OAI22_X1 port map( A1 => n6744, A2 => n4139, B1 => n4147, B2 => 
                           n4138, ZN => n1203);
   U1168 : OAI22_X1 port map( A1 => n5984, A2 => n4139, B1 => n4148, B2 => 
                           n4138, ZN => n1202);
   U1169 : OAI22_X1 port map( A1 => n6231, A2 => n4139, B1 => n4149, B2 => 
                           n4138, ZN => n1201);
   U1170 : OAI22_X1 port map( A1 => n6745, A2 => n4139, B1 => n4150, B2 => 
                           n4138, ZN => n1200);
   U1171 : OAI22_X1 port map( A1 => n6232, A2 => n4139, B1 => n4151, B2 => 
                           n4138, ZN => n1199);
   U1172 : OAI22_X1 port map( A1 => n6481, A2 => n4139, B1 => n4152, B2 => 
                           n4138, ZN => n1198);
   U1173 : OAI22_X1 port map( A1 => n5985, A2 => n4139, B1 => n4153, B2 => 
                           n4138, ZN => n1197);
   U1174 : OAI22_X1 port map( A1 => n5986, A2 => n4139, B1 => n4154, B2 => 
                           n4138, ZN => n1196);
   U1175 : OAI22_X1 port map( A1 => n6482, A2 => n4139, B1 => n4155, B2 => 
                           n4140, ZN => n1195);
   U1176 : OAI22_X1 port map( A1 => n6746, A2 => n4139, B1 => n4156, B2 => 
                           n4140, ZN => n1194);
   U1177 : OAI22_X1 port map( A1 => n6233, A2 => n4139, B1 => n4157, B2 => 
                           n4140, ZN => n1193);
   U1178 : OAI22_X1 port map( A1 => n5987, A2 => n4139, B1 => n4158, B2 => 
                           n4140, ZN => n1192);
   U1179 : OAI22_X1 port map( A1 => n6483, A2 => n4139, B1 => n4159, B2 => 
                           n4140, ZN => n1191);
   U1180 : OAI22_X1 port map( A1 => n5988, A2 => n4139, B1 => n4160, B2 => 
                           n4140, ZN => n1190);
   U1181 : CLKBUF_X1 port map( A => n4139, Z => n4141);
   U1182 : OAI22_X1 port map( A1 => n6747, A2 => n4141, B1 => n4161, B2 => 
                           n4140, ZN => n1189);
   U1183 : OAI22_X1 port map( A1 => n6748, A2 => n4139, B1 => n4162, B2 => 
                           n4140, ZN => n1188);
   U1184 : OAI22_X1 port map( A1 => n6484, A2 => n4139, B1 => n4163, B2 => 
                           n4140, ZN => n1187);
   U1185 : OAI22_X1 port map( A1 => n6234, A2 => n4139, B1 => n4164, B2 => 
                           n4138, ZN => n1186);
   U1186 : OAI22_X1 port map( A1 => n6485, A2 => n4139, B1 => n4165, B2 => 
                           n4138, ZN => n1185);
   U1187 : OAI22_X1 port map( A1 => n5989, A2 => n4139, B1 => n4167, B2 => 
                           n4138, ZN => n1184);
   U1188 : OAI22_X1 port map( A1 => n5990, A2 => n4139, B1 => n4168, B2 => 
                           n4140, ZN => n1183);
   U1189 : OAI22_X1 port map( A1 => n5991, A2 => n4141, B1 => n4170, B2 => 
                           n4140, ZN => n1182);
   U1190 : OAI22_X1 port map( A1 => n6486, A2 => n4141, B1 => n4171, B2 => 
                           n4140, ZN => n1181);
   U1191 : OAI22_X1 port map( A1 => n6235, A2 => n4141, B1 => n4172, B2 => 
                           n4140, ZN => n1180);
   U1192 : OAI22_X1 port map( A1 => n6236, A2 => n4141, B1 => n4173, B2 => 
                           n4140, ZN => n1179);
   U1193 : OAI22_X1 port map( A1 => n5992, A2 => n4141, B1 => n4174, B2 => 
                           n4140, ZN => n1178);
   U1194 : OAI22_X1 port map( A1 => n5993, A2 => n4141, B1 => n4175, B2 => 
                           n4140, ZN => n1177);
   U1195 : OAI22_X1 port map( A1 => n6237, A2 => n4141, B1 => n4176, B2 => 
                           n4140, ZN => n1176);
   U1196 : OAI22_X1 port map( A1 => n6238, A2 => n4141, B1 => n4178, B2 => 
                           n4140, ZN => n1175);
   U1197 : NAND2_X1 port map( A1 => n4143, A2 => n4142, ZN => n4177);
   U1198 : CLKBUF_X1 port map( A => n4177, Z => n4166);
   U1199 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n4166, ZN => n4169);
   U1200 : OAI22_X1 port map( A1 => n5736, A2 => n4169, B1 => n4144, B2 => 
                           n4166, ZN => n1174);
   U1201 : OAI22_X1 port map( A1 => n5994, A2 => n4169, B1 => n4145, B2 => 
                           n4166, ZN => n1173);
   U1202 : OAI22_X1 port map( A1 => n6749, A2 => n4169, B1 => n4146, B2 => 
                           n4166, ZN => n1172);
   U1203 : OAI22_X1 port map( A1 => n5995, A2 => n4169, B1 => n4147, B2 => 
                           n4166, ZN => n1171);
   U1204 : OAI22_X1 port map( A1 => n6750, A2 => n4169, B1 => n4148, B2 => 
                           n4166, ZN => n1170);
   U1205 : OAI22_X1 port map( A1 => n6239, A2 => n4169, B1 => n4149, B2 => 
                           n4166, ZN => n1169);
   U1206 : OAI22_X1 port map( A1 => n6240, A2 => n4169, B1 => n4150, B2 => 
                           n4166, ZN => n1168);
   U1207 : OAI22_X1 port map( A1 => n6487, A2 => n4169, B1 => n4151, B2 => 
                           n4166, ZN => n1167);
   U1208 : OAI22_X1 port map( A1 => n5996, A2 => n4169, B1 => n4152, B2 => 
                           n4166, ZN => n1166);
   U1209 : OAI22_X1 port map( A1 => n6751, A2 => n4169, B1 => n4153, B2 => 
                           n4166, ZN => n1165);
   U1210 : OAI22_X1 port map( A1 => n6488, A2 => n4169, B1 => n4154, B2 => 
                           n4166, ZN => n1164);
   U1211 : OAI22_X1 port map( A1 => n6752, A2 => n4169, B1 => n4155, B2 => 
                           n4177, ZN => n1163);
   U1212 : OAI22_X1 port map( A1 => n6489, A2 => n4169, B1 => n4156, B2 => 
                           n4177, ZN => n1162);
   U1213 : OAI22_X1 port map( A1 => n5997, A2 => n4169, B1 => n4157, B2 => 
                           n4177, ZN => n1161);
   U1214 : OAI22_X1 port map( A1 => n6753, A2 => n4169, B1 => n4158, B2 => 
                           n4177, ZN => n1160);
   U1215 : OAI22_X1 port map( A1 => n5998, A2 => n4169, B1 => n4159, B2 => 
                           n4177, ZN => n1159);
   U1216 : OAI22_X1 port map( A1 => n6754, A2 => n4169, B1 => n4160, B2 => 
                           n4177, ZN => n1158);
   U1217 : CLKBUF_X1 port map( A => n4169, Z => n4179);
   U1218 : OAI22_X1 port map( A1 => n6241, A2 => n4179, B1 => n4161, B2 => 
                           n4177, ZN => n1157);
   U1219 : OAI22_X1 port map( A1 => n6242, A2 => n4169, B1 => n4162, B2 => 
                           n4177, ZN => n1156);
   U1220 : OAI22_X1 port map( A1 => n6755, A2 => n4169, B1 => n4163, B2 => 
                           n4177, ZN => n1155);
   U1221 : OAI22_X1 port map( A1 => n5999, A2 => n4169, B1 => n4164, B2 => 
                           n4166, ZN => n1154);
   U1222 : OAI22_X1 port map( A1 => n6756, A2 => n4169, B1 => n4165, B2 => 
                           n4166, ZN => n1153);
   U1223 : OAI22_X1 port map( A1 => n6243, A2 => n4169, B1 => n4167, B2 => 
                           n4166, ZN => n1152);
   U1224 : OAI22_X1 port map( A1 => n6490, A2 => n4169, B1 => n4168, B2 => 
                           n4177, ZN => n1151);
   U1225 : OAI22_X1 port map( A1 => n6000, A2 => n4179, B1 => n4170, B2 => 
                           n4177, ZN => n1150);
   U1226 : OAI22_X1 port map( A1 => n6244, A2 => n4179, B1 => n4171, B2 => 
                           n4177, ZN => n1149);
   U1227 : OAI22_X1 port map( A1 => n6245, A2 => n4179, B1 => n4172, B2 => 
                           n4177, ZN => n1148);
   U1228 : OAI22_X1 port map( A1 => n6246, A2 => n4179, B1 => n4173, B2 => 
                           n4177, ZN => n1147);
   U1229 : OAI22_X1 port map( A1 => n6491, A2 => n4179, B1 => n4174, B2 => 
                           n4177, ZN => n1146);
   U1230 : OAI22_X1 port map( A1 => n6247, A2 => n4179, B1 => n4175, B2 => 
                           n4177, ZN => n1145);
   U1231 : OAI22_X1 port map( A1 => n6492, A2 => n4179, B1 => n4176, B2 => 
                           n4177, ZN => n1144);
   U1232 : OAI22_X1 port map( A1 => n6248, A2 => n4179, B1 => n4178, B2 => 
                           n4177, ZN => n1143);
   U1233 : INV_X1 port map( A => ADD_RD2(3), ZN => n4202);
   U1234 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n4202, ZN => n4189);
   U1235 : INV_X1 port map( A => ADD_RD2(2), ZN => n4186);
   U1236 : OR3_X1 port map( A1 => n4186, A2 => ADD_RD2(0), A3 => ADD_RD2(1), ZN
                           => n4268);
   U1237 : NOR2_X1 port map( A1 => n4189, A2 => n4268, ZN => n4906);
   U1238 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n4188);
   U1239 : INV_X1 port map( A => ADD_RD2(1), ZN => n4184);
   U1240 : OR3_X1 port map( A1 => n4186, A2 => n4184, A3 => ADD_RD2(0), ZN => 
                           n4291);
   U1241 : NOR2_X1 port map( A1 => n4188, A2 => n4291, ZN => n4754);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n4906, B1 => 
                           REGISTERS_30_31_port, B2 => n4754, ZN => n4183);
   U1243 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), ZN => n4185);
   U1244 : NAND2_X1 port map( A1 => n4185, A2 => ADD_RD2(1), ZN => n4196);
   U1245 : NOR2_X1 port map( A1 => n4188, A2 => n4196, ZN => n4803);
   U1246 : INV_X1 port map( A => ADD_RD2(0), ZN => n4187);
   U1247 : OR3_X1 port map( A1 => n4186, A2 => n4187, A3 => n4184, ZN => n4245)
                           ;
   U1248 : NOR2_X1 port map( A1 => n4188, A2 => n4245, ZN => n4710);
   U1249 : CLKBUF_X1 port map( A => n4710, Z => n4921);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n4803, B1 => 
                           REGISTERS_31_31_port, B2 => n4921, ZN => n4182);
   U1251 : NOR2_X1 port map( A1 => n4189, A2 => n4196, ZN => n4882);
   U1252 : OR3_X1 port map( A1 => n4187, A2 => n4184, A3 => ADD_RD2(2), ZN => 
                           n4314);
   U1253 : NOR2_X1 port map( A1 => n4188, A2 => n4314, ZN => n4621);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_18_31_port, A2 => n4882, B1 => 
                           REGISTERS_27_31_port, B2 => n4621, ZN => n4181);
   U1255 : OR3_X1 port map( A1 => n4187, A2 => ADD_RD2(2), A3 => ADD_RD2(1), ZN
                           => n4225);
   U1256 : NOR2_X1 port map( A1 => n4188, A2 => n4225, ZN => n4825);
   U1257 : NOR2_X1 port map( A1 => n4189, A2 => n4245, ZN => n4905);
   U1258 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n4825, B1 => 
                           REGISTERS_23_31_port, B2 => n4905, ZN => n4180);
   U1259 : NAND4_X1 port map( A1 => n4183, A2 => n4182, A3 => n4181, A4 => 
                           n4180, ZN => n4195);
   U1260 : NAND2_X1 port map( A1 => n4185, A2 => n4184, ZN => n4197);
   U1261 : NOR2_X1 port map( A1 => n4197, A2 => n4189, ZN => n4856);
   U1262 : NOR2_X1 port map( A1 => n4188, A2 => n4268, ZN => n4881);
   U1263 : CLKBUF_X1 port map( A => n4881, Z => n4922);
   U1264 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n4856, B1 => 
                           REGISTERS_28_31_port, B2 => n4922, ZN => n4193);
   U1265 : NOR2_X1 port map( A1 => n4188, A2 => n4197, ZN => n4442);
   U1266 : OR3_X1 port map( A1 => n4187, A2 => n4186, A3 => ADD_RD2(1), ZN => 
                           n4244);
   U1267 : NOR2_X1 port map( A1 => n4188, A2 => n4244, ZN => n4855);
   U1268 : CLKBUF_X1 port map( A => n4855, Z => n4908);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n4442, B1 => 
                           REGISTERS_29_31_port, B2 => n4908, ZN => n4192);
   U1270 : NOR2_X1 port map( A1 => n4244, A2 => n4189, ZN => n4883);
   U1271 : CLKBUF_X1 port map( A => n4883, Z => n4916);
   U1272 : NOR2_X1 port map( A1 => n4189, A2 => n4314, ZN => n4920);
   U1273 : CLKBUF_X1 port map( A => n4920, Z => n4850);
   U1274 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n4916, B1 => 
                           REGISTERS_19_31_port, B2 => n4850, ZN => n4191);
   U1275 : NOR2_X1 port map( A1 => n4189, A2 => n4291, ZN => n4876);
   U1276 : CLKBUF_X1 port map( A => n4876, Z => n4910);
   U1277 : NOR2_X1 port map( A1 => n4189, A2 => n4225, ZN => n4804);
   U1278 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n4910, B1 => 
                           REGISTERS_17_31_port, B2 => n4804, ZN => n4190);
   U1279 : NAND4_X1 port map( A1 => n4193, A2 => n4192, A3 => n4191, A4 => 
                           n4190, ZN => n4194);
   U1280 : NOR2_X1 port map( A1 => n4195, A2 => n4194, ZN => n4210);
   U1281 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n4958, 
                           ZN => n4503);
   U1282 : CLKBUF_X1 port map( A => n4503, Z => n4728);
   U1283 : INV_X1 port map( A => n4314, ZN => n4741);
   U1284 : AOI22_X1 port map( A1 => n4741, A2 => REGISTERS_3_31_port, B1 => 
                           n4933, B2 => REGISTERS_2_31_port, ZN => n4201);
   U1285 : INV_X1 port map( A => n4291, ZN => n4929);
   U1286 : INV_X1 port map( A => n4245, ZN => n4944);
   U1287 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_6_31_port, B1 => 
                           n4944, B2 => REGISTERS_7_31_port, ZN => n4200);
   U1288 : INV_X1 port map( A => n4268, ZN => n4943);
   U1289 : INV_X1 port map( A => n4225, ZN => n4931);
   U1290 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_31_port, B1 => 
                           n4931, B2 => REGISTERS_1_31_port, ZN => n4199);
   U1291 : INV_X1 port map( A => n4244, ZN => n4721);
   U1292 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_31_port, B1 => 
                           n4721, B2 => REGISTERS_5_31_port, ZN => n4198);
   U1293 : NAND4_X1 port map( A1 => n4201, A2 => n4200, A3 => n4199, A4 => 
                           n4198, ZN => n4208);
   U1294 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n4202, A3 => n4958, ZN => 
                           n4434);
   U1295 : CLKBUF_X1 port map( A => n4434, Z => n4953);
   U1296 : INV_X1 port map( A => n4245, ZN => n4932);
   U1297 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_31_port, B1 => 
                           n4932, B2 => REGISTERS_15_31_port, ZN => n4206);
   U1298 : INV_X1 port map( A => n4268, ZN => n4816);
   U1299 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_31_port, B1 => 
                           n4929, B2 => REGISTERS_14_31_port, ZN => n4205);
   U1300 : INV_X1 port map( A => n4244, ZN => n4940);
   U1301 : INV_X1 port map( A => n4225, ZN => n4815);
   U1302 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_31_port, B1 => 
                           n4815, B2 => REGISTERS_9_31_port, ZN => n4204);
   U1303 : AOI22_X1 port map( A1 => n4741, A2 => REGISTERS_11_31_port, B1 => 
                           n4933, B2 => REGISTERS_10_31_port, ZN => n4203);
   U1304 : NAND4_X1 port map( A1 => n4206, A2 => n4205, A3 => n4204, A4 => 
                           n4203, ZN => n4207);
   U1305 : AOI22_X1 port map( A1 => n4728, A2 => n4208, B1 => n4953, B2 => 
                           n4207, ZN => n4209);
   U1306 : OAI21_X1 port map( B1 => n4958, B2 => n4210, A => n4209, ZN => N448)
                           ;
   U1307 : CLKBUF_X1 port map( A => n4906, Z => n4849);
   U1308 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_30_port, B1 => 
                           n4849, B2 => REGISTERS_20_30_port, ZN => n4214);
   U1309 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_30_port, B1 => 
                           n4921, B2 => REGISTERS_31_30_port, ZN => n4213);
   U1310 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_30_port, B1 => 
                           n4850, B2 => REGISTERS_19_30_port, ZN => n4212);
   U1311 : CLKBUF_X1 port map( A => n4754, Z => n4919);
   U1312 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_30_port, B1 => 
                           n4919, B2 => REGISTERS_30_30_port, ZN => n4211);
   U1313 : NAND4_X1 port map( A1 => n4214, A2 => n4213, A3 => n4212, A4 => 
                           n4211, ZN => n4220);
   U1314 : CLKBUF_X1 port map( A => n4803, Z => n4918);
   U1315 : CLKBUF_X1 port map( A => n4621, Z => n4915);
   U1316 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_30_port, B1 => 
                           n4915, B2 => REGISTERS_27_30_port, ZN => n4218);
   U1317 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_30_port, B1 => 
                           n4825, B2 => REGISTERS_25_30_port, ZN => n4217);
   U1318 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_30_port, B1 => 
                           n4905, B2 => REGISTERS_23_30_port, ZN => n4216);
   U1319 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_30_port, B1 => 
                           n4882, B2 => REGISTERS_18_30_port, ZN => n4215);
   U1320 : NAND4_X1 port map( A1 => n4218, A2 => n4217, A3 => n4216, A4 => 
                           n4215, ZN => n4219);
   U1321 : NOR2_X1 port map( A1 => n4220, A2 => n4219, ZN => n4233);
   U1322 : INV_X1 port map( A => n4291, ZN => n4947);
   U1323 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_5_30_port, B1 => 
                           n4947, B2 => REGISTERS_6_30_port, ZN => n4224);
   U1324 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_30_port, B1 => 
                           n4932, B2 => REGISTERS_7_30_port, ZN => n4223);
   U1325 : INV_X1 port map( A => n4314, ZN => n4934);
   U1326 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_1_30_port, B1 => 
                           n4934, B2 => REGISTERS_3_30_port, ZN => n4222);
   U1327 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_30_port, B1 => 
                           n4943, B2 => REGISTERS_4_30_port, ZN => n4221);
   U1328 : NAND4_X1 port map( A1 => n4224, A2 => n4223, A3 => n4222, A4 => 
                           n4221, ZN => n4231);
   U1329 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_30_port, B1 => 
                           n4933, B2 => REGISTERS_10_30_port, ZN => n4229);
   U1330 : INV_X1 port map( A => n4225, ZN => n4942);
   U1331 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_30_port, B1 => 
                           n4741, B2 => REGISTERS_11_30_port, ZN => n4228);
   U1332 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_30_port, B1 => 
                           n4816, B2 => REGISTERS_12_30_port, ZN => n4227);
   U1333 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_30_port, B1 => 
                           n4944, B2 => REGISTERS_15_30_port, ZN => n4226);
   U1334 : NAND4_X1 port map( A1 => n4229, A2 => n4228, A3 => n4227, A4 => 
                           n4226, ZN => n4230);
   U1335 : AOI22_X1 port map( A1 => n4728, A2 => n4231, B1 => n4953, B2 => 
                           n4230, ZN => n4232);
   U1336 : OAI21_X1 port map( B1 => n4958, B2 => n4233, A => n4232, ZN => N447)
                           ;
   U1337 : CLKBUF_X1 port map( A => n4882, Z => n4917);
   U1338 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_29_port, B1 => 
                           n4917, B2 => REGISTERS_18_29_port, ZN => n4237);
   U1339 : CLKBUF_X1 port map( A => n4856, Z => n4903);
   U1340 : CLKBUF_X1 port map( A => n4825, Z => n4907);
   U1341 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_29_port, B1 => 
                           n4907, B2 => REGISTERS_25_29_port, ZN => n4236);
   U1342 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_29_port, B1 => 
                           n4919, B2 => REGISTERS_30_29_port, ZN => n4235);
   U1343 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_29_port, B1 => 
                           n4849, B2 => REGISTERS_20_29_port, ZN => n4234);
   U1344 : NAND4_X1 port map( A1 => n4237, A2 => n4236, A3 => n4235, A4 => 
                           n4234, ZN => n4243);
   U1345 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_29_port, B1 => 
                           n4908, B2 => REGISTERS_29_29_port, ZN => n4241);
   U1346 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_29_port, B1 => 
                           n4621, B2 => REGISTERS_27_29_port, ZN => n4240);
   U1347 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_29_port, B1 => 
                           n4918, B2 => REGISTERS_26_29_port, ZN => n4239);
   U1348 : CLKBUF_X1 port map( A => n4905, Z => n4848);
   U1349 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_29_port, B1 => 
                           n4848, B2 => REGISTERS_23_29_port, ZN => n4238);
   U1350 : NAND4_X1 port map( A1 => n4241, A2 => n4240, A3 => n4239, A4 => 
                           n4238, ZN => n4242);
   U1351 : NOR2_X1 port map( A1 => n4243, A2 => n4242, ZN => n4257);
   U1352 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_6_29_port, B1 => 
                           n4934, B2 => REGISTERS_3_29_port, ZN => n4249);
   U1353 : INV_X1 port map( A => n4244, ZN => n4930);
   U1354 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_29_port, B1 => 
                           n4930, B2 => REGISTERS_5_29_port, ZN => n4248);
   U1355 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_1_29_port, B1 => 
                           n4933, B2 => REGISTERS_2_29_port, ZN => n4247);
   U1356 : INV_X1 port map( A => n4245, ZN => n4586);
   U1357 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_29_port, B1 => 
                           n4586, B2 => REGISTERS_7_29_port, ZN => n4246);
   U1358 : NAND4_X1 port map( A1 => n4249, A2 => n4248, A3 => n4247, A4 => 
                           n4246, ZN => n4255);
   U1359 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_29_port, B1 => 
                           n4932, B2 => REGISTERS_15_29_port, ZN => n4253);
   U1360 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_29_port, B1 => 
                           n4934, B2 => REGISTERS_11_29_port, ZN => n4252);
   U1361 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_29_port, B1 => 
                           n4933, B2 => REGISTERS_10_29_port, ZN => n4251);
   U1362 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_29_port, B1 => 
                           n4942, B2 => REGISTERS_9_29_port, ZN => n4250);
   U1363 : NAND4_X1 port map( A1 => n4253, A2 => n4252, A3 => n4251, A4 => 
                           n4250, ZN => n4254);
   U1364 : AOI22_X1 port map( A1 => n4728, A2 => n4255, B1 => n4953, B2 => 
                           n4254, ZN => n4256);
   U1365 : OAI21_X1 port map( B1 => n4958, B2 => n4257, A => n4256, ZN => N446)
                           ;
   U1366 : CLKBUF_X1 port map( A => n4804, Z => n4909);
   U1367 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_28_port, B1 => 
                           n4909, B2 => REGISTERS_17_28_port, ZN => n4261);
   U1368 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_28_port, B1 => 
                           n4850, B2 => REGISTERS_19_28_port, ZN => n4260);
   U1369 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_28_port, B1 => 
                           n4918, B2 => REGISTERS_26_28_port, ZN => n4259);
   U1370 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_28_port, B1 => 
                           n4907, B2 => REGISTERS_25_28_port, ZN => n4258);
   U1371 : NAND4_X1 port map( A1 => n4261, A2 => n4260, A3 => n4259, A4 => 
                           n4258, ZN => n4267);
   U1372 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_28_port, B1 => 
                           n4848, B2 => REGISTERS_23_28_port, ZN => n4265);
   U1373 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_28_port, B1 => 
                           n4915, B2 => REGISTERS_27_28_port, ZN => n4264);
   U1374 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_28_port, B1 => 
                           n4921, B2 => REGISTERS_31_28_port, ZN => n4263);
   U1375 : AOI22_X1 port map( A1 => n4754, A2 => REGISTERS_30_28_port, B1 => 
                           n4917, B2 => REGISTERS_18_28_port, ZN => n4262);
   U1376 : NAND4_X1 port map( A1 => n4265, A2 => n4264, A3 => n4263, A4 => 
                           n4262, ZN => n4266);
   U1377 : NOR2_X1 port map( A1 => n4267, A2 => n4266, ZN => n4280);
   U1378 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_6_28_port, B1 => 
                           n4741, B2 => REGISTERS_3_28_port, ZN => n4272);
   U1379 : INV_X1 port map( A => n4268, ZN => n4867);
   U1380 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_4_28_port, B1 => 
                           n4931, B2 => REGISTERS_1_28_port, ZN => n4271);
   U1381 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_28_port, B1 => 
                           n4940, B2 => REGISTERS_5_28_port, ZN => n4270);
   U1382 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_28_port, B1 => 
                           n4944, B2 => REGISTERS_7_28_port, ZN => n4269);
   U1383 : NAND4_X1 port map( A1 => n4272, A2 => n4271, A3 => n4270, A4 => 
                           n4269, ZN => n4278);
   U1384 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_28_port, B1 => 
                           n4944, B2 => REGISTERS_15_28_port, ZN => n4276);
   U1385 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_28_port, B1 => 
                           n4815, B2 => REGISTERS_9_28_port, ZN => n4275);
   U1386 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_28_port, B1 => 
                           n4934, B2 => REGISTERS_11_28_port, ZN => n4274);
   U1387 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_28_port, B1 => 
                           n4933, B2 => REGISTERS_10_28_port, ZN => n4273);
   U1388 : NAND4_X1 port map( A1 => n4276, A2 => n4275, A3 => n4274, A4 => 
                           n4273, ZN => n4277);
   U1389 : AOI22_X1 port map( A1 => n4728, A2 => n4278, B1 => n4953, B2 => 
                           n4277, ZN => n4279);
   U1390 : OAI21_X1 port map( B1 => n4958, B2 => n4280, A => n4279, ZN => N445)
                           ;
   U1391 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_27_port, B1 => 
                           n4848, B2 => REGISTERS_23_27_port, ZN => n4284);
   U1392 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_27_port, B1 => 
                           n4907, B2 => REGISTERS_25_27_port, ZN => n4283);
   U1393 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_27_port, B1 => 
                           n4918, B2 => REGISTERS_26_27_port, ZN => n4282);
   U1394 : AOI22_X1 port map( A1 => n4849, A2 => REGISTERS_20_27_port, B1 => 
                           n4919, B2 => REGISTERS_30_27_port, ZN => n4281);
   U1395 : NAND4_X1 port map( A1 => n4284, A2 => n4283, A3 => n4282, A4 => 
                           n4281, ZN => n4290);
   U1396 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_27_port, B1 => 
                           n4621, B2 => REGISTERS_27_27_port, ZN => n4288);
   U1397 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_27_port, B1 => 
                           n4917, B2 => REGISTERS_18_27_port, ZN => n4287);
   U1398 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_27_port, B1 => 
                           n4850, B2 => REGISTERS_19_27_port, ZN => n4286);
   U1399 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_27_port, B1 => 
                           n4909, B2 => REGISTERS_17_27_port, ZN => n4285);
   U1400 : NAND4_X1 port map( A1 => n4288, A2 => n4287, A3 => n4286, A4 => 
                           n4285, ZN => n4289);
   U1401 : NOR2_X1 port map( A1 => n4290, A2 => n4289, ZN => n4303);
   U1402 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_27_port, B1 => 
                           n4932, B2 => REGISTERS_7_27_port, ZN => n4295);
   U1403 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_5_27_port, B1 => 
                           n4934, B2 => REGISTERS_3_27_port, ZN => n4294);
   U1404 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_27_port, B1 => 
                           n4815, B2 => REGISTERS_1_27_port, ZN => n4293);
   U1405 : INV_X1 port map( A => n4291, ZN => n4894);
   U1406 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_27_port, B1 => 
                           n4894, B2 => REGISTERS_6_27_port, ZN => n4292);
   U1407 : NAND4_X1 port map( A1 => n4295, A2 => n4294, A3 => n4293, A4 => 
                           n4292, ZN => n4301);
   U1408 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_27_port, B1 => 
                           n4934, B2 => REGISTERS_11_27_port, ZN => n4299);
   U1409 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_27_port, B1 => 
                           n4815, B2 => REGISTERS_9_27_port, ZN => n4298);
   U1410 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_27_port, B1 => 
                           n4894, B2 => REGISTERS_14_27_port, ZN => n4297);
   U1411 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_10_27_port, B1 => 
                           n4932, B2 => REGISTERS_15_27_port, ZN => n4296);
   U1412 : NAND4_X1 port map( A1 => n4299, A2 => n4298, A3 => n4297, A4 => 
                           n4296, ZN => n4300);
   U1413 : AOI22_X1 port map( A1 => n4728, A2 => n4301, B1 => n4434, B2 => 
                           n4300, ZN => n4302);
   U1414 : OAI21_X1 port map( B1 => n4958, B2 => n4303, A => n4302, ZN => N444)
                           ;
   U1415 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_26_port, B1 => 
                           n4919, B2 => REGISTERS_30_26_port, ZN => n4307);
   U1416 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_26_port, B1 => 
                           n4848, B2 => REGISTERS_23_26_port, ZN => n4306);
   U1417 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_26_port, B1 => 
                           n4917, B2 => REGISTERS_18_26_port, ZN => n4305);
   U1418 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_26_port, B1 => 
                           n4907, B2 => REGISTERS_25_26_port, ZN => n4304);
   U1419 : NAND4_X1 port map( A1 => n4307, A2 => n4306, A3 => n4305, A4 => 
                           n4304, ZN => n4313);
   U1420 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_26_port, B1 => 
                           n4908, B2 => REGISTERS_29_26_port, ZN => n4311);
   U1421 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_26_port, B1 => 
                           n4921, B2 => REGISTERS_31_26_port, ZN => n4310);
   U1422 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_26_port, B1 => 
                           n4849, B2 => REGISTERS_20_26_port, ZN => n4309);
   U1423 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_26_port, B1 => 
                           n4915, B2 => REGISTERS_27_26_port, ZN => n4308);
   U1424 : NAND4_X1 port map( A1 => n4311, A2 => n4310, A3 => n4309, A4 => 
                           n4308, ZN => n4312);
   U1425 : NOR2_X1 port map( A1 => n4313, A2 => n4312, ZN => n4326);
   U1426 : INV_X1 port map( A => n4314, ZN => n4945);
   U1427 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_26_port, B1 => 
                           n4945, B2 => REGISTERS_3_26_port, ZN => n4318);
   U1428 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_26_port, B1 => 
                           n4586, B2 => REGISTERS_7_26_port, ZN => n4317);
   U1429 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_5_26_port, B1 => 
                           n4947, B2 => REGISTERS_6_26_port, ZN => n4316);
   U1430 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_26_port, B1 => 
                           n4933, B2 => REGISTERS_2_26_port, ZN => n4315);
   U1431 : NAND4_X1 port map( A1 => n4318, A2 => n4317, A3 => n4316, A4 => 
                           n4315, ZN => n4324);
   U1432 : AOI22_X1 port map( A1 => n4945, A2 => REGISTERS_11_26_port, B1 => 
                           n4586, B2 => REGISTERS_15_26_port, ZN => n4322);
   U1433 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_12_26_port, B1 => 
                           n4933, B2 => REGISTERS_10_26_port, ZN => n4321);
   U1434 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_26_port, B1 => 
                           n4815, B2 => REGISTERS_9_26_port, ZN => n4320);
   U1435 : CLKBUF_X1 port map( A => n4941, Z => n4935);
   U1436 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_26_port, B1 => 
                           n4894, B2 => REGISTERS_14_26_port, ZN => n4319);
   U1437 : NAND4_X1 port map( A1 => n4322, A2 => n4321, A3 => n4320, A4 => 
                           n4319, ZN => n4323);
   U1438 : AOI22_X1 port map( A1 => n4728, A2 => n4324, B1 => n4434, B2 => 
                           n4323, ZN => n4325);
   U1439 : OAI21_X1 port map( B1 => n4958, B2 => n4326, A => n4325, ZN => N443)
                           ;
   U1440 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_25_port, B1 => 
                           n4849, B2 => REGISTERS_20_25_port, ZN => n4330);
   U1441 : CLKBUF_X1 port map( A => n4442, Z => n4904);
   U1442 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_25_port, B1 => 
                           n4917, B2 => REGISTERS_18_25_port, ZN => n4329);
   U1443 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_25_port, B1 => 
                           n4848, B2 => REGISTERS_23_25_port, ZN => n4328);
   U1444 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_25_port, B1 => 
                           n4907, B2 => REGISTERS_25_25_port, ZN => n4327);
   U1445 : NAND4_X1 port map( A1 => n4330, A2 => n4329, A3 => n4328, A4 => 
                           n4327, ZN => n4336);
   U1446 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_25_port, B1 => 
                           n4850, B2 => REGISTERS_19_25_port, ZN => n4334);
   U1447 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_25_port, B1 => 
                           n4921, B2 => REGISTERS_31_25_port, ZN => n4333);
   U1448 : AOI22_X1 port map( A1 => n4754, A2 => REGISTERS_30_25_port, B1 => 
                           n4621, B2 => REGISTERS_27_25_port, ZN => n4332);
   U1449 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_25_port, B1 => 
                           n4918, B2 => REGISTERS_26_25_port, ZN => n4331);
   U1450 : NAND4_X1 port map( A1 => n4334, A2 => n4333, A3 => n4332, A4 => 
                           n4331, ZN => n4335);
   U1451 : NOR2_X1 port map( A1 => n4336, A2 => n4335, ZN => n4348);
   U1452 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_6_25_port, B1 => 
                           n4933, B2 => REGISTERS_2_25_port, ZN => n4340);
   U1453 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_1_25_port, B1 => 
                           n4586, B2 => REGISTERS_7_25_port, ZN => n4339);
   U1454 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_4_25_port, B1 => 
                           n4741, B2 => REGISTERS_3_25_port, ZN => n4338);
   U1455 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_25_port, B1 => 
                           n4721, B2 => REGISTERS_5_25_port, ZN => n4337);
   U1456 : NAND4_X1 port map( A1 => n4340, A2 => n4339, A3 => n4338, A4 => 
                           n4337, ZN => n4346);
   U1457 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_25_port, B1 => 
                           n4945, B2 => REGISTERS_11_25_port, ZN => n4344);
   U1458 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_25_port, B1 => 
                           n4586, B2 => REGISTERS_15_25_port, ZN => n4343);
   U1459 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_25_port, B1 => 
                           n4815, B2 => REGISTERS_9_25_port, ZN => n4342);
   U1460 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_25_port, B1 => 
                           n4933, B2 => REGISTERS_10_25_port, ZN => n4341);
   U1461 : NAND4_X1 port map( A1 => n4344, A2 => n4343, A3 => n4342, A4 => 
                           n4341, ZN => n4345);
   U1462 : AOI22_X1 port map( A1 => n4728, A2 => n4346, B1 => n4434, B2 => 
                           n4345, ZN => n4347);
   U1463 : OAI21_X1 port map( B1 => n4958, B2 => n4348, A => n4347, ZN => N442)
                           ;
   U1464 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_24_port, B1 => 
                           n4848, B2 => REGISTERS_23_24_port, ZN => n4352);
   U1465 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_24_port, B1 => 
                           n4907, B2 => REGISTERS_25_24_port, ZN => n4351);
   U1466 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_24_port, B1 => 
                           n4918, B2 => REGISTERS_26_24_port, ZN => n4350);
   U1467 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_24_port, B1 => 
                           n4850, B2 => REGISTERS_19_24_port, ZN => n4349);
   U1468 : NAND4_X1 port map( A1 => n4352, A2 => n4351, A3 => n4350, A4 => 
                           n4349, ZN => n4358);
   U1469 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_24_port, B1 => 
                           n4621, B2 => REGISTERS_27_24_port, ZN => n4356);
   U1470 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_24_port, B1 => 
                           n4849, B2 => REGISTERS_20_24_port, ZN => n4355);
   U1471 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_24_port, B1 => 
                           n4754, B2 => REGISTERS_30_24_port, ZN => n4354);
   U1472 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_24_port, B1 => 
                           n4917, B2 => REGISTERS_18_24_port, ZN => n4353);
   U1473 : NAND4_X1 port map( A1 => n4356, A2 => n4355, A3 => n4354, A4 => 
                           n4353, ZN => n4357);
   U1474 : NOR2_X1 port map( A1 => n4358, A2 => n4357, ZN => n4370);
   U1475 : AOI22_X1 port map( A1 => n4934, A2 => REGISTERS_3_24_port, B1 => 
                           n4586, B2 => REGISTERS_7_24_port, ZN => n4362);
   U1476 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_24_port, B1 => 
                           n4815, B2 => REGISTERS_1_24_port, ZN => n4361);
   U1477 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_24_port, B1 => 
                           n4894, B2 => REGISTERS_6_24_port, ZN => n4360);
   U1478 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_24_port, B1 => 
                           n4933, B2 => REGISTERS_2_24_port, ZN => n4359);
   U1479 : NAND4_X1 port map( A1 => n4362, A2 => n4361, A3 => n4360, A4 => 
                           n4359, ZN => n4368);
   U1480 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_24_port, B1 => 
                           n4815, B2 => REGISTERS_9_24_port, ZN => n4366);
   U1481 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_24_port, B1 => 
                           n4934, B2 => REGISTERS_11_24_port, ZN => n4365);
   U1482 : CLKBUF_X1 port map( A => n4933, Z => n4946);
   U1483 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_24_port, B1 => 
                           n4946, B2 => REGISTERS_10_24_port, ZN => n4364);
   U1484 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_24_port, B1 => 
                           n4586, B2 => REGISTERS_15_24_port, ZN => n4363);
   U1485 : NAND4_X1 port map( A1 => n4366, A2 => n4365, A3 => n4364, A4 => 
                           n4363, ZN => n4367);
   U1486 : AOI22_X1 port map( A1 => n4728, A2 => n4368, B1 => n4434, B2 => 
                           n4367, ZN => n4369);
   U1487 : OAI21_X1 port map( B1 => n4958, B2 => n4370, A => n4369, ZN => N441)
                           ;
   U1488 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_23_port, B1 => 
                           n4917, B2 => REGISTERS_18_23_port, ZN => n4374);
   U1489 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_23_port, B1 => 
                           n4903, B2 => REGISTERS_16_23_port, ZN => n4373);
   U1490 : AOI22_X1 port map( A1 => n4919, A2 => REGISTERS_30_23_port, B1 => 
                           n4621, B2 => REGISTERS_27_23_port, ZN => n4372);
   U1491 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_23_port, B1 => 
                           n4921, B2 => REGISTERS_31_23_port, ZN => n4371);
   U1492 : NAND4_X1 port map( A1 => n4374, A2 => n4373, A3 => n4372, A4 => 
                           n4371, ZN => n4380);
   U1493 : AOI22_X1 port map( A1 => n4849, A2 => REGISTERS_20_23_port, B1 => 
                           n4907, B2 => REGISTERS_25_23_port, ZN => n4378);
   U1494 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_23_port, B1 => 
                           n4850, B2 => REGISTERS_19_23_port, ZN => n4377);
   U1495 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_23_port, B1 => 
                           n4848, B2 => REGISTERS_23_23_port, ZN => n4376);
   U1496 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_23_port, B1 => 
                           n4910, B2 => REGISTERS_22_23_port, ZN => n4375);
   U1497 : NAND4_X1 port map( A1 => n4378, A2 => n4377, A3 => n4376, A4 => 
                           n4375, ZN => n4379);
   U1498 : NOR2_X1 port map( A1 => n4380, A2 => n4379, ZN => n4392);
   U1499 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_1_23_port, B1 => 
                           n4586, B2 => REGISTERS_7_23_port, ZN => n4384);
   U1500 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_23_port, B1 => 
                           n4933, B2 => REGISTERS_2_23_port, ZN => n4383);
   U1501 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_5_23_port, B1 => 
                           n4945, B2 => REGISTERS_3_23_port, ZN => n4382);
   U1502 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_23_port, B1 => 
                           n4894, B2 => REGISTERS_6_23_port, ZN => n4381);
   U1503 : NAND4_X1 port map( A1 => n4384, A2 => n4383, A3 => n4382, A4 => 
                           n4381, ZN => n4390);
   U1504 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_23_port, B1 => 
                           n4894, B2 => REGISTERS_14_23_port, ZN => n4388);
   U1505 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_23_port, B1 => 
                           n4934, B2 => REGISTERS_11_23_port, ZN => n4387);
   U1506 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_23_port, B1 => 
                           n4815, B2 => REGISTERS_9_23_port, ZN => n4386);
   U1507 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_10_23_port, B1 => 
                           n4586, B2 => REGISTERS_15_23_port, ZN => n4385);
   U1508 : NAND4_X1 port map( A1 => n4388, A2 => n4387, A3 => n4386, A4 => 
                           n4385, ZN => n4389);
   U1509 : AOI22_X1 port map( A1 => n4728, A2 => n4390, B1 => n4434, B2 => 
                           n4389, ZN => n4391);
   U1510 : OAI21_X1 port map( B1 => n4958, B2 => n4392, A => n4391, ZN => N440)
                           ;
   U1511 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_22_port, B1 => 
                           n4919, B2 => REGISTERS_30_22_port, ZN => n4396);
   U1512 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_22_port, B1 => 
                           n4621, B2 => REGISTERS_27_22_port, ZN => n4395);
   U1513 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_22_port, B1 => 
                           n4909, B2 => REGISTERS_17_22_port, ZN => n4394);
   U1514 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_22_port, B1 => 
                           n4917, B2 => REGISTERS_18_22_port, ZN => n4393);
   U1515 : NAND4_X1 port map( A1 => n4396, A2 => n4395, A3 => n4394, A4 => 
                           n4393, ZN => n4402);
   U1516 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_22_port, B1 => 
                           n4907, B2 => REGISTERS_25_22_port, ZN => n4400);
   U1517 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_22_port, B1 => 
                           n4916, B2 => REGISTERS_21_22_port, ZN => n4399);
   U1518 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_22_port, B1 => 
                           n4848, B2 => REGISTERS_23_22_port, ZN => n4398);
   U1519 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_22_port, B1 => 
                           n4850, B2 => REGISTERS_19_22_port, ZN => n4397);
   U1520 : NAND4_X1 port map( A1 => n4400, A2 => n4399, A3 => n4398, A4 => 
                           n4397, ZN => n4401);
   U1521 : NOR2_X1 port map( A1 => n4402, A2 => n4401, ZN => n4414);
   U1522 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_22_port, B1 => 
                           n4815, B2 => REGISTERS_1_22_port, ZN => n4406);
   U1523 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_5_22_port, B1 => 
                           n4929, B2 => REGISTERS_6_22_port, ZN => n4405);
   U1524 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_22_port, B1 => 
                           n4741, B2 => REGISTERS_3_22_port, ZN => n4404);
   U1525 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_22_port, B1 => 
                           n4586, B2 => REGISTERS_7_22_port, ZN => n4403);
   U1526 : NAND4_X1 port map( A1 => n4406, A2 => n4405, A3 => n4404, A4 => 
                           n4403, ZN => n4412);
   U1527 : AOI22_X1 port map( A1 => n4945, A2 => REGISTERS_11_22_port, B1 => 
                           n4586, B2 => REGISTERS_15_22_port, ZN => n4410);
   U1528 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_22_port, B1 => 
                           n4867, B2 => REGISTERS_12_22_port, ZN => n4409);
   U1529 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_9_22_port, B1 => 
                           n4933, B2 => REGISTERS_10_22_port, ZN => n4408);
   U1530 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_22_port, B1 => 
                           n4894, B2 => REGISTERS_14_22_port, ZN => n4407);
   U1531 : NAND4_X1 port map( A1 => n4410, A2 => n4409, A3 => n4408, A4 => 
                           n4407, ZN => n4411);
   U1532 : AOI22_X1 port map( A1 => n4728, A2 => n4412, B1 => n4434, B2 => 
                           n4411, ZN => n4413);
   U1533 : OAI21_X1 port map( B1 => n4958, B2 => n4414, A => n4413, ZN => N439)
                           ;
   U1534 : AOI22_X1 port map( A1 => n4907, A2 => REGISTERS_25_21_port, B1 => 
                           n4917, B2 => REGISTERS_18_21_port, ZN => n4418);
   U1535 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_21_port, B1 => 
                           n4621, B2 => REGISTERS_27_21_port, ZN => n4417);
   U1536 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_21_port, B1 => 
                           n4909, B2 => REGISTERS_17_21_port, ZN => n4416);
   U1537 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_21_port, B1 => 
                           n4849, B2 => REGISTERS_20_21_port, ZN => n4415);
   U1538 : NAND4_X1 port map( A1 => n4418, A2 => n4417, A3 => n4416, A4 => 
                           n4415, ZN => n4424);
   U1539 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_21_port, B1 => 
                           n4754, B2 => REGISTERS_30_21_port, ZN => n4422);
   U1540 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_21_port, B1 => 
                           n4850, B2 => REGISTERS_19_21_port, ZN => n4421);
   U1541 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_21_port, B1 => 
                           n4848, B2 => REGISTERS_23_21_port, ZN => n4420);
   U1542 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_21_port, B1 => 
                           n4910, B2 => REGISTERS_22_21_port, ZN => n4419);
   U1543 : NAND4_X1 port map( A1 => n4422, A2 => n4421, A3 => n4420, A4 => 
                           n4419, ZN => n4423);
   U1544 : NOR2_X1 port map( A1 => n4424, A2 => n4423, ZN => n4437);
   U1545 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_21_port, B1 => 
                           n4933, B2 => REGISTERS_2_21_port, ZN => n4428);
   U1546 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_6_21_port, B1 => 
                           n4586, B2 => REGISTERS_7_21_port, ZN => n4427);
   U1547 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_21_port, B1 => 
                           n4816, B2 => REGISTERS_4_21_port, ZN => n4426);
   U1548 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_1_21_port, B1 => 
                           n4934, B2 => REGISTERS_3_21_port, ZN => n4425);
   U1549 : NAND4_X1 port map( A1 => n4428, A2 => n4427, A3 => n4426, A4 => 
                           n4425, ZN => n4435);
   U1550 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_21_port, B1 => 
                           n4929, B2 => REGISTERS_14_21_port, ZN => n4432);
   U1551 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_9_21_port, B1 => 
                           n4933, B2 => REGISTERS_10_21_port, ZN => n4431);
   U1552 : AOI22_X1 port map( A1 => n4940, A2 => REGISTERS_13_21_port, B1 => 
                           n4586, B2 => REGISTERS_15_21_port, ZN => n4430);
   U1553 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_21_port, B1 => 
                           n4934, B2 => REGISTERS_11_21_port, ZN => n4429);
   U1554 : NAND4_X1 port map( A1 => n4432, A2 => n4431, A3 => n4430, A4 => 
                           n4429, ZN => n4433);
   U1555 : AOI22_X1 port map( A1 => n4728, A2 => n4435, B1 => n4434, B2 => 
                           n4433, ZN => n4436);
   U1556 : OAI21_X1 port map( B1 => n4958, B2 => n4437, A => n4436, ZN => N438)
                           ;
   U1557 : AOI22_X1 port map( A1 => n4754, A2 => REGISTERS_30_20_port, B1 => 
                           n4825, B2 => REGISTERS_25_20_port, ZN => n4441);
   U1558 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_20_port, B1 => 
                           n4849, B2 => REGISTERS_20_20_port, ZN => n4440);
   U1559 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_20_port, B1 => 
                           n4916, B2 => REGISTERS_21_20_port, ZN => n4439);
   U1560 : AOI22_X1 port map( A1 => n4850, A2 => REGISTERS_19_20_port, B1 => 
                           n4918, B2 => REGISTERS_26_20_port, ZN => n4438);
   U1561 : NAND4_X1 port map( A1 => n4441, A2 => n4440, A3 => n4439, A4 => 
                           n4438, ZN => n4448);
   U1562 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_20_port, B1 => 
                           n4917, B2 => REGISTERS_18_20_port, ZN => n4446);
   U1563 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_20_port, B1 => 
                           n4915, B2 => REGISTERS_27_20_port, ZN => n4445);
   U1564 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_20_port, B1 => 
                           n4909, B2 => REGISTERS_17_20_port, ZN => n4444);
   U1565 : AOI22_X1 port map( A1 => n4442, A2 => REGISTERS_24_20_port, B1 => 
                           n4848, B2 => REGISTERS_23_20_port, ZN => n4443);
   U1566 : NAND4_X1 port map( A1 => n4446, A2 => n4445, A3 => n4444, A4 => 
                           n4443, ZN => n4447);
   U1567 : NOR2_X1 port map( A1 => n4448, A2 => n4447, ZN => n4460);
   U1568 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_20_port, B1 => 
                           n4894, B2 => REGISTERS_6_20_port, ZN => n4452);
   U1569 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_20_port, B1 => 
                           n4586, B2 => REGISTERS_7_20_port, ZN => n4451);
   U1570 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_1_20_port, B1 => 
                           n4933, B2 => REGISTERS_2_20_port, ZN => n4450);
   U1571 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_20_port, B1 => 
                           n4741, B2 => REGISTERS_3_20_port, ZN => n4449);
   U1572 : NAND4_X1 port map( A1 => n4452, A2 => n4451, A3 => n4450, A4 => 
                           n4449, ZN => n4458);
   U1573 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_20_port, B1 => 
                           n4586, B2 => REGISTERS_15_20_port, ZN => n4456);
   U1574 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_20_port, B1 => 
                           n4867, B2 => REGISTERS_12_20_port, ZN => n4455);
   U1575 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_20_port, B1 => 
                           n4741, B2 => REGISTERS_11_20_port, ZN => n4454);
   U1576 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_20_port, B1 => 
                           n4946, B2 => REGISTERS_10_20_port, ZN => n4453);
   U1577 : NAND4_X1 port map( A1 => n4456, A2 => n4455, A3 => n4454, A4 => 
                           n4453, ZN => n4457);
   U1578 : AOI22_X1 port map( A1 => n4728, A2 => n4458, B1 => n4953, B2 => 
                           n4457, ZN => n4459);
   U1579 : OAI21_X1 port map( B1 => n4958, B2 => n4460, A => n4459, ZN => N437)
                           ;
   U1580 : AOI22_X1 port map( A1 => n4919, A2 => REGISTERS_30_19_port, B1 => 
                           n4915, B2 => REGISTERS_27_19_port, ZN => n4464);
   U1581 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_19_port, B1 => 
                           n4917, B2 => REGISTERS_18_19_port, ZN => n4463);
   U1582 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_19_port, B1 => 
                           n4849, B2 => REGISTERS_20_19_port, ZN => n4462);
   U1583 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_19_port, B1 => 
                           n4903, B2 => REGISTERS_16_19_port, ZN => n4461);
   U1584 : NAND4_X1 port map( A1 => n4464, A2 => n4463, A3 => n4462, A4 => 
                           n4461, ZN => n4470);
   U1585 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_19_port, B1 => 
                           n4918, B2 => REGISTERS_26_19_port, ZN => n4468);
   U1586 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_19_port, B1 => 
                           n4804, B2 => REGISTERS_17_19_port, ZN => n4467);
   U1587 : AOI22_X1 port map( A1 => n4825, A2 => REGISTERS_25_19_port, B1 => 
                           n4848, B2 => REGISTERS_23_19_port, ZN => n4466);
   U1588 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_19_port, B1 => 
                           n4850, B2 => REGISTERS_19_19_port, ZN => n4465);
   U1589 : NAND4_X1 port map( A1 => n4468, A2 => n4467, A3 => n4466, A4 => 
                           n4465, ZN => n4469);
   U1590 : NOR2_X1 port map( A1 => n4470, A2 => n4469, ZN => n4482);
   U1591 : CLKBUF_X1 port map( A => n4503, Z => n4955);
   U1592 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_19_port, B1 => 
                           n4944, B2 => REGISTERS_7_19_port, ZN => n4474);
   U1593 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_19_port, B1 => 
                           n4933, B2 => REGISTERS_2_19_port, ZN => n4473);
   U1594 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_19_port, B1 => 
                           n4929, B2 => REGISTERS_6_19_port, ZN => n4472);
   U1595 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_1_19_port, B1 => 
                           n4741, B2 => REGISTERS_3_19_port, ZN => n4471);
   U1596 : NAND4_X1 port map( A1 => n4474, A2 => n4473, A3 => n4472, A4 => 
                           n4471, ZN => n4480);
   U1597 : AOI22_X1 port map( A1 => n4741, A2 => REGISTERS_11_19_port, B1 => 
                           n4586, B2 => REGISTERS_15_19_port, ZN => n4478);
   U1598 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_19_port, B1 => 
                           n4815, B2 => REGISTERS_9_19_port, ZN => n4477);
   U1599 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_19_port, B1 => 
                           n4867, B2 => REGISTERS_12_19_port, ZN => n4476);
   U1600 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_19_port, B1 => 
                           n4933, B2 => REGISTERS_10_19_port, ZN => n4475);
   U1601 : NAND4_X1 port map( A1 => n4478, A2 => n4477, A3 => n4476, A4 => 
                           n4475, ZN => n4479);
   U1602 : AOI22_X1 port map( A1 => n4955, A2 => n4480, B1 => n4953, B2 => 
                           n4479, ZN => n4481);
   U1603 : OAI21_X1 port map( B1 => n4958, B2 => n4482, A => n4481, ZN => N436)
                           ;
   U1604 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_18_port, B1 => 
                           n4921, B2 => REGISTERS_31_18_port, ZN => n4486);
   U1605 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_18_port, B1 => 
                           n4919, B2 => REGISTERS_30_18_port, ZN => n4485);
   U1606 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_18_port, B1 => 
                           n4916, B2 => REGISTERS_21_18_port, ZN => n4484);
   U1607 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_18_port, B1 => 
                           n4910, B2 => REGISTERS_22_18_port, ZN => n4483);
   U1608 : NAND4_X1 port map( A1 => n4486, A2 => n4485, A3 => n4484, A4 => 
                           n4483, ZN => n4492);
   U1609 : AOI22_X1 port map( A1 => n4850, A2 => REGISTERS_19_18_port, B1 => 
                           n4848, B2 => REGISTERS_23_18_port, ZN => n4490);
   U1610 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_18_port, B1 => 
                           n4804, B2 => REGISTERS_17_18_port, ZN => n4489);
   U1611 : AOI22_X1 port map( A1 => n4849, A2 => REGISTERS_20_18_port, B1 => 
                           n4917, B2 => REGISTERS_18_18_port, ZN => n4488);
   U1612 : AOI22_X1 port map( A1 => n4825, A2 => REGISTERS_25_18_port, B1 => 
                           n4621, B2 => REGISTERS_27_18_port, ZN => n4487);
   U1613 : NAND4_X1 port map( A1 => n4490, A2 => n4489, A3 => n4488, A4 => 
                           n4487, ZN => n4491);
   U1614 : NOR2_X1 port map( A1 => n4492, A2 => n4491, ZN => n4505);
   U1615 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_18_port, B1 => 
                           n4940, B2 => REGISTERS_5_18_port, ZN => n4496);
   U1616 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_1_18_port, B1 => 
                           n4932, B2 => REGISTERS_7_18_port, ZN => n4495);
   U1617 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_6_18_port, B1 => 
                           n4741, B2 => REGISTERS_3_18_port, ZN => n4494);
   U1618 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_18_port, B1 => 
                           n4933, B2 => REGISTERS_2_18_port, ZN => n4493);
   U1619 : NAND4_X1 port map( A1 => n4496, A2 => n4495, A3 => n4494, A4 => 
                           n4493, ZN => n4502);
   U1620 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_18_port, B1 => 
                           n4944, B2 => REGISTERS_15_18_port, ZN => n4500);
   U1621 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_18_port, B1 => 
                           n4867, B2 => REGISTERS_12_18_port, ZN => n4499);
   U1622 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_18_port, B1 => 
                           n4946, B2 => REGISTERS_10_18_port, ZN => n4498);
   U1623 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_18_port, B1 => 
                           n4741, B2 => REGISTERS_11_18_port, ZN => n4497);
   U1624 : NAND4_X1 port map( A1 => n4500, A2 => n4499, A3 => n4498, A4 => 
                           n4497, ZN => n4501);
   U1625 : AOI22_X1 port map( A1 => n4503, A2 => n4502, B1 => n4953, B2 => 
                           n4501, ZN => n4504);
   U1626 : OAI21_X1 port map( B1 => n4958, B2 => n4505, A => n4504, ZN => N435)
                           ;
   U1627 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_17_port, B1 => 
                           n4825, B2 => REGISTERS_25_17_port, ZN => n4509);
   U1628 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_17_port, B1 => 
                           n4849, B2 => REGISTERS_20_17_port, ZN => n4508);
   U1629 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_17_port, B1 => 
                           n4919, B2 => REGISTERS_30_17_port, ZN => n4507);
   U1630 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_17_port, B1 => 
                           n4915, B2 => REGISTERS_27_17_port, ZN => n4506);
   U1631 : NAND4_X1 port map( A1 => n4509, A2 => n4508, A3 => n4507, A4 => 
                           n4506, ZN => n4515);
   U1632 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_17_port, B1 => 
                           n4917, B2 => REGISTERS_18_17_port, ZN => n4513);
   U1633 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_17_port, B1 => 
                           n4918, B2 => REGISTERS_26_17_port, ZN => n4512);
   U1634 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_17_port, B1 => 
                           n4922, B2 => REGISTERS_28_17_port, ZN => n4511);
   U1635 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_17_port, B1 => 
                           n4848, B2 => REGISTERS_23_17_port, ZN => n4510);
   U1636 : NAND4_X1 port map( A1 => n4513, A2 => n4512, A3 => n4511, A4 => 
                           n4510, ZN => n4514);
   U1637 : NOR2_X1 port map( A1 => n4515, A2 => n4514, ZN => n4527);
   U1638 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_4_17_port, B1 => 
                           n4932, B2 => REGISTERS_7_17_port, ZN => n4519);
   U1639 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_17_port, B1 => 
                           n4929, B2 => REGISTERS_6_17_port, ZN => n4518);
   U1640 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_17_port, B1 => 
                           n4946, B2 => REGISTERS_2_17_port, ZN => n4517);
   U1641 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_17_port, B1 => 
                           n4741, B2 => REGISTERS_3_17_port, ZN => n4516);
   U1642 : NAND4_X1 port map( A1 => n4519, A2 => n4518, A3 => n4517, A4 => 
                           n4516, ZN => n4525);
   U1643 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_17_port, B1 => 
                           n4816, B2 => REGISTERS_12_17_port, ZN => n4523);
   U1644 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_17_port, B1 => 
                           n4741, B2 => REGISTERS_11_17_port, ZN => n4522);
   U1645 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_17_port, B1 => 
                           n4933, B2 => REGISTERS_10_17_port, ZN => n4521);
   U1646 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_9_17_port, B1 => 
                           n4932, B2 => REGISTERS_15_17_port, ZN => n4520);
   U1647 : NAND4_X1 port map( A1 => n4523, A2 => n4522, A3 => n4521, A4 => 
                           n4520, ZN => n4524);
   U1648 : AOI22_X1 port map( A1 => n4955, A2 => n4525, B1 => n4953, B2 => 
                           n4524, ZN => n4526);
   U1649 : OAI21_X1 port map( B1 => n4958, B2 => n4527, A => n4526, ZN => N434)
                           ;
   U1650 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_16_port, B1 => 
                           n4849, B2 => REGISTERS_20_16_port, ZN => n4531);
   U1651 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_16_port, B1 => 
                           n4917, B2 => REGISTERS_18_16_port, ZN => n4530);
   U1652 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_16_port, B1 => 
                           n4907, B2 => REGISTERS_25_16_port, ZN => n4529);
   U1653 : AOI22_X1 port map( A1 => n4754, A2 => REGISTERS_30_16_port, B1 => 
                           n4915, B2 => REGISTERS_27_16_port, ZN => n4528);
   U1654 : NAND4_X1 port map( A1 => n4531, A2 => n4530, A3 => n4529, A4 => 
                           n4528, ZN => n4537);
   U1655 : AOI22_X1 port map( A1 => n4850, A2 => REGISTERS_19_16_port, B1 => 
                           n4905, B2 => REGISTERS_23_16_port, ZN => n4535);
   U1656 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_16_port, B1 => 
                           n4918, B2 => REGISTERS_26_16_port, ZN => n4534);
   U1657 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_16_port, B1 => 
                           n4710, B2 => REGISTERS_31_16_port, ZN => n4533);
   U1658 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_16_port, B1 => 
                           n4910, B2 => REGISTERS_22_16_port, ZN => n4532);
   U1659 : NAND4_X1 port map( A1 => n4535, A2 => n4534, A3 => n4533, A4 => 
                           n4532, ZN => n4536);
   U1660 : NOR2_X1 port map( A1 => n4537, A2 => n4536, ZN => n4549);
   U1661 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_16_port, B1 => 
                           n4741, B2 => REGISTERS_3_16_port, ZN => n4541);
   U1662 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_16_port, B1 => 
                           n4586, B2 => REGISTERS_7_16_port, ZN => n4540);
   U1663 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_16_port, B1 => 
                           n4933, B2 => REGISTERS_2_16_port, ZN => n4539);
   U1664 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_16_port, B1 => 
                           n4894, B2 => REGISTERS_6_16_port, ZN => n4538);
   U1665 : NAND4_X1 port map( A1 => n4541, A2 => n4540, A3 => n4539, A4 => 
                           n4538, ZN => n4547);
   U1666 : AOI22_X1 port map( A1 => n4945, A2 => REGISTERS_11_16_port, B1 => 
                           n4933, B2 => REGISTERS_10_16_port, ZN => n4545);
   U1667 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_12_16_port, B1 => 
                           n4894, B2 => REGISTERS_14_16_port, ZN => n4544);
   U1668 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_16_port, B1 => 
                           n4815, B2 => REGISTERS_9_16_port, ZN => n4543);
   U1669 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_16_port, B1 => 
                           n4586, B2 => REGISTERS_15_16_port, ZN => n4542);
   U1670 : NAND4_X1 port map( A1 => n4545, A2 => n4544, A3 => n4543, A4 => 
                           n4542, ZN => n4546);
   U1671 : AOI22_X1 port map( A1 => n4728, A2 => n4547, B1 => n4953, B2 => 
                           n4546, ZN => n4548);
   U1672 : OAI21_X1 port map( B1 => n4958, B2 => n4549, A => n4548, ZN => N433)
                           ;
   U1673 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_15_port, B1 => 
                           n4916, B2 => REGISTERS_21_15_port, ZN => n4553);
   U1674 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_15_port, B1 => 
                           n4905, B2 => REGISTERS_23_15_port, ZN => n4552);
   U1675 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_15_port, B1 => 
                           n4919, B2 => REGISTERS_30_15_port, ZN => n4551);
   U1676 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_15_port, B1 => 
                           n4907, B2 => REGISTERS_25_15_port, ZN => n4550);
   U1677 : NAND4_X1 port map( A1 => n4553, A2 => n4552, A3 => n4551, A4 => 
                           n4550, ZN => n4559);
   U1678 : AOI22_X1 port map( A1 => n4849, A2 => REGISTERS_20_15_port, B1 => 
                           n4621, B2 => REGISTERS_27_15_port, ZN => n4557);
   U1679 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_15_port, B1 => 
                           n4803, B2 => REGISTERS_26_15_port, ZN => n4556);
   U1680 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_15_port, B1 => 
                           n4917, B2 => REGISTERS_18_15_port, ZN => n4555);
   U1681 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_15_port, B1 => 
                           n4920, B2 => REGISTERS_19_15_port, ZN => n4554);
   U1682 : NAND4_X1 port map( A1 => n4557, A2 => n4556, A3 => n4555, A4 => 
                           n4554, ZN => n4558);
   U1683 : NOR2_X1 port map( A1 => n4559, A2 => n4558, ZN => n4571);
   U1684 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_15_port, B1 => 
                           n4815, B2 => REGISTERS_1_15_port, ZN => n4563);
   U1685 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_15_port, B1 => 
                           n4940, B2 => REGISTERS_5_15_port, ZN => n4562);
   U1686 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_6_15_port, B1 => 
                           n4946, B2 => REGISTERS_2_15_port, ZN => n4561);
   U1687 : AOI22_X1 port map( A1 => n4741, A2 => REGISTERS_3_15_port, B1 => 
                           n4944, B2 => REGISTERS_7_15_port, ZN => n4560);
   U1688 : NAND4_X1 port map( A1 => n4563, A2 => n4562, A3 => n4561, A4 => 
                           n4560, ZN => n4569);
   U1689 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_15_port, B1 => 
                           n4586, B2 => REGISTERS_15_15_port, ZN => n4567);
   U1690 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_15_port, B1 => 
                           n4815, B2 => REGISTERS_9_15_port, ZN => n4566);
   U1691 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_12_15_port, B1 => 
                           n4933, B2 => REGISTERS_10_15_port, ZN => n4565);
   U1692 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_15_port, B1 => 
                           n4741, B2 => REGISTERS_11_15_port, ZN => n4564);
   U1693 : NAND4_X1 port map( A1 => n4567, A2 => n4566, A3 => n4565, A4 => 
                           n4564, ZN => n4568);
   U1694 : AOI22_X1 port map( A1 => n4955, A2 => n4569, B1 => n4953, B2 => 
                           n4568, ZN => n4570);
   U1695 : OAI21_X1 port map( B1 => n4958, B2 => n4571, A => n4570, ZN => N432)
                           ;
   U1696 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_14_port, B1 => 
                           n4916, B2 => REGISTERS_21_14_port, ZN => n4575);
   U1697 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_14_port, B1 => 
                           n4918, B2 => REGISTERS_26_14_port, ZN => n4574);
   U1698 : AOI22_X1 port map( A1 => n4882, A2 => REGISTERS_18_14_port, B1 => 
                           n4915, B2 => REGISTERS_27_14_port, ZN => n4573);
   U1699 : AOI22_X1 port map( A1 => n4754, A2 => REGISTERS_30_14_port, B1 => 
                           n4848, B2 => REGISTERS_23_14_port, ZN => n4572);
   U1700 : NAND4_X1 port map( A1 => n4575, A2 => n4574, A3 => n4573, A4 => 
                           n4572, ZN => n4581);
   U1701 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_14_port, B1 => 
                           n4920, B2 => REGISTERS_19_14_port, ZN => n4579);
   U1702 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_14_port, B1 => 
                           n4907, B2 => REGISTERS_25_14_port, ZN => n4578);
   U1703 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_14_port, B1 => 
                           n4710, B2 => REGISTERS_31_14_port, ZN => n4577);
   U1704 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_14_port, B1 => 
                           n4906, B2 => REGISTERS_20_14_port, ZN => n4576);
   U1705 : NAND4_X1 port map( A1 => n4579, A2 => n4578, A3 => n4577, A4 => 
                           n4576, ZN => n4580);
   U1706 : NOR2_X1 port map( A1 => n4581, A2 => n4580, ZN => n4594);
   U1707 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_14_port, B1 => 
                           n4946, B2 => REGISTERS_2_14_port, ZN => n4585);
   U1708 : AOI22_X1 port map( A1 => n4934, A2 => REGISTERS_3_14_port, B1 => 
                           n4586, B2 => REGISTERS_7_14_port, ZN => n4584);
   U1709 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_14_port, B1 => 
                           n4940, B2 => REGISTERS_5_14_port, ZN => n4583);
   U1710 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_4_14_port, B1 => 
                           n4894, B2 => REGISTERS_6_14_port, ZN => n4582);
   U1711 : NAND4_X1 port map( A1 => n4585, A2 => n4584, A3 => n4583, A4 => 
                           n4582, ZN => n4592);
   U1712 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_14_port, B1 => 
                           n4946, B2 => REGISTERS_10_14_port, ZN => n4590);
   U1713 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_14_port, B1 => 
                           n4931, B2 => REGISTERS_9_14_port, ZN => n4589);
   U1714 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_14_port, B1 => 
                           n4867, B2 => REGISTERS_12_14_port, ZN => n4588);
   U1715 : AOI22_X1 port map( A1 => n4934, A2 => REGISTERS_11_14_port, B1 => 
                           n4586, B2 => REGISTERS_15_14_port, ZN => n4587);
   U1716 : NAND4_X1 port map( A1 => n4590, A2 => n4589, A3 => n4588, A4 => 
                           n4587, ZN => n4591);
   U1717 : AOI22_X1 port map( A1 => n4728, A2 => n4592, B1 => n4953, B2 => 
                           n4591, ZN => n4593);
   U1718 : OAI21_X1 port map( B1 => n4958, B2 => n4594, A => n4593, ZN => N431)
                           ;
   U1719 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_13_port, B1 => 
                           n4909, B2 => REGISTERS_17_13_port, ZN => n4598);
   U1720 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_13_port, B1 => 
                           n4850, B2 => REGISTERS_19_13_port, ZN => n4597);
   U1721 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_13_port, B1 => 
                           n4849, B2 => REGISTERS_20_13_port, ZN => n4596);
   U1722 : AOI22_X1 port map( A1 => n4848, A2 => REGISTERS_23_13_port, B1 => 
                           n4621, B2 => REGISTERS_27_13_port, ZN => n4595);
   U1723 : NAND4_X1 port map( A1 => n4598, A2 => n4597, A3 => n4596, A4 => 
                           n4595, ZN => n4604);
   U1724 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_13_port, B1 => 
                           n4921, B2 => REGISTERS_31_13_port, ZN => n4602);
   U1725 : AOI22_X1 port map( A1 => n4919, A2 => REGISTERS_30_13_port, B1 => 
                           n4907, B2 => REGISTERS_25_13_port, ZN => n4601);
   U1726 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_13_port, B1 => 
                           n4803, B2 => REGISTERS_26_13_port, ZN => n4600);
   U1727 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_13_port, B1 => 
                           n4917, B2 => REGISTERS_18_13_port, ZN => n4599);
   U1728 : NAND4_X1 port map( A1 => n4602, A2 => n4601, A3 => n4600, A4 => 
                           n4599, ZN => n4603);
   U1729 : NOR2_X1 port map( A1 => n4604, A2 => n4603, ZN => n4616);
   U1730 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_13_port, B1 => 
                           n4741, B2 => REGISTERS_3_13_port, ZN => n4608);
   U1731 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_13_port, B1 => 
                           n4894, B2 => REGISTERS_6_13_port, ZN => n4607);
   U1732 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_4_13_port, B1 => 
                           n4944, B2 => REGISTERS_7_13_port, ZN => n4606);
   U1733 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_13_port, B1 => 
                           n4946, B2 => REGISTERS_2_13_port, ZN => n4605);
   U1734 : NAND4_X1 port map( A1 => n4608, A2 => n4607, A3 => n4606, A4 => 
                           n4605, ZN => n4614);
   U1735 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_13_port, B1 => 
                           n4944, B2 => REGISTERS_15_13_port, ZN => n4612);
   U1736 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_13_port, B1 => 
                           n4946, B2 => REGISTERS_10_13_port, ZN => n4611);
   U1737 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_13_port, B1 => 
                           n4894, B2 => REGISTERS_14_13_port, ZN => n4610);
   U1738 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_13_port, B1 => 
                           n4741, B2 => REGISTERS_11_13_port, ZN => n4609);
   U1739 : NAND4_X1 port map( A1 => n4612, A2 => n4611, A3 => n4610, A4 => 
                           n4609, ZN => n4613);
   U1740 : AOI22_X1 port map( A1 => n4728, A2 => n4614, B1 => n4953, B2 => 
                           n4613, ZN => n4615);
   U1741 : OAI21_X1 port map( B1 => n4958, B2 => n4616, A => n4615, ZN => N430)
                           ;
   U1742 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_12_port, B1 => 
                           n4905, B2 => REGISTERS_23_12_port, ZN => n4620);
   U1743 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_12_port, B1 => 
                           n4910, B2 => REGISTERS_22_12_port, ZN => n4619);
   U1744 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_12_port, B1 => 
                           n4849, B2 => REGISTERS_20_12_port, ZN => n4618);
   U1745 : AOI22_X1 port map( A1 => n4919, A2 => REGISTERS_30_12_port, B1 => 
                           n4917, B2 => REGISTERS_18_12_port, ZN => n4617);
   U1746 : NAND4_X1 port map( A1 => n4620, A2 => n4619, A3 => n4618, A4 => 
                           n4617, ZN => n4627);
   U1747 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_12_port, B1 => 
                           n4916, B2 => REGISTERS_21_12_port, ZN => n4625);
   U1748 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_12_port, B1 => 
                           n4907, B2 => REGISTERS_25_12_port, ZN => n4624);
   U1749 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_12_port, B1 => 
                           n4920, B2 => REGISTERS_19_12_port, ZN => n4623);
   U1750 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_12_port, B1 => 
                           n4621, B2 => REGISTERS_27_12_port, ZN => n4622);
   U1751 : NAND4_X1 port map( A1 => n4625, A2 => n4624, A3 => n4623, A4 => 
                           n4622, ZN => n4626);
   U1752 : NOR2_X1 port map( A1 => n4627, A2 => n4626, ZN => n4639);
   U1753 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_12_port, B1 => 
                           n4931, B2 => REGISTERS_1_12_port, ZN => n4631);
   U1754 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_12_port, B1 => 
                           n4944, B2 => REGISTERS_7_12_port, ZN => n4630);
   U1755 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_6_12_port, B1 => 
                           n4946, B2 => REGISTERS_2_12_port, ZN => n4629);
   U1756 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_12_port, B1 => 
                           n4945, B2 => REGISTERS_3_12_port, ZN => n4628);
   U1757 : NAND4_X1 port map( A1 => n4631, A2 => n4630, A3 => n4629, A4 => 
                           n4628, ZN => n4637);
   U1758 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_12_port, B1 => 
                           n4945, B2 => REGISTERS_11_12_port, ZN => n4635);
   U1759 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_12_port, B1 => 
                           n4944, B2 => REGISTERS_15_12_port, ZN => n4634);
   U1760 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_12_port, B1 => 
                           n4931, B2 => REGISTERS_9_12_port, ZN => n4633);
   U1761 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_12_port, B1 => 
                           n4946, B2 => REGISTERS_10_12_port, ZN => n4632);
   U1762 : NAND4_X1 port map( A1 => n4635, A2 => n4634, A3 => n4633, A4 => 
                           n4632, ZN => n4636);
   U1763 : AOI22_X1 port map( A1 => n4728, A2 => n4637, B1 => n4953, B2 => 
                           n4636, ZN => n4638);
   U1764 : OAI21_X1 port map( B1 => n4958, B2 => n4639, A => n4638, ZN => N429)
                           ;
   U1765 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_11_port, B1 => 
                           n4905, B2 => REGISTERS_23_11_port, ZN => n4643);
   U1766 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_11_port, B1 => 
                           n4849, B2 => REGISTERS_20_11_port, ZN => n4642);
   U1767 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_11_port, B1 => 
                           n4915, B2 => REGISTERS_27_11_port, ZN => n4641);
   U1768 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_11_port, B1 => 
                           n4850, B2 => REGISTERS_19_11_port, ZN => n4640);
   U1769 : NAND4_X1 port map( A1 => n4643, A2 => n4642, A3 => n4641, A4 => 
                           n4640, ZN => n4649);
   U1770 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_11_port, B1 => 
                           n4907, B2 => REGISTERS_25_11_port, ZN => n4647);
   U1771 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_11_port, B1 => 
                           n4754, B2 => REGISTERS_30_11_port, ZN => n4646);
   U1772 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_11_port, B1 => 
                           n4710, B2 => REGISTERS_31_11_port, ZN => n4645);
   U1773 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_11_port, B1 => 
                           n4917, B2 => REGISTERS_18_11_port, ZN => n4644);
   U1774 : NAND4_X1 port map( A1 => n4647, A2 => n4646, A3 => n4645, A4 => 
                           n4644, ZN => n4648);
   U1775 : NOR2_X1 port map( A1 => n4649, A2 => n4648, ZN => n4661);
   U1776 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_6_11_port, B1 => 
                           n4945, B2 => REGISTERS_3_11_port, ZN => n4653);
   U1777 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_11_port, B1 => 
                           n4931, B2 => REGISTERS_1_11_port, ZN => n4652);
   U1778 : AOI22_X1 port map( A1 => n4946, A2 => REGISTERS_2_11_port, B1 => 
                           n4944, B2 => REGISTERS_7_11_port, ZN => n4651);
   U1779 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_5_11_port, B1 => 
                           n4867, B2 => REGISTERS_4_11_port, ZN => n4650);
   U1780 : NAND4_X1 port map( A1 => n4653, A2 => n4652, A3 => n4651, A4 => 
                           n4650, ZN => n4659);
   U1781 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_11_port, B1 => 
                           n4944, B2 => REGISTERS_15_11_port, ZN => n4657);
   U1782 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_11_port, B1 => 
                           n4894, B2 => REGISTERS_14_11_port, ZN => n4656);
   U1783 : AOI22_X1 port map( A1 => n4741, A2 => REGISTERS_11_11_port, B1 => 
                           n4946, B2 => REGISTERS_10_11_port, ZN => n4655);
   U1784 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_11_port, B1 => 
                           n4931, B2 => REGISTERS_9_11_port, ZN => n4654);
   U1785 : NAND4_X1 port map( A1 => n4657, A2 => n4656, A3 => n4655, A4 => 
                           n4654, ZN => n4658);
   U1786 : AOI22_X1 port map( A1 => n4728, A2 => n4659, B1 => n4953, B2 => 
                           n4658, ZN => n4660);
   U1787 : OAI21_X1 port map( B1 => n4958, B2 => n4661, A => n4660, ZN => N428)
                           ;
   U1788 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_10_port, B1 => 
                           n4916, B2 => REGISTERS_21_10_port, ZN => n4665);
   U1789 : AOI22_X1 port map( A1 => n4849, A2 => REGISTERS_20_10_port, B1 => 
                           n4907, B2 => REGISTERS_25_10_port, ZN => n4664);
   U1790 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_10_port, B1 => 
                           n4903, B2 => REGISTERS_16_10_port, ZN => n4663);
   U1791 : AOI22_X1 port map( A1 => n4919, A2 => REGISTERS_30_10_port, B1 => 
                           n4905, B2 => REGISTERS_23_10_port, ZN => n4662);
   U1792 : NAND4_X1 port map( A1 => n4665, A2 => n4664, A3 => n4663, A4 => 
                           n4662, ZN => n4671);
   U1793 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_10_port, B1 => 
                           n4915, B2 => REGISTERS_27_10_port, ZN => n4669);
   U1794 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_10_port, B1 => 
                           n4909, B2 => REGISTERS_17_10_port, ZN => n4668);
   U1795 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_10_port, B1 => 
                           n4803, B2 => REGISTERS_26_10_port, ZN => n4667);
   U1796 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_10_port, B1 => 
                           n4882, B2 => REGISTERS_18_10_port, ZN => n4666);
   U1797 : NAND4_X1 port map( A1 => n4669, A2 => n4668, A3 => n4667, A4 => 
                           n4666, ZN => n4670);
   U1798 : NOR2_X1 port map( A1 => n4671, A2 => n4670, ZN => n4683);
   U1799 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_10_port, B1 => 
                           n4946, B2 => REGISTERS_2_10_port, ZN => n4675);
   U1800 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_10_port, B1 => 
                           n4931, B2 => REGISTERS_1_10_port, ZN => n4674);
   U1801 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_10_port, B1 => 
                           n4929, B2 => REGISTERS_6_10_port, ZN => n4673);
   U1802 : AOI22_X1 port map( A1 => n4945, A2 => REGISTERS_3_10_port, B1 => 
                           n4944, B2 => REGISTERS_7_10_port, ZN => n4672);
   U1803 : NAND4_X1 port map( A1 => n4675, A2 => n4674, A3 => n4673, A4 => 
                           n4672, ZN => n4681);
   U1804 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_10_port, B1 => 
                           n4946, B2 => REGISTERS_10_10_port, ZN => n4679);
   U1805 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_10_port, B1 => 
                           n4867, B2 => REGISTERS_12_10_port, ZN => n4678);
   U1806 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_10_port, B1 => 
                           n4945, B2 => REGISTERS_11_10_port, ZN => n4677);
   U1807 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_10_port, B1 => 
                           n4944, B2 => REGISTERS_15_10_port, ZN => n4676);
   U1808 : NAND4_X1 port map( A1 => n4679, A2 => n4678, A3 => n4677, A4 => 
                           n4676, ZN => n4680);
   U1809 : AOI22_X1 port map( A1 => n4728, A2 => n4681, B1 => n4953, B2 => 
                           n4680, ZN => n4682);
   U1810 : OAI21_X1 port map( B1 => n4958, B2 => n4683, A => n4682, ZN => N427)
                           ;
   U1811 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_9_port, B1 => 
                           n4922, B2 => REGISTERS_28_9_port, ZN => n4687);
   U1812 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_9_port, B1 => 
                           n4915, B2 => REGISTERS_27_9_port, ZN => n4686);
   U1813 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_9_port, B1 => 
                           n4907, B2 => REGISTERS_25_9_port, ZN => n4685);
   U1814 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_9_port, B1 => 
                           n4848, B2 => REGISTERS_23_9_port, ZN => n4684);
   U1815 : NAND4_X1 port map( A1 => n4687, A2 => n4686, A3 => n4685, A4 => 
                           n4684, ZN => n4693);
   U1816 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_9_port, B1 => 
                           n4850, B2 => REGISTERS_19_9_port, ZN => n4691);
   U1817 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_9_port, B1 => 
                           n4710, B2 => REGISTERS_31_9_port, ZN => n4690);
   U1818 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_9_port, B1 => 
                           n4754, B2 => REGISTERS_30_9_port, ZN => n4689);
   U1819 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_9_port, B1 => 
                           n4882, B2 => REGISTERS_18_9_port, ZN => n4688);
   U1820 : NAND4_X1 port map( A1 => n4691, A2 => n4690, A3 => n4689, A4 => 
                           n4688, ZN => n4692);
   U1821 : NOR2_X1 port map( A1 => n4693, A2 => n4692, ZN => n4705);
   U1822 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_9_port, B1 => 
                           n4946, B2 => REGISTERS_2_9_port, ZN => n4697);
   U1823 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_9_port, B1 => 
                           n4947, B2 => REGISTERS_6_9_port, ZN => n4696);
   U1824 : AOI22_X1 port map( A1 => n4867, A2 => REGISTERS_4_9_port, B1 => 
                           n4945, B2 => REGISTERS_3_9_port, ZN => n4695);
   U1825 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_9_port, B1 => 
                           n4944, B2 => REGISTERS_7_9_port, ZN => n4694);
   U1826 : NAND4_X1 port map( A1 => n4697, A2 => n4696, A3 => n4695, A4 => 
                           n4694, ZN => n4703);
   U1827 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_9_9_port, B1 => 
                           n4946, B2 => REGISTERS_10_9_port, ZN => n4701);
   U1828 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_9_port, B1 => 
                           n4944, B2 => REGISTERS_15_9_port, ZN => n4700);
   U1829 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_9_port, B1 => 
                           n4945, B2 => REGISTERS_11_9_port, ZN => n4699);
   U1830 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_9_port, B1 => 
                           n4867, B2 => REGISTERS_12_9_port, ZN => n4698);
   U1831 : NAND4_X1 port map( A1 => n4701, A2 => n4700, A3 => n4699, A4 => 
                           n4698, ZN => n4702);
   U1832 : AOI22_X1 port map( A1 => n4728, A2 => n4703, B1 => n4953, B2 => 
                           n4702, ZN => n4704);
   U1833 : OAI21_X1 port map( B1 => n4958, B2 => n4705, A => n4704, ZN => N426)
                           ;
   U1834 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_8_port, B1 => 
                           n4918, B2 => REGISTERS_26_8_port, ZN => n4709);
   U1835 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_8_port, B1 => 
                           n4919, B2 => REGISTERS_30_8_port, ZN => n4708);
   U1836 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_8_port, B1 => 
                           n4850, B2 => REGISTERS_19_8_port, ZN => n4707);
   U1837 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_8_port, B1 => 
                           n4917, B2 => REGISTERS_18_8_port, ZN => n4706);
   U1838 : NAND4_X1 port map( A1 => n4709, A2 => n4708, A3 => n4707, A4 => 
                           n4706, ZN => n4716);
   U1839 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_8_port, B1 => 
                           n4915, B2 => REGISTERS_27_8_port, ZN => n4714);
   U1840 : AOI22_X1 port map( A1 => n4825, A2 => REGISTERS_25_8_port, B1 => 
                           n4905, B2 => REGISTERS_23_8_port, ZN => n4713);
   U1841 : AOI22_X1 port map( A1 => n4903, A2 => REGISTERS_16_8_port, B1 => 
                           n4804, B2 => REGISTERS_17_8_port, ZN => n4712);
   U1842 : AOI22_X1 port map( A1 => n4710, A2 => REGISTERS_31_8_port, B1 => 
                           n4906, B2 => REGISTERS_20_8_port, ZN => n4711);
   U1843 : NAND4_X1 port map( A1 => n4714, A2 => n4713, A3 => n4712, A4 => 
                           n4711, ZN => n4715);
   U1844 : NOR2_X1 port map( A1 => n4716, A2 => n4715, ZN => n4730);
   U1845 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_8_port, B1 => 
                           n4944, B2 => REGISTERS_7_8_port, ZN => n4720);
   U1846 : AOI22_X1 port map( A1 => n4894, A2 => REGISTERS_6_8_port, B1 => 
                           n4946, B2 => REGISTERS_2_8_port, ZN => n4719);
   U1847 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_0_8_port, B1 => 
                           n4931, B2 => REGISTERS_1_8_port, ZN => n4718);
   U1848 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_8_port, B1 => 
                           n4945, B2 => REGISTERS_3_8_port, ZN => n4717);
   U1849 : NAND4_X1 port map( A1 => n4720, A2 => n4719, A3 => n4718, A4 => 
                           n4717, ZN => n4727);
   U1850 : AOI22_X1 port map( A1 => n4721, A2 => REGISTERS_13_8_port, B1 => 
                           n4944, B2 => REGISTERS_15_8_port, ZN => n4725);
   U1851 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_8_port, B1 => 
                           n4933, B2 => REGISTERS_10_8_port, ZN => n4724);
   U1852 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_8_port, B1 => 
                           n4741, B2 => REGISTERS_11_8_port, ZN => n4723);
   U1853 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_8_port, B1 => 
                           n4867, B2 => REGISTERS_12_8_port, ZN => n4722);
   U1854 : NAND4_X1 port map( A1 => n4725, A2 => n4724, A3 => n4723, A4 => 
                           n4722, ZN => n4726);
   U1855 : AOI22_X1 port map( A1 => n4728, A2 => n4727, B1 => n4953, B2 => 
                           n4726, ZN => n4729);
   U1856 : OAI21_X1 port map( B1 => n4958, B2 => n4730, A => n4729, ZN => N425)
                           ;
   U1857 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_7_port, B1 => 
                           n4907, B2 => REGISTERS_25_7_port, ZN => n4734);
   U1858 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_7_port, B1 => 
                           n4882, B2 => REGISTERS_18_7_port, ZN => n4733);
   U1859 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_7_port, B1 => 
                           n4921, B2 => REGISTERS_31_7_port, ZN => n4732);
   U1860 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_7_port, B1 => 
                           n4919, B2 => REGISTERS_30_7_port, ZN => n4731);
   U1861 : NAND4_X1 port map( A1 => n4734, A2 => n4733, A3 => n4732, A4 => 
                           n4731, ZN => n4740);
   U1862 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_7_port, B1 => 
                           n4916, B2 => REGISTERS_21_7_port, ZN => n4738);
   U1863 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_7_port, B1 => 
                           n4905, B2 => REGISTERS_23_7_port, ZN => n4737);
   U1864 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_7_port, B1 => 
                           n4920, B2 => REGISTERS_19_7_port, ZN => n4736);
   U1865 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_7_port, B1 => 
                           n4915, B2 => REGISTERS_27_7_port, ZN => n4735);
   U1866 : NAND4_X1 port map( A1 => n4738, A2 => n4737, A3 => n4736, A4 => 
                           n4735, ZN => n4739);
   U1867 : NOR2_X1 port map( A1 => n4740, A2 => n4739, ZN => n4753);
   U1868 : AOI22_X1 port map( A1 => n4741, A2 => REGISTERS_3_7_port, B1 => 
                           n4932, B2 => REGISTERS_7_7_port, ZN => n4745);
   U1869 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_7_port, B1 => 
                           n4894, B2 => REGISTERS_6_7_port, ZN => n4744);
   U1870 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_7_port, B1 => 
                           n4933, B2 => REGISTERS_2_7_port, ZN => n4743);
   U1871 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_7_port, B1 => 
                           n4931, B2 => REGISTERS_1_7_port, ZN => n4742);
   U1872 : NAND4_X1 port map( A1 => n4745, A2 => n4744, A3 => n4743, A4 => 
                           n4742, ZN => n4751);
   U1873 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_7_port, B1 => 
                           n4945, B2 => REGISTERS_11_7_port, ZN => n4749);
   U1874 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_7_port, B1 => 
                           n4932, B2 => REGISTERS_15_7_port, ZN => n4748);
   U1875 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_7_port, B1 => 
                           n4933, B2 => REGISTERS_10_7_port, ZN => n4747);
   U1876 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_7_port, B1 => 
                           n4894, B2 => REGISTERS_14_7_port, ZN => n4746);
   U1877 : NAND4_X1 port map( A1 => n4749, A2 => n4748, A3 => n4747, A4 => 
                           n4746, ZN => n4750);
   U1878 : AOI22_X1 port map( A1 => n4955, A2 => n4751, B1 => n4953, B2 => 
                           n4750, ZN => n4752);
   U1879 : OAI21_X1 port map( B1 => n4958, B2 => n4753, A => n4752, ZN => N424)
                           ;
   U1880 : AOI22_X1 port map( A1 => n4754, A2 => REGISTERS_30_6_port, B1 => 
                           n4882, B2 => REGISTERS_18_6_port, ZN => n4758);
   U1881 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_6_port, B1 => 
                           n4849, B2 => REGISTERS_20_6_port, ZN => n4757);
   U1882 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_6_port, B1 => 
                           n4922, B2 => REGISTERS_28_6_port, ZN => n4756);
   U1883 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_6_port, B1 => 
                           n4850, B2 => REGISTERS_19_6_port, ZN => n4755);
   U1884 : NAND4_X1 port map( A1 => n4758, A2 => n4757, A3 => n4756, A4 => 
                           n4755, ZN => n4764);
   U1885 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_6_port, B1 => 
                           n4921, B2 => REGISTERS_31_6_port, ZN => n4762);
   U1886 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_6_port, B1 => 
                           n4825, B2 => REGISTERS_25_6_port, ZN => n4761);
   U1887 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_6_port, B1 => 
                           n4908, B2 => REGISTERS_29_6_port, ZN => n4760);
   U1888 : AOI22_X1 port map( A1 => n4848, A2 => REGISTERS_23_6_port, B1 => 
                           n4915, B2 => REGISTERS_27_6_port, ZN => n4759);
   U1889 : NAND4_X1 port map( A1 => n4762, A2 => n4761, A3 => n4760, A4 => 
                           n4759, ZN => n4763);
   U1890 : NOR2_X1 port map( A1 => n4764, A2 => n4763, ZN => n4776);
   U1891 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_6_port, B1 => 
                           n4933, B2 => REGISTERS_2_6_port, ZN => n4768);
   U1892 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_6_port, B1 => 
                           n4940, B2 => REGISTERS_5_6_port, ZN => n4767);
   U1893 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_6_6_port, B1 => 
                           n4945, B2 => REGISTERS_3_6_port, ZN => n4766);
   U1894 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_1_6_port, B1 => 
                           n4932, B2 => REGISTERS_7_6_port, ZN => n4765);
   U1895 : NAND4_X1 port map( A1 => n4768, A2 => n4767, A3 => n4766, A4 => 
                           n4765, ZN => n4774);
   U1896 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_6_port, B1 => 
                           n4934, B2 => REGISTERS_11_6_port, ZN => n4772);
   U1897 : AOI22_X1 port map( A1 => n4931, A2 => REGISTERS_9_6_port, B1 => 
                           n4933, B2 => REGISTERS_10_6_port, ZN => n4771);
   U1898 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_6_port, B1 => 
                           n4932, B2 => REGISTERS_15_6_port, ZN => n4770);
   U1899 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_6_port, B1 => 
                           n4894, B2 => REGISTERS_14_6_port, ZN => n4769);
   U1900 : NAND4_X1 port map( A1 => n4772, A2 => n4771, A3 => n4770, A4 => 
                           n4769, ZN => n4773);
   U1901 : AOI22_X1 port map( A1 => n4955, A2 => n4774, B1 => n4953, B2 => 
                           n4773, ZN => n4775);
   U1902 : OAI21_X1 port map( B1 => n4958, B2 => n4776, A => n4775, ZN => N423)
                           ;
   U1903 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_5_port, B1 => 
                           n4918, B2 => REGISTERS_26_5_port, ZN => n4780);
   U1904 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_5_port, B1 => 
                           n4848, B2 => REGISTERS_23_5_port, ZN => n4779);
   U1905 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_5_port, B1 => 
                           n4910, B2 => REGISTERS_22_5_port, ZN => n4778);
   U1906 : AOI22_X1 port map( A1 => n4850, A2 => REGISTERS_19_5_port, B1 => 
                           n4921, B2 => REGISTERS_31_5_port, ZN => n4777);
   U1907 : NAND4_X1 port map( A1 => n4780, A2 => n4779, A3 => n4778, A4 => 
                           n4777, ZN => n4786);
   U1908 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_5_port, B1 => 
                           n4825, B2 => REGISTERS_25_5_port, ZN => n4784);
   U1909 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_5_port, B1 => 
                           n4915, B2 => REGISTERS_27_5_port, ZN => n4783);
   U1910 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_5_port, B1 => 
                           n4919, B2 => REGISTERS_30_5_port, ZN => n4782);
   U1911 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_5_port, B1 => 
                           n4882, B2 => REGISTERS_18_5_port, ZN => n4781);
   U1912 : NAND4_X1 port map( A1 => n4784, A2 => n4783, A3 => n4782, A4 => 
                           n4781, ZN => n4785);
   U1913 : NOR2_X1 port map( A1 => n4786, A2 => n4785, ZN => n4798);
   U1914 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_5_port, B1 => 
                           n4945, B2 => REGISTERS_3_5_port, ZN => n4790);
   U1915 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_5_port, B1 => 
                           n4932, B2 => REGISTERS_7_5_port, ZN => n4789);
   U1916 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_5_port, B1 => 
                           n4894, B2 => REGISTERS_6_5_port, ZN => n4788);
   U1917 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_5_port, B1 => 
                           n4867, B2 => REGISTERS_4_5_port, ZN => n4787);
   U1918 : NAND4_X1 port map( A1 => n4790, A2 => n4789, A3 => n4788, A4 => 
                           n4787, ZN => n4796);
   U1919 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_5_port, B1 => 
                           n4867, B2 => REGISTERS_12_5_port, ZN => n4794);
   U1920 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_5_port, B1 => 
                           n4932, B2 => REGISTERS_15_5_port, ZN => n4793);
   U1921 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_5_port, B1 => 
                           n4933, B2 => REGISTERS_10_5_port, ZN => n4792);
   U1922 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_9_5_port, B1 => 
                           n4934, B2 => REGISTERS_11_5_port, ZN => n4791);
   U1923 : NAND4_X1 port map( A1 => n4794, A2 => n4793, A3 => n4792, A4 => 
                           n4791, ZN => n4795);
   U1924 : AOI22_X1 port map( A1 => n4955, A2 => n4796, B1 => n4953, B2 => 
                           n4795, ZN => n4797);
   U1925 : OAI21_X1 port map( B1 => n4958, B2 => n4798, A => n4797, ZN => N422)
                           ;
   U1926 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_4_port, B1 => 
                           n4850, B2 => REGISTERS_19_4_port, ZN => n4802);
   U1927 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_4_port, B1 => 
                           n4849, B2 => REGISTERS_20_4_port, ZN => n4801);
   U1928 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_4_port, B1 => 
                           n4848, B2 => REGISTERS_23_4_port, ZN => n4800);
   U1929 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_4_port, B1 => 
                           n4882, B2 => REGISTERS_18_4_port, ZN => n4799);
   U1930 : NAND4_X1 port map( A1 => n4802, A2 => n4801, A3 => n4800, A4 => 
                           n4799, ZN => n4810);
   U1931 : AOI22_X1 port map( A1 => n4803, A2 => REGISTERS_26_4_port, B1 => 
                           n4919, B2 => REGISTERS_30_4_port, ZN => n4808);
   U1932 : AOI22_X1 port map( A1 => n4804, A2 => REGISTERS_17_4_port, B1 => 
                           n4825, B2 => REGISTERS_25_4_port, ZN => n4807);
   U1933 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_4_port, B1 => 
                           n4915, B2 => REGISTERS_27_4_port, ZN => n4806);
   U1934 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_4_port, B1 => 
                           n4921, B2 => REGISTERS_31_4_port, ZN => n4805);
   U1935 : NAND4_X1 port map( A1 => n4808, A2 => n4807, A3 => n4806, A4 => 
                           n4805, ZN => n4809);
   U1936 : NOR2_X1 port map( A1 => n4810, A2 => n4809, ZN => n4824);
   U1937 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_4_port, B1 => 
                           n4931, B2 => REGISTERS_1_4_port, ZN => n4814);
   U1938 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_4_port, B1 => 
                           n4932, B2 => REGISTERS_7_4_port, ZN => n4813);
   U1939 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_4_port, B1 => 
                           n4947, B2 => REGISTERS_6_4_port, ZN => n4812);
   U1940 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_4_port, B1 => 
                           n4945, B2 => REGISTERS_3_4_port, ZN => n4811);
   U1941 : NAND4_X1 port map( A1 => n4814, A2 => n4813, A3 => n4812, A4 => 
                           n4811, ZN => n4822);
   U1942 : AOI22_X1 port map( A1 => n4815, A2 => REGISTERS_9_4_port, B1 => 
                           n4934, B2 => REGISTERS_11_4_port, ZN => n4820);
   U1943 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_4_port, B1 => 
                           n4932, B2 => REGISTERS_15_4_port, ZN => n4819);
   U1944 : AOI22_X1 port map( A1 => n4816, A2 => REGISTERS_12_4_port, B1 => 
                           n4894, B2 => REGISTERS_14_4_port, ZN => n4818);
   U1945 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_4_port, B1 => 
                           n4933, B2 => REGISTERS_10_4_port, ZN => n4817);
   U1946 : NAND4_X1 port map( A1 => n4820, A2 => n4819, A3 => n4818, A4 => 
                           n4817, ZN => n4821);
   U1947 : AOI22_X1 port map( A1 => n4955, A2 => n4822, B1 => n4953, B2 => 
                           n4821, ZN => n4823);
   U1948 : OAI21_X1 port map( B1 => n4958, B2 => n4824, A => n4823, ZN => N421)
                           ;
   U1949 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_3_port, B1 => 
                           n4882, B2 => REGISTERS_18_3_port, ZN => n4829);
   U1950 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_3_port, B1 => 
                           n4825, B2 => REGISTERS_25_3_port, ZN => n4828);
   U1951 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_3_port, B1 => 
                           n4919, B2 => REGISTERS_30_3_port, ZN => n4827);
   U1952 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_3_port, B1 => 
                           n4915, B2 => REGISTERS_27_3_port, ZN => n4826);
   U1953 : NAND4_X1 port map( A1 => n4829, A2 => n4828, A3 => n4827, A4 => 
                           n4826, ZN => n4835);
   U1954 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_3_port, B1 => 
                           n4909, B2 => REGISTERS_17_3_port, ZN => n4833);
   U1955 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_3_port, B1 => 
                           n4918, B2 => REGISTERS_26_3_port, ZN => n4832);
   U1956 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_3_port, B1 => 
                           n4910, B2 => REGISTERS_22_3_port, ZN => n4831);
   U1957 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_3_port, B1 => 
                           n4905, B2 => REGISTERS_23_3_port, ZN => n4830);
   U1958 : NAND4_X1 port map( A1 => n4833, A2 => n4832, A3 => n4831, A4 => 
                           n4830, ZN => n4834);
   U1959 : NOR2_X1 port map( A1 => n4835, A2 => n4834, ZN => n4847);
   U1960 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_3_port, B1 => 
                           n4934, B2 => REGISTERS_3_3_port, ZN => n4839);
   U1961 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_3_port, B1 => 
                           n4933, B2 => REGISTERS_2_3_port, ZN => n4838);
   U1962 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_3_port, B1 => 
                           n4947, B2 => REGISTERS_6_3_port, ZN => n4837);
   U1963 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_3_port, B1 => 
                           n4932, B2 => REGISTERS_7_3_port, ZN => n4836);
   U1964 : NAND4_X1 port map( A1 => n4839, A2 => n4838, A3 => n4837, A4 => 
                           n4836, ZN => n4845);
   U1965 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_3_port, B1 => 
                           n4940, B2 => REGISTERS_13_3_port, ZN => n4843);
   U1966 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_3_port, B1 => 
                           n4932, B2 => REGISTERS_15_3_port, ZN => n4842);
   U1967 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_3_port, B1 => 
                           n4933, B2 => REGISTERS_10_3_port, ZN => n4841);
   U1968 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_3_port, B1 => 
                           n4934, B2 => REGISTERS_11_3_port, ZN => n4840);
   U1969 : NAND4_X1 port map( A1 => n4843, A2 => n4842, A3 => n4841, A4 => 
                           n4840, ZN => n4844);
   U1970 : AOI22_X1 port map( A1 => n4955, A2 => n4845, B1 => n4953, B2 => 
                           n4844, ZN => n4846);
   U1971 : OAI21_X1 port map( B1 => n4958, B2 => n4847, A => n4846, ZN => N420)
                           ;
   U1972 : AOI22_X1 port map( A1 => n4909, A2 => REGISTERS_17_2_port, B1 => 
                           n4919, B2 => REGISTERS_30_2_port, ZN => n4854);
   U1973 : AOI22_X1 port map( A1 => n4848, A2 => REGISTERS_23_2_port, B1 => 
                           n4882, B2 => REGISTERS_18_2_port, ZN => n4853);
   U1974 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_2_port, B1 => 
                           n4849, B2 => REGISTERS_20_2_port, ZN => n4852);
   U1975 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_2_port, B1 => 
                           n4850, B2 => REGISTERS_19_2_port, ZN => n4851);
   U1976 : NAND4_X1 port map( A1 => n4854, A2 => n4853, A3 => n4852, A4 => 
                           n4851, ZN => n4862);
   U1977 : AOI22_X1 port map( A1 => n4855, A2 => REGISTERS_29_2_port, B1 => 
                           n4916, B2 => REGISTERS_21_2_port, ZN => n4860);
   U1978 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_2_port, B1 => 
                           n4907, B2 => REGISTERS_25_2_port, ZN => n4859);
   U1979 : AOI22_X1 port map( A1 => n4856, A2 => REGISTERS_16_2_port, B1 => 
                           n4915, B2 => REGISTERS_27_2_port, ZN => n4858);
   U1980 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_2_port, B1 => 
                           n4921, B2 => REGISTERS_31_2_port, ZN => n4857);
   U1981 : NAND4_X1 port map( A1 => n4860, A2 => n4859, A3 => n4858, A4 => 
                           n4857, ZN => n4861);
   U1982 : NOR2_X1 port map( A1 => n4862, A2 => n4861, ZN => n4875);
   U1983 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_2_port, B1 => 
                           n4932, B2 => REGISTERS_7_2_port, ZN => n4866);
   U1984 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_2_port, B1 => 
                           n4934, B2 => REGISTERS_3_2_port, ZN => n4865);
   U1985 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_2_port, B1 => 
                           n4867, B2 => REGISTERS_4_2_port, ZN => n4864);
   U1986 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_6_2_port, B1 => 
                           n4942, B2 => REGISTERS_1_2_port, ZN => n4863);
   U1987 : NAND4_X1 port map( A1 => n4866, A2 => n4865, A3 => n4864, A4 => 
                           n4863, ZN => n4873);
   U1988 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_9_2_port, B1 => 
                           n4933, B2 => REGISTERS_10_2_port, ZN => n4871);
   U1989 : AOI22_X1 port map( A1 => n4929, A2 => REGISTERS_14_2_port, B1 => 
                           n4932, B2 => REGISTERS_15_2_port, ZN => n4870);
   U1990 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_8_2_port, B1 => 
                           n4934, B2 => REGISTERS_11_2_port, ZN => n4869);
   U1991 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_2_port, B1 => 
                           n4867, B2 => REGISTERS_12_2_port, ZN => n4868);
   U1992 : NAND4_X1 port map( A1 => n4871, A2 => n4870, A3 => n4869, A4 => 
                           n4868, ZN => n4872);
   U1993 : AOI22_X1 port map( A1 => n4955, A2 => n4873, B1 => n4953, B2 => 
                           n4872, ZN => n4874);
   U1994 : OAI21_X1 port map( B1 => n4958, B2 => n4875, A => n4874, ZN => N419)
                           ;
   U1995 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_1_port, B1 => 
                           n4909, B2 => REGISTERS_17_1_port, ZN => n4880);
   U1996 : AOI22_X1 port map( A1 => n4876, A2 => REGISTERS_22_1_port, B1 => 
                           n4918, B2 => REGISTERS_26_1_port, ZN => n4879);
   U1997 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_1_port, B1 => 
                           n4903, B2 => REGISTERS_16_1_port, ZN => n4878);
   U1998 : AOI22_X1 port map( A1 => n4921, A2 => REGISTERS_31_1_port, B1 => 
                           n4905, B2 => REGISTERS_23_1_port, ZN => n4877);
   U1999 : NAND4_X1 port map( A1 => n4880, A2 => n4879, A3 => n4878, A4 => 
                           n4877, ZN => n4889);
   U2000 : AOI22_X1 port map( A1 => n4907, A2 => REGISTERS_25_1_port, B1 => 
                           n4915, B2 => REGISTERS_27_1_port, ZN => n4887);
   U2001 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_1_port, B1 => 
                           n4919, B2 => REGISTERS_30_1_port, ZN => n4886);
   U2002 : AOI22_X1 port map( A1 => n4881, A2 => REGISTERS_28_1_port, B1 => 
                           n4906, B2 => REGISTERS_20_1_port, ZN => n4885);
   U2003 : AOI22_X1 port map( A1 => n4883, A2 => REGISTERS_21_1_port, B1 => 
                           n4882, B2 => REGISTERS_18_1_port, ZN => n4884);
   U2004 : NAND4_X1 port map( A1 => n4887, A2 => n4886, A3 => n4885, A4 => 
                           n4884, ZN => n4888);
   U2005 : NOR2_X1 port map( A1 => n4889, A2 => n4888, ZN => n4902);
   U2006 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_1_port, B1 => 
                           n4944, B2 => REGISTERS_7_1_port, ZN => n4893);
   U2007 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_1_port, B1 => 
                           n4943, B2 => REGISTERS_4_1_port, ZN => n4892);
   U2008 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_6_1_port, B1 => 
                           n4934, B2 => REGISTERS_3_1_port, ZN => n4891);
   U2009 : AOI22_X1 port map( A1 => n4942, A2 => REGISTERS_1_1_port, B1 => 
                           n4933, B2 => REGISTERS_2_1_port, ZN => n4890);
   U2010 : NAND4_X1 port map( A1 => n4893, A2 => n4892, A3 => n4891, A4 => 
                           n4890, ZN => n4900);
   U2011 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_13_1_port, B1 => 
                           n4931, B2 => REGISTERS_9_1_port, ZN => n4898);
   U2012 : AOI22_X1 port map( A1 => n4946, A2 => REGISTERS_10_1_port, B1 => 
                           n4932, B2 => REGISTERS_15_1_port, ZN => n4897);
   U2013 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_1_port, B1 => 
                           n4894, B2 => REGISTERS_14_1_port, ZN => n4896);
   U2014 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_1_port, B1 => 
                           n4945, B2 => REGISTERS_11_1_port, ZN => n4895);
   U2015 : NAND4_X1 port map( A1 => n4898, A2 => n4897, A3 => n4896, A4 => 
                           n4895, ZN => n4899);
   U2016 : AOI22_X1 port map( A1 => n4955, A2 => n4900, B1 => n4953, B2 => 
                           n4899, ZN => n4901);
   U2017 : OAI21_X1 port map( B1 => n4958, B2 => n4902, A => n4901, ZN => N418)
                           ;
   U2018 : AOI22_X1 port map( A1 => n4904, A2 => REGISTERS_24_0_port, B1 => 
                           n4903, B2 => REGISTERS_16_0_port, ZN => n4914);
   U2019 : AOI22_X1 port map( A1 => n4906, A2 => REGISTERS_20_0_port, B1 => 
                           n4905, B2 => REGISTERS_23_0_port, ZN => n4913);
   U2020 : AOI22_X1 port map( A1 => n4908, A2 => REGISTERS_29_0_port, B1 => 
                           n4907, B2 => REGISTERS_25_0_port, ZN => n4912);
   U2021 : AOI22_X1 port map( A1 => n4910, A2 => REGISTERS_22_0_port, B1 => 
                           n4909, B2 => REGISTERS_17_0_port, ZN => n4911);
   U2022 : NAND4_X1 port map( A1 => n4914, A2 => n4913, A3 => n4912, A4 => 
                           n4911, ZN => n4928);
   U2023 : AOI22_X1 port map( A1 => n4916, A2 => REGISTERS_21_0_port, B1 => 
                           n4915, B2 => REGISTERS_27_0_port, ZN => n4926);
   U2024 : AOI22_X1 port map( A1 => n4918, A2 => REGISTERS_26_0_port, B1 => 
                           n4917, B2 => REGISTERS_18_0_port, ZN => n4925);
   U2025 : AOI22_X1 port map( A1 => n4920, A2 => REGISTERS_19_0_port, B1 => 
                           n4919, B2 => REGISTERS_30_0_port, ZN => n4924);
   U2026 : AOI22_X1 port map( A1 => n4922, A2 => REGISTERS_28_0_port, B1 => 
                           n4921, B2 => REGISTERS_31_0_port, ZN => n4923);
   U2027 : NAND4_X1 port map( A1 => n4926, A2 => n4925, A3 => n4924, A4 => 
                           n4923, ZN => n4927);
   U2028 : NOR2_X1 port map( A1 => n4928, A2 => n4927, ZN => n4957);
   U2029 : AOI22_X1 port map( A1 => n4930, A2 => REGISTERS_5_0_port, B1 => 
                           n4929, B2 => REGISTERS_6_0_port, ZN => n4939);
   U2030 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_4_0_port, B1 => 
                           n4931, B2 => REGISTERS_1_0_port, ZN => n4938);
   U2031 : AOI22_X1 port map( A1 => n4933, A2 => REGISTERS_2_0_port, B1 => 
                           n4932, B2 => REGISTERS_7_0_port, ZN => n4937);
   U2032 : AOI22_X1 port map( A1 => n4935, A2 => REGISTERS_0_0_port, B1 => 
                           n4934, B2 => REGISTERS_3_0_port, ZN => n4936);
   U2033 : NAND4_X1 port map( A1 => n4939, A2 => n4938, A3 => n4937, A4 => 
                           n4936, ZN => n4954);
   U2034 : AOI22_X1 port map( A1 => n4941, A2 => REGISTERS_8_0_port, B1 => 
                           n4940, B2 => REGISTERS_13_0_port, ZN => n4951);
   U2035 : AOI22_X1 port map( A1 => n4943, A2 => REGISTERS_12_0_port, B1 => 
                           n4942, B2 => REGISTERS_9_0_port, ZN => n4950);
   U2036 : AOI22_X1 port map( A1 => n4945, A2 => REGISTERS_11_0_port, B1 => 
                           n4944, B2 => REGISTERS_15_0_port, ZN => n4949);
   U2037 : AOI22_X1 port map( A1 => n4947, A2 => REGISTERS_14_0_port, B1 => 
                           n4946, B2 => REGISTERS_10_0_port, ZN => n4948);
   U2038 : NAND4_X1 port map( A1 => n4951, A2 => n4950, A3 => n4949, A4 => 
                           n4948, ZN => n4952);
   U2039 : AOI22_X1 port map( A1 => n4955, A2 => n4954, B1 => n4953, B2 => 
                           n4952, ZN => n4956);
   U2040 : OAI21_X1 port map( B1 => n4958, B2 => n4957, A => n4956, ZN => N417)
                           ;
   U2041 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n4967);
   U2042 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), ZN => n4959);
   U2043 : INV_X1 port map( A => ADD_RD1(1), ZN => n4965);
   U2044 : NAND2_X1 port map( A1 => n4959, A2 => n4965, ZN => n4975);
   U2045 : NOR2_X1 port map( A1 => n4967, A2 => n4975, ZN => n5699);
   U2046 : INV_X1 port map( A => ADD_RD1(3), ZN => n4984);
   U2047 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n4984, ZN => n4966);
   U2048 : INV_X1 port map( A => ADD_RD1(2), ZN => n4964);
   U2049 : OR3_X1 port map( A1 => n4964, A2 => ADD_RD1(1), A3 => ADD_RD1(0), ZN
                           => n5047);
   U2050 : NOR2_X1 port map( A1 => n4966, A2 => n5047, ZN => n5599);
   U2051 : CLKBUF_X1 port map( A => n5599, Z => n5683);
   U2052 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n5699, B1 => 
                           REGISTERS_20_31_port, B2 => n5683, ZN => n4963);
   U2053 : NOR2_X1 port map( A1 => n4966, A2 => n4975, ZN => n5700);
   U2054 : NAND2_X1 port map( A1 => ADD_RD1(1), A2 => n4959, ZN => n4977);
   U2055 : NOR2_X1 port map( A1 => n4967, A2 => n4977, ZN => n5688);
   U2056 : CLKBUF_X1 port map( A => n5688, Z => n5657);
   U2057 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n5700, B1 => 
                           REGISTERS_26_31_port, B2 => n5657, ZN => n4962);
   U2058 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n4965, 
                           ZN => n4978);
   U2059 : NOR2_X1 port map( A1 => n4966, A2 => n4978, ZN => n5654);
   U2060 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => 
                           ADD_RD1(2), ZN => n4979);
   U2061 : NOR2_X1 port map( A1 => n4966, A2 => n4979, ZN => n5697);
   U2062 : CLKBUF_X1 port map( A => n5697, Z => n5656);
   U2063 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n5654, B1 => 
                           REGISTERS_23_31_port, B2 => n5656, ZN => n4961);
   U2064 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n4964, 
                           ZN => n4976);
   U2065 : NOR2_X1 port map( A1 => n4966, A2 => n4976, ZN => n5686);
   U2066 : NOR2_X1 port map( A1 => n4966, A2 => n4977, ZN => n5645);
   U2067 : CLKBUF_X1 port map( A => n5645, Z => n5684);
   U2068 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n5686, B1 => 
                           REGISTERS_18_31_port, B2 => n5684, ZN => n4960);
   U2069 : NAND4_X1 port map( A1 => n4963, A2 => n4962, A3 => n4961, A4 => 
                           n4960, ZN => n4973);
   U2070 : NOR2_X1 port map( A1 => n4967, A2 => n5047, ZN => n5648);
   U2071 : NOR2_X1 port map( A1 => n4967, A2 => n4979, ZN => n5624);
   U2072 : CLKBUF_X1 port map( A => n5624, Z => n5698);
   U2073 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n5648, B1 => 
                           REGISTERS_31_31_port, B2 => n5698, ZN => n4971);
   U2074 : OR3_X1 port map( A1 => n4965, A2 => n4964, A3 => ADD_RD1(0), ZN => 
                           n5070);
   U2075 : NOR2_X1 port map( A1 => n5070, A2 => n4966, ZN => n5594);
   U2076 : NOR2_X1 port map( A1 => n5070, A2 => n4967, ZN => n5696);
   U2077 : CLKBUF_X1 port map( A => n5696, Z => n5619);
   U2078 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n5594, B1 => 
                           REGISTERS_30_31_port, B2 => n5619, ZN => n4970);
   U2079 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n4965, A3 => n4964, ZN =>
                           n4974);
   U2080 : NOR2_X1 port map( A1 => n4966, A2 => n4974, ZN => n5570);
   U2081 : NOR2_X1 port map( A1 => n4967, A2 => n4976, ZN => n5694);
   U2082 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n5570, B1 => 
                           REGISTERS_27_31_port, B2 => n5694, ZN => n4969);
   U2083 : NOR2_X1 port map( A1 => n4967, A2 => n4978, ZN => n5655);
   U2084 : NOR2_X1 port map( A1 => n4967, A2 => n4974, ZN => n5625);
   U2085 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n5655, B1 => 
                           REGISTERS_25_31_port, B2 => n5625, ZN => n4968);
   U2086 : NAND4_X1 port map( A1 => n4971, A2 => n4970, A3 => n4969, A4 => 
                           n4968, ZN => n4972);
   U2087 : NOR2_X1 port map( A1 => n4973, A2 => n4972, ZN => n4992);
   U2088 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n5732, 
                           ZN => n5302);
   U2089 : CLKBUF_X1 port map( A => n5302, Z => n5501);
   U2090 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n5708, B1 => 
                           REGISTERS_0_31_port, B2 => n5720, ZN => n4983);
   U2091 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n5717, B1 => 
                           REGISTERS_2_31_port, B2 => n5707, ZN => n4982);
   U2092 : INV_X1 port map( A => n5047, ZN => n5721);
   U2093 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n5721, B1 => 
                           REGISTERS_5_31_port, B2 => n5718, ZN => n4981);
   U2094 : INV_X1 port map( A => n5070, ZN => n5716);
   U2095 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n5671, B1 => 
                           REGISTERS_6_31_port, B2 => n5716, ZN => n4980);
   U2096 : NAND4_X1 port map( A1 => n4983, A2 => n4982, A3 => n4981, A4 => 
                           n4980, ZN => n4990);
   U2097 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n4984, A3 => n5732, ZN => 
                           n5212);
   U2098 : CLKBUF_X1 port map( A => n5212, Z => n5727);
   U2099 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n5718, B1 => 
                           REGISTERS_10_31_port, B2 => n5707, ZN => n4988);
   U2100 : CLKBUF_X1 port map( A => n5720, Z => n5668);
   U2101 : INV_X1 port map( A => n5070, ZN => n5670);
   U2102 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n5668, B1 => 
                           REGISTERS_14_31_port, B2 => n5670, ZN => n4987);
   U2103 : INV_X1 port map( A => n5047, ZN => n5610);
   U2104 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n5610, B1 => 
                           REGISTERS_9_31_port, B2 => n5708, ZN => n4986);
   U2105 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n5671, B1 => 
                           REGISTERS_11_31_port, B2 => n5717, ZN => n4985);
   U2106 : NAND4_X1 port map( A1 => n4988, A2 => n4987, A3 => n4986, A4 => 
                           n4985, ZN => n4989);
   U2107 : AOI22_X1 port map( A1 => n5501, A2 => n4990, B1 => n5727, B2 => 
                           n4989, ZN => n4991);
   U2108 : OAI21_X1 port map( B1 => n5732, B2 => n4992, A => n4991, ZN => N416)
                           ;
   U2109 : CLKBUF_X1 port map( A => n5625, Z => n5693);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n5693, B1 => 
                           REGISTERS_31_30_port, B2 => n5698, ZN => n4996);
   U2111 : CLKBUF_X1 port map( A => n5655, Z => n5685);
   U2112 : CLKBUF_X1 port map( A => n5686, Z => n5626);
   U2113 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n5685, B1 => 
                           REGISTERS_19_30_port, B2 => n5626, ZN => n4995);
   U2114 : CLKBUF_X1 port map( A => n5694, Z => n5646);
   U2115 : CLKBUF_X1 port map( A => n5654, Z => n5687);
   U2116 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n5646, B1 => 
                           REGISTERS_21_30_port, B2 => n5687, ZN => n4994);
   U2117 : CLKBUF_X1 port map( A => n5594, Z => n5681);
   U2118 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n5699, B1 => 
                           REGISTERS_22_30_port, B2 => n5681, ZN => n4993);
   U2119 : NAND4_X1 port map( A1 => n4996, A2 => n4995, A3 => n4994, A4 => 
                           n4993, ZN => n5002);
   U2120 : CLKBUF_X1 port map( A => n5648, Z => n5682);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n5570, B1 => 
                           REGISTERS_28_30_port, B2 => n5682, ZN => n5000);
   U2122 : CLKBUF_X1 port map( A => n5700, Z => n5647);
   U2123 : AOI22_X1 port map( A1 => REGISTERS_26_30_port, A2 => n5688, B1 => 
                           REGISTERS_16_30_port, B2 => n5647, ZN => n4999);
   U2124 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n5656, B1 => 
                           REGISTERS_20_30_port, B2 => n5683, ZN => n4998);
   U2125 : AOI22_X1 port map( A1 => REGISTERS_18_30_port, A2 => n5684, B1 => 
                           REGISTERS_30_30_port, B2 => n5696, ZN => n4997);
   U2126 : NAND4_X1 port map( A1 => n5000, A2 => n4999, A3 => n4998, A4 => 
                           n4997, ZN => n5001);
   U2127 : NOR2_X1 port map( A1 => n5002, A2 => n5001, ZN => n5014);
   U2128 : AOI22_X1 port map( A1 => REGISTERS_6_30_port, A2 => n5716, B1 => 
                           REGISTERS_7_30_port, B2 => n5671, ZN => n5006);
   U2129 : CLKBUF_X1 port map( A => n5717, Z => n5710);
   U2130 : AOI22_X1 port map( A1 => REGISTERS_2_30_port, A2 => n5707, B1 => 
                           REGISTERS_3_30_port, B2 => n5710, ZN => n5005);
   U2131 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n5708, B1 => 
                           REGISTERS_4_30_port, B2 => n5721, ZN => n5004);
   U2132 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n5718, B1 => 
                           REGISTERS_0_30_port, B2 => n5668, ZN => n5003);
   U2133 : NAND4_X1 port map( A1 => n5006, A2 => n5005, A3 => n5004, A4 => 
                           n5003, ZN => n5012);
   U2134 : AOI22_X1 port map( A1 => REGISTERS_14_30_port, A2 => n5716, B1 => 
                           REGISTERS_13_30_port, B2 => n5718, ZN => n5010);
   U2135 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n5708, B1 => 
                           REGISTERS_12_30_port, B2 => n5721, ZN => n5009);
   U2136 : CLKBUF_X1 port map( A => n5671, Z => n5711);
   U2137 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n5720, B1 => 
                           REGISTERS_15_30_port, B2 => n5711, ZN => n5008);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_10_30_port, A2 => n5707, B1 => 
                           REGISTERS_11_30_port, B2 => n5710, ZN => n5007);
   U2139 : NAND4_X1 port map( A1 => n5010, A2 => n5009, A3 => n5008, A4 => 
                           n5007, ZN => n5011);
   U2140 : AOI22_X1 port map( A1 => n5501, A2 => n5012, B1 => n5727, B2 => 
                           n5011, ZN => n5013);
   U2141 : OAI21_X1 port map( B1 => n5732, B2 => n5014, A => n5013, ZN => N415)
                           ;
   U2142 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n5682, B1 => 
                           REGISTERS_21_29_port, B2 => n5687, ZN => n5018);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n5685, B1 => 
                           REGISTERS_25_29_port, B2 => n5693, ZN => n5017);
   U2144 : CLKBUF_X1 port map( A => n5570, Z => n5695);
   U2145 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n5626, B1 => 
                           REGISTERS_17_29_port, B2 => n5695, ZN => n5016);
   U2146 : AOI22_X1 port map( A1 => REGISTERS_18_29_port, A2 => n5684, B1 => 
                           REGISTERS_20_29_port, B2 => n5683, ZN => n5015);
   U2147 : NAND4_X1 port map( A1 => n5018, A2 => n5017, A3 => n5016, A4 => 
                           n5015, ZN => n5024);
   U2148 : AOI22_X1 port map( A1 => REGISTERS_22_29_port, A2 => n5681, B1 => 
                           REGISTERS_26_29_port, B2 => n5657, ZN => n5022);
   U2149 : CLKBUF_X1 port map( A => n5699, Z => n5653);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n5694, B1 => 
                           REGISTERS_24_29_port, B2 => n5653, ZN => n5021);
   U2151 : AOI22_X1 port map( A1 => REGISTERS_31_29_port, A2 => n5698, B1 => 
                           REGISTERS_30_29_port, B2 => n5619, ZN => n5020);
   U2152 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n5697, B1 => 
                           REGISTERS_16_29_port, B2 => n5647, ZN => n5019);
   U2153 : NAND4_X1 port map( A1 => n5022, A2 => n5021, A3 => n5020, A4 => 
                           n5019, ZN => n5023);
   U2154 : NOR2_X1 port map( A1 => n5024, A2 => n5023, ZN => n5036);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_2_29_port, A2 => n5707, B1 => 
                           REGISTERS_7_29_port, B2 => n5671, ZN => n5028);
   U2156 : CLKBUF_X1 port map( A => n5718, Z => n5581);
   U2157 : AOI22_X1 port map( A1 => REGISTERS_6_29_port, A2 => n5670, B1 => 
                           REGISTERS_5_29_port, B2 => n5581, ZN => n5027);
   U2158 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n5717, B1 => 
                           REGISTERS_4_29_port, B2 => n5721, ZN => n5026);
   U2159 : CLKBUF_X1 port map( A => n5708, Z => n5719);
   U2160 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n5720, B1 => 
                           REGISTERS_1_29_port, B2 => n5719, ZN => n5025);
   U2161 : NAND4_X1 port map( A1 => n5028, A2 => n5027, A3 => n5026, A4 => 
                           n5025, ZN => n5034);
   U2162 : CLKBUF_X1 port map( A => n5707, Z => n5672);
   U2163 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n5717, B1 => 
                           REGISTERS_10_29_port, B2 => n5672, ZN => n5032);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n5610, B1 => 
                           REGISTERS_8_29_port, B2 => n5720, ZN => n5031);
   U2165 : AOI22_X1 port map( A1 => REGISTERS_14_29_port, A2 => n5716, B1 => 
                           REGISTERS_9_29_port, B2 => n5719, ZN => n5030);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n5711, B1 => 
                           REGISTERS_13_29_port, B2 => n5718, ZN => n5029);
   U2167 : NAND4_X1 port map( A1 => n5032, A2 => n5031, A3 => n5030, A4 => 
                           n5029, ZN => n5033);
   U2168 : AOI22_X1 port map( A1 => n5501, A2 => n5034, B1 => n5727, B2 => 
                           n5033, ZN => n5035);
   U2169 : OAI21_X1 port map( B1 => n5732, B2 => n5036, A => n5035, ZN => N414)
                           ;
   U2170 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n5570, B1 => 
                           REGISTERS_25_28_port, B2 => n5693, ZN => n5040);
   U2171 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n5647, B1 => 
                           REGISTERS_28_28_port, B2 => n5682, ZN => n5039);
   U2172 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n5694, B1 => 
                           REGISTERS_21_28_port, B2 => n5687, ZN => n5038);
   U2173 : AOI22_X1 port map( A1 => REGISTERS_18_28_port, A2 => n5684, B1 => 
                           REGISTERS_19_28_port, B2 => n5626, ZN => n5037);
   U2174 : NAND4_X1 port map( A1 => n5040, A2 => n5039, A3 => n5038, A4 => 
                           n5037, ZN => n5046);
   U2175 : AOI22_X1 port map( A1 => REGISTERS_30_28_port, A2 => n5696, B1 => 
                           REGISTERS_31_28_port, B2 => n5698, ZN => n5044);
   U2176 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n5699, B1 => 
                           REGISTERS_26_28_port, B2 => n5657, ZN => n5043);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n5599, B1 => 
                           REGISTERS_29_28_port, B2 => n5685, ZN => n5042);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_23_28_port, A2 => n5697, B1 => 
                           REGISTERS_22_28_port, B2 => n5681, ZN => n5041);
   U2179 : NAND4_X1 port map( A1 => n5044, A2 => n5043, A3 => n5042, A4 => 
                           n5041, ZN => n5045);
   U2180 : NOR2_X1 port map( A1 => n5046, A2 => n5045, ZN => n5059);
   U2181 : INV_X1 port map( A => n5047, ZN => n5669);
   U2182 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n5669, B1 => 
                           REGISTERS_0_28_port, B2 => n5720, ZN => n5051);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n5718, B1 => 
                           REGISTERS_2_28_port, B2 => n5707, ZN => n5050);
   U2184 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n5717, B1 => 
                           REGISTERS_1_28_port, B2 => n5719, ZN => n5049);
   U2185 : AOI22_X1 port map( A1 => REGISTERS_6_28_port, A2 => n5716, B1 => 
                           REGISTERS_7_28_port, B2 => n5671, ZN => n5048);
   U2186 : NAND4_X1 port map( A1 => n5051, A2 => n5050, A3 => n5049, A4 => 
                           n5048, ZN => n5057);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n5718, B1 => 
                           REGISTERS_14_28_port, B2 => n5716, ZN => n5055);
   U2188 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n5717, B1 => 
                           REGISTERS_10_28_port, B2 => n5707, ZN => n5054);
   U2189 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n5671, B1 => 
                           REGISTERS_8_28_port, B2 => n5668, ZN => n5053);
   U2190 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n5708, B1 => 
                           REGISTERS_12_28_port, B2 => n5610, ZN => n5052);
   U2191 : NAND4_X1 port map( A1 => n5055, A2 => n5054, A3 => n5053, A4 => 
                           n5052, ZN => n5056);
   U2192 : AOI22_X1 port map( A1 => n5501, A2 => n5057, B1 => n5727, B2 => 
                           n5056, ZN => n5058);
   U2193 : OAI21_X1 port map( B1 => n5732, B2 => n5059, A => n5058, ZN => N413)
                           ;
   U2194 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n5699, B1 => 
                           REGISTERS_19_27_port, B2 => n5626, ZN => n5063);
   U2195 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n5687, B1 => 
                           REGISTERS_17_27_port, B2 => n5695, ZN => n5062);
   U2196 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n5693, B1 => 
                           REGISTERS_20_27_port, B2 => n5683, ZN => n5061);
   U2197 : AOI22_X1 port map( A1 => REGISTERS_18_27_port, A2 => n5684, B1 => 
                           REGISTERS_16_27_port, B2 => n5647, ZN => n5060);
   U2198 : NAND4_X1 port map( A1 => n5063, A2 => n5062, A3 => n5061, A4 => 
                           n5060, ZN => n5069);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n5697, B1 => 
                           REGISTERS_30_27_port, B2 => n5619, ZN => n5067);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n5698, B1 => 
                           REGISTERS_28_27_port, B2 => n5682, ZN => n5066);
   U2201 : AOI22_X1 port map( A1 => REGISTERS_22_27_port, A2 => n5681, B1 => 
                           REGISTERS_29_27_port, B2 => n5655, ZN => n5065);
   U2202 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n5694, B1 => 
                           REGISTERS_26_27_port, B2 => n5657, ZN => n5064);
   U2203 : NAND4_X1 port map( A1 => n5067, A2 => n5066, A3 => n5065, A4 => 
                           n5064, ZN => n5068);
   U2204 : NOR2_X1 port map( A1 => n5069, A2 => n5068, ZN => n5082);
   U2205 : INV_X1 port map( A => n5070, ZN => n5709);
   U2206 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n5708, B1 => 
                           REGISTERS_6_27_port, B2 => n5709, ZN => n5074);
   U2207 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n5671, B1 => 
                           REGISTERS_3_27_port, B2 => n5710, ZN => n5073);
   U2208 : AOI22_X1 port map( A1 => REGISTERS_2_27_port, A2 => n5707, B1 => 
                           REGISTERS_5_27_port, B2 => n5581, ZN => n5072);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n5720, B1 => 
                           REGISTERS_4_27_port, B2 => n5610, ZN => n5071);
   U2210 : NAND4_X1 port map( A1 => n5074, A2 => n5073, A3 => n5072, A4 => 
                           n5071, ZN => n5080);
   U2211 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n5717, B1 => 
                           REGISTERS_15_27_port, B2 => n5671, ZN => n5078);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n5720, B1 => 
                           REGISTERS_12_27_port, B2 => n5669, ZN => n5077);
   U2213 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n5719, B1 => 
                           REGISTERS_13_27_port, B2 => n5581, ZN => n5076);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_14_27_port, A2 => n5716, B1 => 
                           REGISTERS_10_27_port, B2 => n5707, ZN => n5075);
   U2215 : NAND4_X1 port map( A1 => n5078, A2 => n5077, A3 => n5076, A4 => 
                           n5075, ZN => n5079);
   U2216 : AOI22_X1 port map( A1 => n5501, A2 => n5080, B1 => n5212, B2 => 
                           n5079, ZN => n5081);
   U2217 : OAI21_X1 port map( B1 => n5732, B2 => n5082, A => n5081, ZN => N412)
                           ;
   U2218 : AOI22_X1 port map( A1 => REGISTERS_31_26_port, A2 => n5698, B1 => 
                           REGISTERS_16_26_port, B2 => n5647, ZN => n5086);
   U2219 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n5694, B1 => 
                           REGISTERS_21_26_port, B2 => n5687, ZN => n5085);
   U2220 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n5699, B1 => 
                           REGISTERS_26_26_port, B2 => n5657, ZN => n5084);
   U2221 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n5685, B1 => 
                           REGISTERS_23_26_port, B2 => n5656, ZN => n5083);
   U2222 : NAND4_X1 port map( A1 => n5086, A2 => n5085, A3 => n5084, A4 => 
                           n5083, ZN => n5092);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n5682, B1 => 
                           REGISTERS_18_26_port, B2 => n5684, ZN => n5090);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n5570, B1 => 
                           REGISTERS_20_26_port, B2 => n5683, ZN => n5089);
   U2225 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n5626, B1 => 
                           REGISTERS_25_26_port, B2 => n5693, ZN => n5088);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_30_26_port, A2 => n5696, B1 => 
                           REGISTERS_22_26_port, B2 => n5594, ZN => n5087);
   U2227 : NAND4_X1 port map( A1 => n5090, A2 => n5089, A3 => n5088, A4 => 
                           n5087, ZN => n5091);
   U2228 : NOR2_X1 port map( A1 => n5092, A2 => n5091, ZN => n5104);
   U2229 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n5719, B1 => 
                           REGISTERS_6_26_port, B2 => n5716, ZN => n5096);
   U2230 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n5717, B1 => 
                           REGISTERS_5_26_port, B2 => n5581, ZN => n5095);
   U2231 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n5720, B1 => 
                           REGISTERS_2_26_port, B2 => n5707, ZN => n5094);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n5671, B1 => 
                           REGISTERS_4_26_port, B2 => n5669, ZN => n5093);
   U2233 : NAND4_X1 port map( A1 => n5096, A2 => n5095, A3 => n5094, A4 => 
                           n5093, ZN => n5102);
   U2234 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n5717, B1 => 
                           REGISTERS_10_26_port, B2 => n5707, ZN => n5100);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n5711, B1 => 
                           REGISTERS_9_26_port, B2 => n5719, ZN => n5099);
   U2236 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n5718, B1 => 
                           REGISTERS_8_26_port, B2 => n5720, ZN => n5098);
   U2237 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n5610, B1 => 
                           REGISTERS_14_26_port, B2 => n5709, ZN => n5097);
   U2238 : NAND4_X1 port map( A1 => n5100, A2 => n5099, A3 => n5098, A4 => 
                           n5097, ZN => n5101);
   U2239 : AOI22_X1 port map( A1 => n5501, A2 => n5102, B1 => n5212, B2 => 
                           n5101, ZN => n5103);
   U2240 : OAI21_X1 port map( B1 => n5732, B2 => n5104, A => n5103, ZN => N411)
                           ;
   U2241 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n5682, B1 => 
                           REGISTERS_27_25_port, B2 => n5646, ZN => n5108);
   U2242 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n5687, B1 => 
                           REGISTERS_20_25_port, B2 => n5683, ZN => n5107);
   U2243 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n5626, B1 => 
                           REGISTERS_29_25_port, B2 => n5685, ZN => n5106);
   U2244 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n5698, B1 => 
                           REGISTERS_22_25_port, B2 => n5594, ZN => n5105);
   U2245 : NAND4_X1 port map( A1 => n5108, A2 => n5107, A3 => n5106, A4 => 
                           n5105, ZN => n5114);
   U2246 : AOI22_X1 port map( A1 => REGISTERS_18_25_port, A2 => n5684, B1 => 
                           REGISTERS_23_25_port, B2 => n5656, ZN => n5112);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n5570, B1 => 
                           REGISTERS_25_25_port, B2 => n5693, ZN => n5111);
   U2248 : AOI22_X1 port map( A1 => REGISTERS_30_25_port, A2 => n5696, B1 => 
                           REGISTERS_24_25_port, B2 => n5653, ZN => n5110);
   U2249 : AOI22_X1 port map( A1 => REGISTERS_26_25_port, A2 => n5657, B1 => 
                           REGISTERS_16_25_port, B2 => n5647, ZN => n5109);
   U2250 : NAND4_X1 port map( A1 => n5112, A2 => n5111, A3 => n5110, A4 => 
                           n5109, ZN => n5113);
   U2251 : NOR2_X1 port map( A1 => n5114, A2 => n5113, ZN => n5126);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n5708, B1 => 
                           REGISTERS_4_25_port, B2 => n5669, ZN => n5118);
   U2253 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n5717, B1 => 
                           REGISTERS_5_25_port, B2 => n5581, ZN => n5117);
   U2254 : AOI22_X1 port map( A1 => REGISTERS_2_25_port, A2 => n5707, B1 => 
                           REGISTERS_7_25_port, B2 => n5671, ZN => n5116);
   U2255 : AOI22_X1 port map( A1 => REGISTERS_6_25_port, A2 => n5709, B1 => 
                           REGISTERS_0_25_port, B2 => n5720, ZN => n5115);
   U2256 : NAND4_X1 port map( A1 => n5118, A2 => n5117, A3 => n5116, A4 => 
                           n5115, ZN => n5124);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_14_25_port, A2 => n5670, B1 => 
                           REGISTERS_9_25_port, B2 => n5708, ZN => n5122);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n5671, B1 => 
                           REGISTERS_12_25_port, B2 => n5669, ZN => n5121);
   U2259 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n5710, B1 => 
                           REGISTERS_13_25_port, B2 => n5581, ZN => n5120);
   U2260 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n5720, B1 => 
                           REGISTERS_10_25_port, B2 => n5707, ZN => n5119);
   U2261 : NAND4_X1 port map( A1 => n5122, A2 => n5121, A3 => n5120, A4 => 
                           n5119, ZN => n5123);
   U2262 : AOI22_X1 port map( A1 => n5501, A2 => n5124, B1 => n5212, B2 => 
                           n5123, ZN => n5125);
   U2263 : OAI21_X1 port map( B1 => n5732, B2 => n5126, A => n5125, ZN => N410)
                           ;
   U2264 : AOI22_X1 port map( A1 => REGISTERS_30_24_port, A2 => n5696, B1 => 
                           REGISTERS_19_24_port, B2 => n5626, ZN => n5130);
   U2265 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n5684, B1 => 
                           REGISTERS_23_24_port, B2 => n5656, ZN => n5129);
   U2266 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n5599, B1 => 
                           REGISTERS_28_24_port, B2 => n5682, ZN => n5128);
   U2267 : AOI22_X1 port map( A1 => REGISTERS_22_24_port, A2 => n5681, B1 => 
                           REGISTERS_31_24_port, B2 => n5698, ZN => n5127);
   U2268 : NAND4_X1 port map( A1 => n5130, A2 => n5129, A3 => n5128, A4 => 
                           n5127, ZN => n5136);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n5700, B1 => 
                           REGISTERS_25_24_port, B2 => n5693, ZN => n5134);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n5687, B1 => 
                           REGISTERS_26_24_port, B2 => n5657, ZN => n5133);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n5646, B1 => 
                           REGISTERS_17_24_port, B2 => n5695, ZN => n5132);
   U2272 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n5685, B1 => 
                           REGISTERS_24_24_port, B2 => n5653, ZN => n5131);
   U2273 : NAND4_X1 port map( A1 => n5134, A2 => n5133, A3 => n5132, A4 => 
                           n5131, ZN => n5135);
   U2274 : NOR2_X1 port map( A1 => n5136, A2 => n5135, ZN => n5148);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n5708, B1 => 
                           REGISTERS_6_24_port, B2 => n5709, ZN => n5140);
   U2276 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n5717, B1 => 
                           REGISTERS_5_24_port, B2 => n5581, ZN => n5139);
   U2277 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n5671, B1 => 
                           REGISTERS_2_24_port, B2 => n5672, ZN => n5138);
   U2278 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n5610, B1 => 
                           REGISTERS_0_24_port, B2 => n5668, ZN => n5137);
   U2279 : NAND4_X1 port map( A1 => n5140, A2 => n5139, A3 => n5138, A4 => 
                           n5137, ZN => n5146);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_10_24_port, A2 => n5707, B1 => 
                           REGISTERS_8_24_port, B2 => n5720, ZN => n5144);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n5717, B1 => 
                           REGISTERS_13_24_port, B2 => n5581, ZN => n5143);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n5610, B1 => 
                           REGISTERS_15_24_port, B2 => n5711, ZN => n5142);
   U2283 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n5719, B1 => 
                           REGISTERS_14_24_port, B2 => n5709, ZN => n5141);
   U2284 : NAND4_X1 port map( A1 => n5144, A2 => n5143, A3 => n5142, A4 => 
                           n5141, ZN => n5145);
   U2285 : AOI22_X1 port map( A1 => n5501, A2 => n5146, B1 => n5212, B2 => 
                           n5145, ZN => n5147);
   U2286 : OAI21_X1 port map( B1 => n5732, B2 => n5148, A => n5147, ZN => N409)
                           ;
   U2287 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n5685, B1 => 
                           REGISTERS_31_23_port, B2 => n5698, ZN => n5152);
   U2288 : AOI22_X1 port map( A1 => REGISTERS_22_23_port, A2 => n5681, B1 => 
                           REGISTERS_23_23_port, B2 => n5656, ZN => n5151);
   U2289 : AOI22_X1 port map( A1 => REGISTERS_18_23_port, A2 => n5645, B1 => 
                           REGISTERS_27_23_port, B2 => n5646, ZN => n5150);
   U2290 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n5626, B1 => 
                           REGISTERS_30_23_port, B2 => n5619, ZN => n5149);
   U2291 : NAND4_X1 port map( A1 => n5152, A2 => n5151, A3 => n5150, A4 => 
                           n5149, ZN => n5158);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n5683, B1 => 
                           REGISTERS_25_23_port, B2 => n5693, ZN => n5156);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n5687, B1 => 
                           REGISTERS_26_23_port, B2 => n5657, ZN => n5155);
   U2294 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n5695, B1 => 
                           REGISTERS_24_23_port, B2 => n5653, ZN => n5154);
   U2295 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n5682, B1 => 
                           REGISTERS_16_23_port, B2 => n5700, ZN => n5153);
   U2296 : NAND4_X1 port map( A1 => n5156, A2 => n5155, A3 => n5154, A4 => 
                           n5153, ZN => n5157);
   U2297 : NOR2_X1 port map( A1 => n5158, A2 => n5157, ZN => n5170);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n5708, B1 => 
                           REGISTERS_0_23_port, B2 => n5720, ZN => n5162);
   U2299 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n5718, B1 => 
                           REGISTERS_4_23_port, B2 => n5610, ZN => n5161);
   U2300 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n5671, B1 => 
                           REGISTERS_3_23_port, B2 => n5717, ZN => n5160);
   U2301 : AOI22_X1 port map( A1 => REGISTERS_2_23_port, A2 => n5707, B1 => 
                           REGISTERS_6_23_port, B2 => n5709, ZN => n5159);
   U2302 : NAND4_X1 port map( A1 => n5162, A2 => n5161, A3 => n5160, A4 => 
                           n5159, ZN => n5168);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_14_23_port, A2 => n5670, B1 => 
                           REGISTERS_8_23_port, B2 => n5720, ZN => n5166);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n5718, B1 => 
                           REGISTERS_12_23_port, B2 => n5669, ZN => n5165);
   U2305 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n5717, B1 => 
                           REGISTERS_15_23_port, B2 => n5711, ZN => n5164);
   U2306 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n5708, B1 => 
                           REGISTERS_10_23_port, B2 => n5707, ZN => n5163);
   U2307 : NAND4_X1 port map( A1 => n5166, A2 => n5165, A3 => n5164, A4 => 
                           n5163, ZN => n5167);
   U2308 : AOI22_X1 port map( A1 => n5501, A2 => n5168, B1 => n5212, B2 => 
                           n5167, ZN => n5169);
   U2309 : OAI21_X1 port map( B1 => n5732, B2 => n5170, A => n5169, ZN => N408)
                           ;
   U2310 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n5687, B1 => 
                           REGISTERS_28_22_port, B2 => n5682, ZN => n5174);
   U2311 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n5698, B1 => 
                           REGISTERS_30_22_port, B2 => n5619, ZN => n5173);
   U2312 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n5700, B1 => 
                           REGISTERS_27_22_port, B2 => n5646, ZN => n5172);
   U2313 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n5625, B1 => 
                           REGISTERS_22_22_port, B2 => n5681, ZN => n5171);
   U2314 : NAND4_X1 port map( A1 => n5174, A2 => n5173, A3 => n5172, A4 => 
                           n5171, ZN => n5180);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n5699, B1 => 
                           REGISTERS_26_22_port, B2 => n5657, ZN => n5178);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n5683, B1 => 
                           REGISTERS_18_22_port, B2 => n5645, ZN => n5177);
   U2317 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n5685, B1 => 
                           REGISTERS_17_22_port, B2 => n5695, ZN => n5176);
   U2318 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n5626, B1 => 
                           REGISTERS_23_22_port, B2 => n5656, ZN => n5175);
   U2319 : NAND4_X1 port map( A1 => n5178, A2 => n5177, A3 => n5176, A4 => 
                           n5175, ZN => n5179);
   U2320 : NOR2_X1 port map( A1 => n5180, A2 => n5179, ZN => n5192);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n5717, B1 => 
                           REGISTERS_0_22_port, B2 => n5668, ZN => n5184);
   U2322 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n5721, B1 => 
                           REGISTERS_5_22_port, B2 => n5581, ZN => n5183);
   U2323 : AOI22_X1 port map( A1 => REGISTERS_6_22_port, A2 => n5709, B1 => 
                           REGISTERS_2_22_port, B2 => n5707, ZN => n5182);
   U2324 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n5719, B1 => 
                           REGISTERS_7_22_port, B2 => n5711, ZN => n5181);
   U2325 : NAND4_X1 port map( A1 => n5184, A2 => n5183, A3 => n5182, A4 => 
                           n5181, ZN => n5190);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n5669, B1 => 
                           REGISTERS_8_22_port, B2 => n5720, ZN => n5188);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n5671, B1 => 
                           REGISTERS_9_22_port, B2 => n5708, ZN => n5187);
   U2328 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n5718, B1 => 
                           REGISTERS_10_22_port, B2 => n5707, ZN => n5186);
   U2329 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n5717, B1 => 
                           REGISTERS_14_22_port, B2 => n5709, ZN => n5185);
   U2330 : NAND4_X1 port map( A1 => n5188, A2 => n5187, A3 => n5186, A4 => 
                           n5185, ZN => n5189);
   U2331 : AOI22_X1 port map( A1 => n5501, A2 => n5190, B1 => n5212, B2 => 
                           n5189, ZN => n5191);
   U2332 : OAI21_X1 port map( B1 => n5732, B2 => n5192, A => n5191, ZN => N407)
                           ;
   U2333 : AOI22_X1 port map( A1 => REGISTERS_27_21_port, A2 => n5694, B1 => 
                           REGISTERS_20_21_port, B2 => n5683, ZN => n5196);
   U2334 : AOI22_X1 port map( A1 => REGISTERS_23_21_port, A2 => n5697, B1 => 
                           REGISTERS_18_21_port, B2 => n5684, ZN => n5195);
   U2335 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n5626, B1 => 
                           REGISTERS_30_21_port, B2 => n5619, ZN => n5194);
   U2336 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n5687, B1 => 
                           REGISTERS_17_21_port, B2 => n5695, ZN => n5193);
   U2337 : NAND4_X1 port map( A1 => n5196, A2 => n5195, A3 => n5194, A4 => 
                           n5193, ZN => n5202);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n5681, B1 => 
                           REGISTERS_26_21_port, B2 => n5657, ZN => n5200);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n5655, B1 => 
                           REGISTERS_25_21_port, B2 => n5693, ZN => n5199);
   U2340 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n5682, B1 => 
                           REGISTERS_31_21_port, B2 => n5624, ZN => n5198);
   U2341 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n5653, B1 => 
                           REGISTERS_16_21_port, B2 => n5647, ZN => n5197);
   U2342 : NAND4_X1 port map( A1 => n5200, A2 => n5199, A3 => n5198, A4 => 
                           n5197, ZN => n5201);
   U2343 : NOR2_X1 port map( A1 => n5202, A2 => n5201, ZN => n5215);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n5671, B1 => 
                           REGISTERS_5_21_port, B2 => n5581, ZN => n5206);
   U2345 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n5720, B1 => 
                           REGISTERS_3_21_port, B2 => n5717, ZN => n5205);
   U2346 : AOI22_X1 port map( A1 => REGISTERS_6_21_port, A2 => n5670, B1 => 
                           REGISTERS_4_21_port, B2 => n5669, ZN => n5204);
   U2347 : AOI22_X1 port map( A1 => REGISTERS_2_21_port, A2 => n5707, B1 => 
                           REGISTERS_1_21_port, B2 => n5708, ZN => n5203);
   U2348 : NAND4_X1 port map( A1 => n5206, A2 => n5205, A3 => n5204, A4 => 
                           n5203, ZN => n5213);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_14_21_port, A2 => n5709, B1 => 
                           REGISTERS_13_21_port, B2 => n5581, ZN => n5210);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_10_21_port, A2 => n5707, B1 => 
                           REGISTERS_15_21_port, B2 => n5671, ZN => n5209);
   U2351 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n5708, B1 => 
                           REGISTERS_11_21_port, B2 => n5717, ZN => n5208);
   U2352 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n5720, B1 => 
                           REGISTERS_12_21_port, B2 => n5669, ZN => n5207);
   U2353 : NAND4_X1 port map( A1 => n5210, A2 => n5209, A3 => n5208, A4 => 
                           n5207, ZN => n5211);
   U2354 : AOI22_X1 port map( A1 => n5501, A2 => n5213, B1 => n5212, B2 => 
                           n5211, ZN => n5214);
   U2355 : OAI21_X1 port map( B1 => n5732, B2 => n5215, A => n5214, ZN => N406)
                           ;
   U2356 : AOI22_X1 port map( A1 => REGISTERS_31_20_port, A2 => n5698, B1 => 
                           REGISTERS_23_20_port, B2 => n5656, ZN => n5219);
   U2357 : AOI22_X1 port map( A1 => REGISTERS_22_20_port, A2 => n5681, B1 => 
                           REGISTERS_17_20_port, B2 => n5695, ZN => n5218);
   U2358 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n5682, B1 => 
                           REGISTERS_24_20_port, B2 => n5653, ZN => n5217);
   U2359 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n5646, B1 => 
                           REGISTERS_25_20_port, B2 => n5693, ZN => n5216);
   U2360 : NAND4_X1 port map( A1 => n5219, A2 => n5218, A3 => n5217, A4 => 
                           n5216, ZN => n5225);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n5685, B1 => 
                           REGISTERS_30_20_port, B2 => n5619, ZN => n5223);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_18_20_port, A2 => n5645, B1 => 
                           REGISTERS_21_20_port, B2 => n5687, ZN => n5222);
   U2363 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n5626, B1 => 
                           REGISTERS_26_20_port, B2 => n5657, ZN => n5221);
   U2364 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n5599, B1 => 
                           REGISTERS_16_20_port, B2 => n5647, ZN => n5220);
   U2365 : NAND4_X1 port map( A1 => n5223, A2 => n5222, A3 => n5221, A4 => 
                           n5220, ZN => n5224);
   U2366 : NOR2_X1 port map( A1 => n5225, A2 => n5224, ZN => n5237);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_6_20_port, A2 => n5709, B1 => 
                           REGISTERS_2_20_port, B2 => n5707, ZN => n5229);
   U2368 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n5671, B1 => 
                           REGISTERS_3_20_port, B2 => n5717, ZN => n5228);
   U2369 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n5719, B1 => 
                           REGISTERS_4_20_port, B2 => n5669, ZN => n5227);
   U2370 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n5720, B1 => 
                           REGISTERS_5_20_port, B2 => n5581, ZN => n5226);
   U2371 : NAND4_X1 port map( A1 => n5229, A2 => n5228, A3 => n5227, A4 => 
                           n5226, ZN => n5235);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n5720, B1 => 
                           REGISTERS_12_20_port, B2 => n5669, ZN => n5233);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n5671, B1 => 
                           REGISTERS_14_20_port, B2 => n5709, ZN => n5232);
   U2374 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n5708, B1 => 
                           REGISTERS_10_20_port, B2 => n5707, ZN => n5231);
   U2375 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n5717, B1 => 
                           REGISTERS_13_20_port, B2 => n5581, ZN => n5230);
   U2376 : NAND4_X1 port map( A1 => n5233, A2 => n5232, A3 => n5231, A4 => 
                           n5230, ZN => n5234);
   U2377 : AOI22_X1 port map( A1 => n5501, A2 => n5235, B1 => n5727, B2 => 
                           n5234, ZN => n5236);
   U2378 : OAI21_X1 port map( B1 => n5732, B2 => n5237, A => n5236, ZN => N405)
                           ;
   U2379 : AOI22_X1 port map( A1 => REGISTERS_22_19_port, A2 => n5594, B1 => 
                           REGISTERS_31_19_port, B2 => n5698, ZN => n5241);
   U2380 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n5656, B1 => 
                           REGISTERS_18_19_port, B2 => n5684, ZN => n5240);
   U2381 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n5686, B1 => 
                           REGISTERS_27_19_port, B2 => n5646, ZN => n5239);
   U2382 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n5687, B1 => 
                           REGISTERS_16_19_port, B2 => n5647, ZN => n5238);
   U2383 : NAND4_X1 port map( A1 => n5241, A2 => n5240, A3 => n5239, A4 => 
                           n5238, ZN => n5247);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_30_19_port, A2 => n5619, B1 => 
                           REGISTERS_29_19_port, B2 => n5685, ZN => n5245);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n5570, B1 => 
                           REGISTERS_25_19_port, B2 => n5693, ZN => n5244);
   U2386 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n5682, B1 => 
                           REGISTERS_20_19_port, B2 => n5683, ZN => n5243);
   U2387 : AOI22_X1 port map( A1 => REGISTERS_26_19_port, A2 => n5657, B1 => 
                           REGISTERS_24_19_port, B2 => n5653, ZN => n5242);
   U2388 : NAND4_X1 port map( A1 => n5245, A2 => n5244, A3 => n5243, A4 => 
                           n5242, ZN => n5246);
   U2389 : NOR2_X1 port map( A1 => n5247, A2 => n5246, ZN => n5259);
   U2390 : CLKBUF_X1 port map( A => n5302, Z => n5729);
   U2391 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n5671, B1 => 
                           REGISTERS_1_19_port, B2 => n5708, ZN => n5251);
   U2392 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n5718, B1 => 
                           REGISTERS_6_19_port, B2 => n5709, ZN => n5250);
   U2393 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n5668, B1 => 
                           REGISTERS_2_19_port, B2 => n5672, ZN => n5249);
   U2394 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n5669, B1 => 
                           REGISTERS_3_19_port, B2 => n5717, ZN => n5248);
   U2395 : NAND4_X1 port map( A1 => n5251, A2 => n5250, A3 => n5249, A4 => 
                           n5248, ZN => n5257);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_14_19_port, A2 => n5709, B1 => 
                           REGISTERS_8_19_port, B2 => n5720, ZN => n5255);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n5721, B1 => 
                           REGISTERS_13_19_port, B2 => n5581, ZN => n5254);
   U2398 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n5711, B1 => 
                           REGISTERS_10_19_port, B2 => n5707, ZN => n5253);
   U2399 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n5717, B1 => 
                           REGISTERS_9_19_port, B2 => n5708, ZN => n5252);
   U2400 : NAND4_X1 port map( A1 => n5255, A2 => n5254, A3 => n5253, A4 => 
                           n5252, ZN => n5256);
   U2401 : AOI22_X1 port map( A1 => n5729, A2 => n5257, B1 => n5727, B2 => 
                           n5256, ZN => n5258);
   U2402 : OAI21_X1 port map( B1 => n5732, B2 => n5259, A => n5258, ZN => N404)
                           ;
   U2403 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n5626, B1 => 
                           REGISTERS_22_18_port, B2 => n5681, ZN => n5263);
   U2404 : AOI22_X1 port map( A1 => REGISTERS_26_18_port, A2 => n5688, B1 => 
                           REGISTERS_24_18_port, B2 => n5653, ZN => n5262);
   U2405 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n5682, B1 => 
                           REGISTERS_18_18_port, B2 => n5645, ZN => n5261);
   U2406 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n5697, B1 => 
                           REGISTERS_20_18_port, B2 => n5683, ZN => n5260);
   U2407 : NAND4_X1 port map( A1 => n5263, A2 => n5262, A3 => n5261, A4 => 
                           n5260, ZN => n5269);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n5694, B1 => 
                           REGISTERS_25_18_port, B2 => n5693, ZN => n5267);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_30_18_port, A2 => n5619, B1 => 
                           REGISTERS_31_18_port, B2 => n5624, ZN => n5266);
   U2410 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n5647, B1 => 
                           REGISTERS_21_18_port, B2 => n5654, ZN => n5265);
   U2411 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n5570, B1 => 
                           REGISTERS_29_18_port, B2 => n5685, ZN => n5264);
   U2412 : NAND4_X1 port map( A1 => n5267, A2 => n5266, A3 => n5265, A4 => 
                           n5264, ZN => n5268);
   U2413 : NOR2_X1 port map( A1 => n5269, A2 => n5268, ZN => n5281);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n5708, B1 => 
                           REGISTERS_2_18_port, B2 => n5707, ZN => n5273);
   U2415 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n5720, B1 => 
                           REGISTERS_7_18_port, B2 => n5711, ZN => n5272);
   U2416 : AOI22_X1 port map( A1 => REGISTERS_6_18_port, A2 => n5670, B1 => 
                           REGISTERS_4_18_port, B2 => n5669, ZN => n5271);
   U2417 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n5718, B1 => 
                           REGISTERS_3_18_port, B2 => n5717, ZN => n5270);
   U2418 : NAND4_X1 port map( A1 => n5273, A2 => n5272, A3 => n5271, A4 => 
                           n5270, ZN => n5279);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_14_18_port, A2 => n5670, B1 => 
                           REGISTERS_10_18_port, B2 => n5707, ZN => n5277);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n5671, B1 => 
                           REGISTERS_11_18_port, B2 => n5717, ZN => n5276);
   U2421 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n5719, B1 => 
                           REGISTERS_12_18_port, B2 => n5669, ZN => n5275);
   U2422 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n5718, B1 => 
                           REGISTERS_8_18_port, B2 => n5720, ZN => n5274);
   U2423 : NAND4_X1 port map( A1 => n5277, A2 => n5276, A3 => n5275, A4 => 
                           n5274, ZN => n5278);
   U2424 : AOI22_X1 port map( A1 => n5729, A2 => n5279, B1 => n5727, B2 => 
                           n5278, ZN => n5280);
   U2425 : OAI21_X1 port map( B1 => n5732, B2 => n5281, A => n5280, ZN => N403)
                           ;
   U2426 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n5624, B1 => 
                           REGISTERS_30_17_port, B2 => n5619, ZN => n5285);
   U2427 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n5697, B1 => 
                           REGISTERS_28_17_port, B2 => n5648, ZN => n5284);
   U2428 : AOI22_X1 port map( A1 => REGISTERS_22_17_port, A2 => n5681, B1 => 
                           REGISTERS_27_17_port, B2 => n5646, ZN => n5283);
   U2429 : AOI22_X1 port map( A1 => REGISTERS_18_17_port, A2 => n5645, B1 => 
                           REGISTERS_25_17_port, B2 => n5625, ZN => n5282);
   U2430 : NAND4_X1 port map( A1 => n5285, A2 => n5284, A3 => n5283, A4 => 
                           n5282, ZN => n5291);
   U2431 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n5687, B1 => 
                           REGISTERS_17_17_port, B2 => n5695, ZN => n5289);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_26_17_port, A2 => n5657, B1 => 
                           REGISTERS_16_17_port, B2 => n5647, ZN => n5288);
   U2433 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n5655, B1 => 
                           REGISTERS_19_17_port, B2 => n5686, ZN => n5287);
   U2434 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n5683, B1 => 
                           REGISTERS_24_17_port, B2 => n5653, ZN => n5286);
   U2435 : NAND4_X1 port map( A1 => n5289, A2 => n5288, A3 => n5287, A4 => 
                           n5286, ZN => n5290);
   U2436 : NOR2_X1 port map( A1 => n5291, A2 => n5290, ZN => n5304);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n5670, B1 => 
                           REGISTERS_1_17_port, B2 => n5708, ZN => n5295);
   U2438 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n5671, B1 => 
                           REGISTERS_5_17_port, B2 => n5581, ZN => n5294);
   U2439 : AOI22_X1 port map( A1 => REGISTERS_2_17_port, A2 => n5707, B1 => 
                           REGISTERS_3_17_port, B2 => n5717, ZN => n5293);
   U2440 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n5610, B1 => 
                           REGISTERS_0_17_port, B2 => n5668, ZN => n5292);
   U2441 : NAND4_X1 port map( A1 => n5295, A2 => n5294, A3 => n5293, A4 => 
                           n5292, ZN => n5301);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n5721, B1 => 
                           REGISTERS_8_17_port, B2 => n5720, ZN => n5299);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n5710, B1 => 
                           REGISTERS_9_17_port, B2 => n5708, ZN => n5298);
   U2444 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n5718, B1 => 
                           REGISTERS_14_17_port, B2 => n5709, ZN => n5297);
   U2445 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n5707, B1 => 
                           REGISTERS_15_17_port, B2 => n5711, ZN => n5296);
   U2446 : NAND4_X1 port map( A1 => n5299, A2 => n5298, A3 => n5297, A4 => 
                           n5296, ZN => n5300);
   U2447 : AOI22_X1 port map( A1 => n5302, A2 => n5301, B1 => n5727, B2 => 
                           n5300, ZN => n5303);
   U2448 : OAI21_X1 port map( B1 => n5732, B2 => n5304, A => n5303, ZN => N402)
                           ;
   U2449 : AOI22_X1 port map( A1 => REGISTERS_26_16_port, A2 => n5657, B1 => 
                           REGISTERS_23_16_port, B2 => n5656, ZN => n5308);
   U2450 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n5648, B1 => 
                           REGISTERS_27_16_port, B2 => n5646, ZN => n5307);
   U2451 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n5655, B1 => 
                           REGISTERS_25_16_port, B2 => n5693, ZN => n5306);
   U2452 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n5681, B1 => 
                           REGISTERS_30_16_port, B2 => n5619, ZN => n5305);
   U2453 : NAND4_X1 port map( A1 => n5308, A2 => n5307, A3 => n5306, A4 => 
                           n5305, ZN => n5314);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n5695, B1 => 
                           REGISTERS_24_16_port, B2 => n5653, ZN => n5312);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n5700, B1 => 
                           REGISTERS_31_16_port, B2 => n5624, ZN => n5311);
   U2456 : AOI22_X1 port map( A1 => REGISTERS_18_16_port, A2 => n5684, B1 => 
                           REGISTERS_21_16_port, B2 => n5654, ZN => n5310);
   U2457 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n5626, B1 => 
                           REGISTERS_20_16_port, B2 => n5599, ZN => n5309);
   U2458 : NAND4_X1 port map( A1 => n5312, A2 => n5311, A3 => n5310, A4 => 
                           n5309, ZN => n5313);
   U2459 : NOR2_X1 port map( A1 => n5314, A2 => n5313, ZN => n5326);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n5720, B1 => 
                           REGISTERS_6_16_port, B2 => n5709, ZN => n5318);
   U2461 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n5671, B1 => 
                           REGISTERS_2_16_port, B2 => n5707, ZN => n5317);
   U2462 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n5708, B1 => 
                           REGISTERS_4_16_port, B2 => n5669, ZN => n5316);
   U2463 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n5717, B1 => 
                           REGISTERS_5_16_port, B2 => n5718, ZN => n5315);
   U2464 : NAND4_X1 port map( A1 => n5318, A2 => n5317, A3 => n5316, A4 => 
                           n5315, ZN => n5324);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n5717, B1 => 
                           REGISTERS_13_16_port, B2 => n5718, ZN => n5322);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n5669, B1 => 
                           REGISTERS_8_16_port, B2 => n5668, ZN => n5321);
   U2467 : AOI22_X1 port map( A1 => REGISTERS_14_16_port, A2 => n5670, B1 => 
                           REGISTERS_15_16_port, B2 => n5671, ZN => n5320);
   U2468 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n5672, B1 => 
                           REGISTERS_9_16_port, B2 => n5708, ZN => n5319);
   U2469 : NAND4_X1 port map( A1 => n5322, A2 => n5321, A3 => n5320, A4 => 
                           n5319, ZN => n5323);
   U2470 : AOI22_X1 port map( A1 => n5729, A2 => n5324, B1 => n5727, B2 => 
                           n5323, ZN => n5325);
   U2471 : OAI21_X1 port map( B1 => n5732, B2 => n5326, A => n5325, ZN => N401)
                           ;
   U2472 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n5687, B1 => 
                           REGISTERS_24_15_port, B2 => n5653, ZN => n5330);
   U2473 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n5599, B1 => 
                           REGISTERS_29_15_port, B2 => n5685, ZN => n5329);
   U2474 : AOI22_X1 port map( A1 => REGISTERS_18_15_port, A2 => n5645, B1 => 
                           REGISTERS_22_15_port, B2 => n5594, ZN => n5328);
   U2475 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n5624, B1 => 
                           REGISTERS_17_15_port, B2 => n5695, ZN => n5327);
   U2476 : NAND4_X1 port map( A1 => n5330, A2 => n5329, A3 => n5328, A4 => 
                           n5327, ZN => n5336);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n5646, B1 => 
                           REGISTERS_23_15_port, B2 => n5656, ZN => n5334);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n5647, B1 => 
                           REGISTERS_25_15_port, B2 => n5693, ZN => n5333);
   U2479 : AOI22_X1 port map( A1 => REGISTERS_26_15_port, A2 => n5657, B1 => 
                           REGISTERS_28_15_port, B2 => n5648, ZN => n5332);
   U2480 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n5686, B1 => 
                           REGISTERS_30_15_port, B2 => n5696, ZN => n5331);
   U2481 : NAND4_X1 port map( A1 => n5334, A2 => n5333, A3 => n5332, A4 => 
                           n5331, ZN => n5335);
   U2482 : NOR2_X1 port map( A1 => n5336, A2 => n5335, ZN => n5348);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n5721, B1 => 
                           REGISTERS_3_15_port, B2 => n5710, ZN => n5340);
   U2484 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n5719, B1 => 
                           REGISTERS_0_15_port, B2 => n5668, ZN => n5339);
   U2485 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n5581, B1 => 
                           REGISTERS_6_15_port, B2 => n5709, ZN => n5338);
   U2486 : AOI22_X1 port map( A1 => REGISTERS_2_15_port, A2 => n5672, B1 => 
                           REGISTERS_7_15_port, B2 => n5711, ZN => n5337);
   U2487 : NAND4_X1 port map( A1 => n5340, A2 => n5339, A3 => n5338, A4 => 
                           n5337, ZN => n5346);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n5720, B1 => 
                           REGISTERS_14_15_port, B2 => n5709, ZN => n5344);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n5718, B1 => 
                           REGISTERS_12_15_port, B2 => n5610, ZN => n5343);
   U2490 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n5671, B1 => 
                           REGISTERS_10_15_port, B2 => n5707, ZN => n5342);
   U2491 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n5708, B1 => 
                           REGISTERS_11_15_port, B2 => n5717, ZN => n5341);
   U2492 : NAND4_X1 port map( A1 => n5344, A2 => n5343, A3 => n5342, A4 => 
                           n5341, ZN => n5345);
   U2493 : AOI22_X1 port map( A1 => n5501, A2 => n5346, B1 => n5727, B2 => 
                           n5345, ZN => n5347);
   U2494 : OAI21_X1 port map( B1 => n5732, B2 => n5348, A => n5347, ZN => N400)
                           ;
   U2495 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n5594, B1 => 
                           REGISTERS_23_14_port, B2 => n5656, ZN => n5352);
   U2496 : AOI22_X1 port map( A1 => REGISTERS_31_14_port, A2 => n5624, B1 => 
                           REGISTERS_26_14_port, B2 => n5657, ZN => n5351);
   U2497 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n5695, B1 => 
                           REGISTERS_21_14_port, B2 => n5687, ZN => n5350);
   U2498 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n5686, B1 => 
                           REGISTERS_18_14_port, B2 => n5684, ZN => n5349);
   U2499 : NAND4_X1 port map( A1 => n5352, A2 => n5351, A3 => n5350, A4 => 
                           n5349, ZN => n5358);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n5683, B1 => 
                           REGISTERS_16_14_port, B2 => n5647, ZN => n5356);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n5648, B1 => 
                           REGISTERS_25_14_port, B2 => n5693, ZN => n5355);
   U2502 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n5655, B1 => 
                           REGISTERS_24_14_port, B2 => n5699, ZN => n5354);
   U2503 : AOI22_X1 port map( A1 => REGISTERS_30_14_port, A2 => n5619, B1 => 
                           REGISTERS_27_14_port, B2 => n5646, ZN => n5353);
   U2504 : NAND4_X1 port map( A1 => n5356, A2 => n5355, A3 => n5354, A4 => 
                           n5353, ZN => n5357);
   U2505 : NOR2_X1 port map( A1 => n5358, A2 => n5357, ZN => n5370);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n5717, B1 => 
                           REGISTERS_0_14_port, B2 => n5668, ZN => n5362);
   U2507 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n5708, B1 => 
                           REGISTERS_7_14_port, B2 => n5711, ZN => n5361);
   U2508 : AOI22_X1 port map( A1 => REGISTERS_6_14_port, A2 => n5670, B1 => 
                           REGISTERS_4_14_port, B2 => n5610, ZN => n5360);
   U2509 : AOI22_X1 port map( A1 => REGISTERS_2_14_port, A2 => n5672, B1 => 
                           REGISTERS_5_14_port, B2 => n5718, ZN => n5359);
   U2510 : NAND4_X1 port map( A1 => n5362, A2 => n5361, A3 => n5360, A4 => 
                           n5359, ZN => n5368);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n5668, B1 => 
                           REGISTERS_11_14_port, B2 => n5710, ZN => n5366);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_14_14_port, A2 => n5670, B1 => 
                           REGISTERS_12_14_port, B2 => n5610, ZN => n5365);
   U2513 : AOI22_X1 port map( A1 => REGISTERS_10_14_port, A2 => n5672, B1 => 
                           REGISTERS_9_14_port, B2 => n5708, ZN => n5364);
   U2514 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n5718, B1 => 
                           REGISTERS_15_14_port, B2 => n5711, ZN => n5363);
   U2515 : NAND4_X1 port map( A1 => n5366, A2 => n5365, A3 => n5364, A4 => 
                           n5363, ZN => n5367);
   U2516 : AOI22_X1 port map( A1 => n5501, A2 => n5368, B1 => n5727, B2 => 
                           n5367, ZN => n5369);
   U2517 : OAI21_X1 port map( B1 => n5732, B2 => n5370, A => n5369, ZN => N399)
                           ;
   U2518 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n5654, B1 => 
                           REGISTERS_27_13_port, B2 => n5646, ZN => n5374);
   U2519 : AOI22_X1 port map( A1 => REGISTERS_30_13_port, A2 => n5619, B1 => 
                           REGISTERS_22_13_port, B2 => n5681, ZN => n5373);
   U2520 : AOI22_X1 port map( A1 => REGISTERS_31_13_port, A2 => n5624, B1 => 
                           REGISTERS_19_13_port, B2 => n5626, ZN => n5372);
   U2521 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n5653, B1 => 
                           REGISTERS_20_13_port, B2 => n5683, ZN => n5371);
   U2522 : NAND4_X1 port map( A1 => n5374, A2 => n5373, A3 => n5372, A4 => 
                           n5371, ZN => n5380);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n5647, B1 => 
                           REGISTERS_17_13_port, B2 => n5695, ZN => n5378);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_18_13_port, A2 => n5645, B1 => 
                           REGISTERS_28_13_port, B2 => n5648, ZN => n5377);
   U2525 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n5656, B1 => 
                           REGISTERS_29_13_port, B2 => n5655, ZN => n5376);
   U2526 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n5625, B1 => 
                           REGISTERS_26_13_port, B2 => n5688, ZN => n5375);
   U2527 : NAND4_X1 port map( A1 => n5378, A2 => n5377, A3 => n5376, A4 => 
                           n5375, ZN => n5379);
   U2528 : NOR2_X1 port map( A1 => n5380, A2 => n5379, ZN => n5392);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_6_13_port, A2 => n5716, B1 => 
                           REGISTERS_1_13_port, B2 => n5708, ZN => n5384);
   U2530 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n5671, B1 => 
                           REGISTERS_2_13_port, B2 => n5707, ZN => n5383);
   U2531 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n5581, B1 => 
                           REGISTERS_4_13_port, B2 => n5610, ZN => n5382);
   U2532 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n5720, B1 => 
                           REGISTERS_3_13_port, B2 => n5710, ZN => n5381);
   U2533 : NAND4_X1 port map( A1 => n5384, A2 => n5383, A3 => n5382, A4 => 
                           n5381, ZN => n5390);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_14_13_port, A2 => n5709, B1 => 
                           REGISTERS_9_13_port, B2 => n5708, ZN => n5388);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n5718, B1 => 
                           REGISTERS_11_13_port, B2 => n5717, ZN => n5387);
   U2536 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n5671, B1 => 
                           REGISTERS_12_13_port, B2 => n5610, ZN => n5386);
   U2537 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n5720, B1 => 
                           REGISTERS_10_13_port, B2 => n5707, ZN => n5385);
   U2538 : NAND4_X1 port map( A1 => n5388, A2 => n5387, A3 => n5386, A4 => 
                           n5385, ZN => n5389);
   U2539 : AOI22_X1 port map( A1 => n5501, A2 => n5390, B1 => n5727, B2 => 
                           n5389, ZN => n5391);
   U2540 : OAI21_X1 port map( B1 => n5732, B2 => n5392, A => n5391, ZN => N398)
                           ;
   U2541 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n5699, B1 => 
                           REGISTERS_20_12_port, B2 => n5683, ZN => n5396);
   U2542 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n5693, B1 => 
                           REGISTERS_17_12_port, B2 => n5695, ZN => n5395);
   U2543 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n5654, B1 => 
                           REGISTERS_30_12_port, B2 => n5619, ZN => n5394);
   U2544 : AOI22_X1 port map( A1 => REGISTERS_31_12_port, A2 => n5698, B1 => 
                           REGISTERS_27_12_port, B2 => n5646, ZN => n5393);
   U2545 : NAND4_X1 port map( A1 => n5396, A2 => n5395, A3 => n5394, A4 => 
                           n5393, ZN => n5402);
   U2546 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n5655, B1 => 
                           REGISTERS_26_12_port, B2 => n5688, ZN => n5400);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n5648, B1 => 
                           REGISTERS_16_12_port, B2 => n5647, ZN => n5399);
   U2548 : AOI22_X1 port map( A1 => REGISTERS_19_12_port, A2 => n5686, B1 => 
                           REGISTERS_23_12_port, B2 => n5656, ZN => n5398);
   U2549 : AOI22_X1 port map( A1 => REGISTERS_22_12_port, A2 => n5681, B1 => 
                           REGISTERS_18_12_port, B2 => n5684, ZN => n5397);
   U2550 : NAND4_X1 port map( A1 => n5400, A2 => n5399, A3 => n5398, A4 => 
                           n5397, ZN => n5401);
   U2551 : NOR2_X1 port map( A1 => n5402, A2 => n5401, ZN => n5414);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n5721, B1 => 
                           REGISTERS_7_12_port, B2 => n5711, ZN => n5406);
   U2553 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n5708, B1 => 
                           REGISTERS_3_12_port, B2 => n5717, ZN => n5405);
   U2554 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n5581, B1 => 
                           REGISTERS_6_12_port, B2 => n5709, ZN => n5404);
   U2555 : AOI22_X1 port map( A1 => REGISTERS_2_12_port, A2 => n5672, B1 => 
                           REGISTERS_0_12_port, B2 => n5668, ZN => n5403);
   U2556 : NAND4_X1 port map( A1 => n5406, A2 => n5405, A3 => n5404, A4 => 
                           n5403, ZN => n5412);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n5708, B1 => 
                           REGISTERS_12_12_port, B2 => n5610, ZN => n5410);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n5720, B1 => 
                           REGISTERS_13_12_port, B2 => n5718, ZN => n5409);
   U2559 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n5710, B1 => 
                           REGISTERS_15_12_port, B2 => n5671, ZN => n5408);
   U2560 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n5670, B1 => 
                           REGISTERS_10_12_port, B2 => n5707, ZN => n5407);
   U2561 : NAND4_X1 port map( A1 => n5410, A2 => n5409, A3 => n5408, A4 => 
                           n5407, ZN => n5411);
   U2562 : AOI22_X1 port map( A1 => n5501, A2 => n5412, B1 => n5727, B2 => 
                           n5411, ZN => n5413);
   U2563 : OAI21_X1 port map( B1 => n5732, B2 => n5414, A => n5413, ZN => N397)
                           ;
   U2564 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n5686, B1 => 
                           REGISTERS_17_11_port, B2 => n5695, ZN => n5418);
   U2565 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n5693, B1 => 
                           REGISTERS_29_11_port, B2 => n5685, ZN => n5417);
   U2566 : AOI22_X1 port map( A1 => REGISTERS_22_11_port, A2 => n5594, B1 => 
                           REGISTERS_31_11_port, B2 => n5698, ZN => n5416);
   U2567 : AOI22_X1 port map( A1 => REGISTERS_26_11_port, A2 => n5657, B1 => 
                           REGISTERS_20_11_port, B2 => n5683, ZN => n5415);
   U2568 : NAND4_X1 port map( A1 => n5418, A2 => n5417, A3 => n5416, A4 => 
                           n5415, ZN => n5424);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_30_11_port, A2 => n5619, B1 => 
                           REGISTERS_28_11_port, B2 => n5682, ZN => n5422);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_18_11_port, A2 => n5645, B1 => 
                           REGISTERS_24_11_port, B2 => n5653, ZN => n5421);
   U2571 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n5647, B1 => 
                           REGISTERS_23_11_port, B2 => n5697, ZN => n5420);
   U2572 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n5687, B1 => 
                           REGISTERS_27_11_port, B2 => n5694, ZN => n5419);
   U2573 : NAND4_X1 port map( A1 => n5422, A2 => n5421, A3 => n5420, A4 => 
                           n5419, ZN => n5423);
   U2574 : NOR2_X1 port map( A1 => n5424, A2 => n5423, ZN => n5436);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n5720, B1 => 
                           REGISTERS_2_11_port, B2 => n5707, ZN => n5428);
   U2576 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n5717, B1 => 
                           REGISTERS_7_11_port, B2 => n5711, ZN => n5427);
   U2577 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n5708, B1 => 
                           REGISTERS_4_11_port, B2 => n5610, ZN => n5426);
   U2578 : AOI22_X1 port map( A1 => REGISTERS_6_11_port, A2 => n5670, B1 => 
                           REGISTERS_5_11_port, B2 => n5718, ZN => n5425);
   U2579 : NAND4_X1 port map( A1 => n5428, A2 => n5427, A3 => n5426, A4 => 
                           n5425, ZN => n5434);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_15_11_port, A2 => n5671, B1 => 
                           REGISTERS_12_11_port, B2 => n5610, ZN => n5432);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n5718, B1 => 
                           REGISTERS_11_11_port, B2 => n5717, ZN => n5431);
   U2582 : AOI22_X1 port map( A1 => REGISTERS_14_11_port, A2 => n5670, B1 => 
                           REGISTERS_9_11_port, B2 => n5708, ZN => n5430);
   U2583 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n5672, B1 => 
                           REGISTERS_8_11_port, B2 => n5668, ZN => n5429);
   U2584 : NAND4_X1 port map( A1 => n5432, A2 => n5431, A3 => n5430, A4 => 
                           n5429, ZN => n5433);
   U2585 : AOI22_X1 port map( A1 => n5501, A2 => n5434, B1 => n5727, B2 => 
                           n5433, ZN => n5435);
   U2586 : OAI21_X1 port map( B1 => n5732, B2 => n5436, A => n5435, ZN => N396)
                           ;
   U2587 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n5695, B1 => 
                           REGISTERS_22_10_port, B2 => n5681, ZN => n5440);
   U2588 : AOI22_X1 port map( A1 => REGISTERS_26_10_port, A2 => n5657, B1 => 
                           REGISTERS_25_10_port, B2 => n5625, ZN => n5439);
   U2589 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n5698, B1 => 
                           REGISTERS_23_10_port, B2 => n5656, ZN => n5438);
   U2590 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n5699, B1 => 
                           REGISTERS_30_10_port, B2 => n5619, ZN => n5437);
   U2591 : NAND4_X1 port map( A1 => n5440, A2 => n5439, A3 => n5438, A4 => 
                           n5437, ZN => n5446);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n5686, B1 => 
                           REGISTERS_21_10_port, B2 => n5687, ZN => n5444);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n5648, B1 => 
                           REGISTERS_18_10_port, B2 => n5684, ZN => n5443);
   U2594 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n5685, B1 => 
                           REGISTERS_16_10_port, B2 => n5647, ZN => n5442);
   U2595 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n5646, B1 => 
                           REGISTERS_20_10_port, B2 => n5599, ZN => n5441);
   U2596 : NAND4_X1 port map( A1 => n5444, A2 => n5443, A3 => n5442, A4 => 
                           n5441, ZN => n5445);
   U2597 : NOR2_X1 port map( A1 => n5446, A2 => n5445, ZN => n5458);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n5718, B1 => 
                           REGISTERS_1_10_port, B2 => n5708, ZN => n5450);
   U2599 : AOI22_X1 port map( A1 => REGISTERS_6_10_port, A2 => n5670, B1 => 
                           REGISTERS_7_10_port, B2 => n5671, ZN => n5449);
   U2600 : AOI22_X1 port map( A1 => REGISTERS_2_10_port, A2 => n5672, B1 => 
                           REGISTERS_0_10_port, B2 => n5668, ZN => n5448);
   U2601 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n5721, B1 => 
                           REGISTERS_3_10_port, B2 => n5717, ZN => n5447);
   U2602 : NAND4_X1 port map( A1 => n5450, A2 => n5449, A3 => n5448, A4 => 
                           n5447, ZN => n5456);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n5708, B1 => 
                           REGISTERS_11_10_port, B2 => n5710, ZN => n5454);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n5669, B1 => 
                           REGISTERS_8_10_port, B2 => n5668, ZN => n5453);
   U2605 : AOI22_X1 port map( A1 => REGISTERS_14_10_port, A2 => n5670, B1 => 
                           REGISTERS_13_10_port, B2 => n5718, ZN => n5452);
   U2606 : AOI22_X1 port map( A1 => REGISTERS_10_10_port, A2 => n5707, B1 => 
                           REGISTERS_15_10_port, B2 => n5711, ZN => n5451);
   U2607 : NAND4_X1 port map( A1 => n5454, A2 => n5453, A3 => n5452, A4 => 
                           n5451, ZN => n5455);
   U2608 : AOI22_X1 port map( A1 => n5501, A2 => n5456, B1 => n5727, B2 => 
                           n5455, ZN => n5457);
   U2609 : OAI21_X1 port map( B1 => n5732, B2 => n5458, A => n5457, ZN => N395)
                           ;
   U2610 : AOI22_X1 port map( A1 => REGISTERS_18_9_port, A2 => n5684, B1 => 
                           REGISTERS_24_9_port, B2 => n5653, ZN => n5462);
   U2611 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n5656, B1 => 
                           REGISTERS_29_9_port, B2 => n5685, ZN => n5461);
   U2612 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n5654, B1 => 
                           REGISTERS_30_9_port, B2 => n5619, ZN => n5460);
   U2613 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n5698, B1 => 
                           REGISTERS_20_9_port, B2 => n5683, ZN => n5459);
   U2614 : NAND4_X1 port map( A1 => n5462, A2 => n5461, A3 => n5460, A4 => 
                           n5459, ZN => n5468);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_22_9_port, A2 => n5594, B1 => 
                           REGISTERS_27_9_port, B2 => n5646, ZN => n5466);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_26_9_port, A2 => n5657, B1 => 
                           REGISTERS_19_9_port, B2 => n5686, ZN => n5465);
   U2617 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n5648, B1 => 
                           REGISTERS_17_9_port, B2 => n5570, ZN => n5464);
   U2618 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n5647, B1 => 
                           REGISTERS_25_9_port, B2 => n5693, ZN => n5463);
   U2619 : NAND4_X1 port map( A1 => n5466, A2 => n5465, A3 => n5464, A4 => 
                           n5463, ZN => n5467);
   U2620 : NOR2_X1 port map( A1 => n5468, A2 => n5467, ZN => n5480);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_6_9_port, A2 => n5670, B1 => 
                           REGISTERS_4_9_port, B2 => n5610, ZN => n5472);
   U2622 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n5671, B1 => 
                           REGISTERS_0_9_port, B2 => n5668, ZN => n5471);
   U2623 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n5708, B1 => 
                           REGISTERS_5_9_port, B2 => n5718, ZN => n5470);
   U2624 : AOI22_X1 port map( A1 => REGISTERS_2_9_port, A2 => n5707, B1 => 
                           REGISTERS_3_9_port, B2 => n5717, ZN => n5469);
   U2625 : NAND4_X1 port map( A1 => n5472, A2 => n5471, A3 => n5470, A4 => 
                           n5469, ZN => n5478);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n5718, B1 => 
                           REGISTERS_11_9_port, B2 => n5710, ZN => n5476);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_10_9_port, A2 => n5707, B1 => 
                           REGISTERS_12_9_port, B2 => n5610, ZN => n5475);
   U2628 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n5708, B1 => 
                           REGISTERS_14_9_port, B2 => n5716, ZN => n5474);
   U2629 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n5671, B1 => 
                           REGISTERS_8_9_port, B2 => n5668, ZN => n5473);
   U2630 : NAND4_X1 port map( A1 => n5476, A2 => n5475, A3 => n5474, A4 => 
                           n5473, ZN => n5477);
   U2631 : AOI22_X1 port map( A1 => n5501, A2 => n5478, B1 => n5727, B2 => 
                           n5477, ZN => n5479);
   U2632 : OAI21_X1 port map( B1 => n5732, B2 => n5480, A => n5479, ZN => N394)
                           ;
   U2633 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n5648, B1 => 
                           REGISTERS_30_8_port, B2 => n5619, ZN => n5484);
   U2634 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n5687, B1 => 
                           REGISTERS_17_8_port, B2 => n5695, ZN => n5483);
   U2635 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n5646, B1 => 
                           REGISTERS_22_8_port, B2 => n5681, ZN => n5482);
   U2636 : AOI22_X1 port map( A1 => REGISTERS_26_8_port, A2 => n5688, B1 => 
                           REGISTERS_18_8_port, B2 => n5684, ZN => n5481);
   U2637 : NAND4_X1 port map( A1 => n5484, A2 => n5483, A3 => n5482, A4 => 
                           n5481, ZN => n5490);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n5700, B1 => 
                           REGISTERS_29_8_port, B2 => n5685, ZN => n5488);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n5653, B1 => 
                           REGISTERS_19_8_port, B2 => n5626, ZN => n5487);
   U2640 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n5656, B1 => 
                           REGISTERS_25_8_port, B2 => n5625, ZN => n5486);
   U2641 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n5599, B1 => 
                           REGISTERS_31_8_port, B2 => n5698, ZN => n5485);
   U2642 : NAND4_X1 port map( A1 => n5488, A2 => n5487, A3 => n5486, A4 => 
                           n5485, ZN => n5489);
   U2643 : NOR2_X1 port map( A1 => n5490, A2 => n5489, ZN => n5503);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n5720, B1 => 
                           REGISTERS_4_8_port, B2 => n5610, ZN => n5494);
   U2645 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n5581, B1 => 
                           REGISTERS_1_8_port, B2 => n5708, ZN => n5493);
   U2646 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n5711, B1 => 
                           REGISTERS_2_8_port, B2 => n5672, ZN => n5492);
   U2647 : AOI22_X1 port map( A1 => REGISTERS_6_8_port, A2 => n5670, B1 => 
                           REGISTERS_3_8_port, B2 => n5710, ZN => n5491);
   U2648 : NAND4_X1 port map( A1 => n5494, A2 => n5493, A3 => n5492, A4 => 
                           n5491, ZN => n5500);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n5718, B1 => 
                           REGISTERS_10_8_port, B2 => n5707, ZN => n5498);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n5671, B1 => 
                           REGISTERS_8_8_port, B2 => n5668, ZN => n5497);
   U2651 : AOI22_X1 port map( A1 => REGISTERS_14_8_port, A2 => n5670, B1 => 
                           REGISTERS_11_8_port, B2 => n5710, ZN => n5496);
   U2652 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n5719, B1 => 
                           REGISTERS_12_8_port, B2 => n5721, ZN => n5495);
   U2653 : NAND4_X1 port map( A1 => n5498, A2 => n5497, A3 => n5496, A4 => 
                           n5495, ZN => n5499);
   U2654 : AOI22_X1 port map( A1 => n5501, A2 => n5500, B1 => n5727, B2 => 
                           n5499, ZN => n5502);
   U2655 : OAI21_X1 port map( B1 => n5732, B2 => n5503, A => n5502, ZN => N393)
                           ;
   U2656 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n5654, B1 => 
                           REGISTERS_27_7_port, B2 => n5646, ZN => n5507);
   U2657 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n5599, B1 => 
                           REGISTERS_25_7_port, B2 => n5625, ZN => n5506);
   U2658 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n5700, B1 => 
                           REGISTERS_30_7_port, B2 => n5619, ZN => n5505);
   U2659 : AOI22_X1 port map( A1 => REGISTERS_26_7_port, A2 => n5688, B1 => 
                           REGISTERS_18_7_port, B2 => n5684, ZN => n5504);
   U2660 : NAND4_X1 port map( A1 => n5507, A2 => n5506, A3 => n5505, A4 => 
                           n5504, ZN => n5513);
   U2661 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n5682, B1 => 
                           REGISTERS_24_7_port, B2 => n5653, ZN => n5511);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n5570, B1 => 
                           REGISTERS_31_7_port, B2 => n5698, ZN => n5510);
   U2663 : AOI22_X1 port map( A1 => REGISTERS_23_7_port, A2 => n5656, B1 => 
                           REGISTERS_19_7_port, B2 => n5626, ZN => n5509);
   U2664 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n5594, B1 => 
                           REGISTERS_29_7_port, B2 => n5685, ZN => n5508);
   U2665 : NAND4_X1 port map( A1 => n5511, A2 => n5510, A3 => n5509, A4 => 
                           n5508, ZN => n5512);
   U2666 : NOR2_X1 port map( A1 => n5513, A2 => n5512, ZN => n5525);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n5717, B1 => 
                           REGISTERS_7_7_port, B2 => n5671, ZN => n5517);
   U2668 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n5718, B1 => 
                           REGISTERS_4_7_port, B2 => n5721, ZN => n5516);
   U2669 : AOI22_X1 port map( A1 => REGISTERS_2_7_port, A2 => n5672, B1 => 
                           REGISTERS_1_7_port, B2 => n5719, ZN => n5515);
   U2670 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n5720, B1 => 
                           REGISTERS_6_7_port, B2 => n5716, ZN => n5514);
   U2671 : NAND4_X1 port map( A1 => n5517, A2 => n5516, A3 => n5515, A4 => 
                           n5514, ZN => n5523);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n5708, B1 => 
                           REGISTERS_14_7_port, B2 => n5716, ZN => n5521);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n5717, B1 => 
                           REGISTERS_15_7_port, B2 => n5671, ZN => n5520);
   U2674 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n5669, B1 => 
                           REGISTERS_13_7_port, B2 => n5718, ZN => n5519);
   U2675 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n5720, B1 => 
                           REGISTERS_10_7_port, B2 => n5672, ZN => n5518);
   U2676 : NAND4_X1 port map( A1 => n5521, A2 => n5520, A3 => n5519, A4 => 
                           n5518, ZN => n5522);
   U2677 : AOI22_X1 port map( A1 => n5729, A2 => n5523, B1 => n5727, B2 => 
                           n5522, ZN => n5524);
   U2678 : OAI21_X1 port map( B1 => n5732, B2 => n5525, A => n5524, ZN => N392)
                           ;
   U2679 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n5655, B1 => 
                           REGISTERS_21_6_port, B2 => n5687, ZN => n5529);
   U2680 : AOI22_X1 port map( A1 => REGISTERS_18_6_port, A2 => n5645, B1 => 
                           REGISTERS_19_6_port, B2 => n5626, ZN => n5528);
   U2681 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n5695, B1 => 
                           REGISTERS_28_6_port, B2 => n5682, ZN => n5527);
   U2682 : AOI22_X1 port map( A1 => REGISTERS_22_6_port, A2 => n5681, B1 => 
                           REGISTERS_20_6_port, B2 => n5683, ZN => n5526);
   U2683 : NAND4_X1 port map( A1 => n5529, A2 => n5528, A3 => n5527, A4 => 
                           n5526, ZN => n5535);
   U2684 : AOI22_X1 port map( A1 => REGISTERS_26_6_port, A2 => n5688, B1 => 
                           REGISTERS_16_6_port, B2 => n5647, ZN => n5533);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n5625, B1 => 
                           REGISTERS_23_6_port, B2 => n5656, ZN => n5532);
   U2686 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n5653, B1 => 
                           REGISTERS_30_6_port, B2 => n5696, ZN => n5531);
   U2687 : AOI22_X1 port map( A1 => REGISTERS_31_6_port, A2 => n5624, B1 => 
                           REGISTERS_27_6_port, B2 => n5694, ZN => n5530);
   U2688 : NAND4_X1 port map( A1 => n5533, A2 => n5532, A3 => n5531, A4 => 
                           n5530, ZN => n5534);
   U2689 : NOR2_X1 port map( A1 => n5535, A2 => n5534, ZN => n5547);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n5720, B1 => 
                           REGISTERS_3_6_port, B2 => n5710, ZN => n5539);
   U2691 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n5718, B1 => 
                           REGISTERS_7_6_port, B2 => n5671, ZN => n5538);
   U2692 : AOI22_X1 port map( A1 => REGISTERS_6_6_port, A2 => n5670, B1 => 
                           REGISTERS_1_6_port, B2 => n5719, ZN => n5537);
   U2693 : AOI22_X1 port map( A1 => REGISTERS_2_6_port, A2 => n5707, B1 => 
                           REGISTERS_4_6_port, B2 => n5721, ZN => n5536);
   U2694 : NAND4_X1 port map( A1 => n5539, A2 => n5538, A3 => n5537, A4 => 
                           n5536, ZN => n5545);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n5671, B1 => 
                           REGISTERS_12_6_port, B2 => n5721, ZN => n5543);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n5717, B1 => 
                           REGISTERS_14_6_port, B2 => n5716, ZN => n5542);
   U2697 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n5708, B1 => 
                           REGISTERS_10_6_port, B2 => n5672, ZN => n5541);
   U2698 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n5718, B1 => 
                           REGISTERS_8_6_port, B2 => n5720, ZN => n5540);
   U2699 : NAND4_X1 port map( A1 => n5543, A2 => n5542, A3 => n5541, A4 => 
                           n5540, ZN => n5544);
   U2700 : AOI22_X1 port map( A1 => n5729, A2 => n5545, B1 => n5727, B2 => 
                           n5544, ZN => n5546);
   U2701 : OAI21_X1 port map( B1 => n5732, B2 => n5547, A => n5546, ZN => N391)
                           ;
   U2702 : AOI22_X1 port map( A1 => REGISTERS_30_5_port, A2 => n5696, B1 => 
                           REGISTERS_22_5_port, B2 => n5681, ZN => n5551);
   U2703 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n5697, B1 => 
                           REGISTERS_26_5_port, B2 => n5657, ZN => n5550);
   U2704 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n5654, B1 => 
                           REGISTERS_19_5_port, B2 => n5626, ZN => n5549);
   U2705 : AOI22_X1 port map( A1 => REGISTERS_18_5_port, A2 => n5645, B1 => 
                           REGISTERS_28_5_port, B2 => n5682, ZN => n5548);
   U2706 : NAND4_X1 port map( A1 => n5551, A2 => n5550, A3 => n5549, A4 => 
                           n5548, ZN => n5557);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n5599, B1 => 
                           REGISTERS_24_5_port, B2 => n5653, ZN => n5555);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n5625, B1 => 
                           REGISTERS_29_5_port, B2 => n5685, ZN => n5554);
   U2709 : AOI22_X1 port map( A1 => REGISTERS_31_5_port, A2 => n5624, B1 => 
                           REGISTERS_16_5_port, B2 => n5700, ZN => n5553);
   U2710 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n5646, B1 => 
                           REGISTERS_17_5_port, B2 => n5570, ZN => n5552);
   U2711 : NAND4_X1 port map( A1 => n5555, A2 => n5554, A3 => n5553, A4 => 
                           n5552, ZN => n5556);
   U2712 : NOR2_X1 port map( A1 => n5557, A2 => n5556, ZN => n5569);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n5708, B1 => 
                           REGISTERS_4_5_port, B2 => n5721, ZN => n5561);
   U2714 : AOI22_X1 port map( A1 => REGISTERS_3_5_port, A2 => n5717, B1 => 
                           REGISTERS_0_5_port, B2 => n5720, ZN => n5560);
   U2715 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n5671, B1 => 
                           REGISTERS_5_5_port, B2 => n5718, ZN => n5559);
   U2716 : AOI22_X1 port map( A1 => REGISTERS_2_5_port, A2 => n5672, B1 => 
                           REGISTERS_6_5_port, B2 => n5716, ZN => n5558);
   U2717 : NAND4_X1 port map( A1 => n5561, A2 => n5560, A3 => n5559, A4 => 
                           n5558, ZN => n5567);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n5669, B1 => 
                           REGISTERS_9_5_port, B2 => n5719, ZN => n5565);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n5718, B1 => 
                           REGISTERS_10_5_port, B2 => n5672, ZN => n5564);
   U2720 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n5720, B1 => 
                           REGISTERS_14_5_port, B2 => n5716, ZN => n5563);
   U2721 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n5671, B1 => 
                           REGISTERS_11_5_port, B2 => n5710, ZN => n5562);
   U2722 : NAND4_X1 port map( A1 => n5565, A2 => n5564, A3 => n5563, A4 => 
                           n5562, ZN => n5566);
   U2723 : AOI22_X1 port map( A1 => n5729, A2 => n5567, B1 => n5727, B2 => 
                           n5566, ZN => n5568);
   U2724 : OAI21_X1 port map( B1 => n5732, B2 => n5569, A => n5568, ZN => N390)
                           ;
   U2725 : AOI22_X1 port map( A1 => REGISTERS_31_4_port, A2 => n5624, B1 => 
                           REGISTERS_27_4_port, B2 => n5646, ZN => n5574);
   U2726 : AOI22_X1 port map( A1 => REGISTERS_26_4_port, A2 => n5688, B1 => 
                           REGISTERS_18_4_port, B2 => n5684, ZN => n5573);
   U2727 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n5654, B1 => 
                           REGISTERS_29_4_port, B2 => n5685, ZN => n5572);
   U2728 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n5570, B1 => 
                           REGISTERS_25_4_port, B2 => n5625, ZN => n5571);
   U2729 : NAND4_X1 port map( A1 => n5574, A2 => n5573, A3 => n5572, A4 => 
                           n5571, ZN => n5580);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_30_4_port, A2 => n5619, B1 => 
                           REGISTERS_24_4_port, B2 => n5653, ZN => n5578);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n5700, B1 => 
                           REGISTERS_23_4_port, B2 => n5656, ZN => n5577);
   U2732 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n5594, B1 => 
                           REGISTERS_20_4_port, B2 => n5599, ZN => n5576);
   U2733 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n5682, B1 => 
                           REGISTERS_19_4_port, B2 => n5626, ZN => n5575);
   U2734 : NAND4_X1 port map( A1 => n5578, A2 => n5577, A3 => n5576, A4 => 
                           n5575, ZN => n5579);
   U2735 : NOR2_X1 port map( A1 => n5580, A2 => n5579, ZN => n5593);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_2_4_port, A2 => n5707, B1 => 
                           REGISTERS_0_4_port, B2 => n5720, ZN => n5585);
   U2737 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n5711, B1 => 
                           REGISTERS_5_4_port, B2 => n5581, ZN => n5584);
   U2738 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n5721, B1 => 
                           REGISTERS_1_4_port, B2 => n5719, ZN => n5583);
   U2739 : AOI22_X1 port map( A1 => REGISTERS_6_4_port, A2 => n5709, B1 => 
                           REGISTERS_3_4_port, B2 => n5710, ZN => n5582);
   U2740 : NAND4_X1 port map( A1 => n5585, A2 => n5584, A3 => n5583, A4 => 
                           n5582, ZN => n5591);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n5708, B1 => 
                           REGISTERS_10_4_port, B2 => n5672, ZN => n5589);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n5671, B1 => 
                           REGISTERS_14_4_port, B2 => n5716, ZN => n5588);
   U2743 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n5610, B1 => 
                           REGISTERS_8_4_port, B2 => n5720, ZN => n5587);
   U2744 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n5710, B1 => 
                           REGISTERS_13_4_port, B2 => n5718, ZN => n5586);
   U2745 : NAND4_X1 port map( A1 => n5589, A2 => n5588, A3 => n5587, A4 => 
                           n5586, ZN => n5590);
   U2746 : AOI22_X1 port map( A1 => n5729, A2 => n5591, B1 => n5727, B2 => 
                           n5590, ZN => n5592);
   U2747 : OAI21_X1 port map( B1 => n5732, B2 => n5593, A => n5592, ZN => N389)
                           ;
   U2748 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n5653, B1 => 
                           REGISTERS_19_3_port, B2 => n5626, ZN => n5598);
   U2749 : AOI22_X1 port map( A1 => REGISTERS_26_3_port, A2 => n5688, B1 => 
                           REGISTERS_17_3_port, B2 => n5695, ZN => n5597);
   U2750 : AOI22_X1 port map( A1 => REGISTERS_22_3_port, A2 => n5594, B1 => 
                           REGISTERS_27_3_port, B2 => n5646, ZN => n5596);
   U2751 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n5697, B1 => 
                           REGISTERS_31_3_port, B2 => n5698, ZN => n5595);
   U2752 : NAND4_X1 port map( A1 => n5598, A2 => n5597, A3 => n5596, A4 => 
                           n5595, ZN => n5605);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n5682, B1 => 
                           REGISTERS_16_3_port, B2 => n5647, ZN => n5603);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n5655, B1 => 
                           REGISTERS_25_3_port, B2 => n5693, ZN => n5602);
   U2755 : AOI22_X1 port map( A1 => REGISTERS_18_3_port, A2 => n5684, B1 => 
                           REGISTERS_30_3_port, B2 => n5696, ZN => n5601);
   U2756 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n5599, B1 => 
                           REGISTERS_21_3_port, B2 => n5687, ZN => n5600);
   U2757 : NAND4_X1 port map( A1 => n5603, A2 => n5602, A3 => n5601, A4 => 
                           n5600, ZN => n5604);
   U2758 : NOR2_X1 port map( A1 => n5605, A2 => n5604, ZN => n5618);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n5707, B1 => 
                           REGISTERS_6_3_port, B2 => n5716, ZN => n5609);
   U2760 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n5669, B1 => 
                           REGISTERS_1_3_port, B2 => n5719, ZN => n5608);
   U2761 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n5717, B1 => 
                           REGISTERS_5_3_port, B2 => n5718, ZN => n5607);
   U2762 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n5720, B1 => 
                           REGISTERS_7_3_port, B2 => n5671, ZN => n5606);
   U2763 : NAND4_X1 port map( A1 => n5609, A2 => n5608, A3 => n5607, A4 => 
                           n5606, ZN => n5616);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n5718, B1 => 
                           REGISTERS_14_3_port, B2 => n5716, ZN => n5614);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n5717, B1 => 
                           REGISTERS_9_3_port, B2 => n5719, ZN => n5613);
   U2766 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n5720, B1 => 
                           REGISTERS_15_3_port, B2 => n5671, ZN => n5612);
   U2767 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n5610, B1 => 
                           REGISTERS_10_3_port, B2 => n5672, ZN => n5611);
   U2768 : NAND4_X1 port map( A1 => n5614, A2 => n5613, A3 => n5612, A4 => 
                           n5611, ZN => n5615);
   U2769 : AOI22_X1 port map( A1 => n5729, A2 => n5616, B1 => n5727, B2 => 
                           n5615, ZN => n5617);
   U2770 : OAI21_X1 port map( B1 => n5732, B2 => n5618, A => n5617, ZN => N388)
                           ;
   U2771 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n5697, B1 => 
                           REGISTERS_30_2_port, B2 => n5619, ZN => n5623);
   U2772 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n5694, B1 => 
                           REGISTERS_20_2_port, B2 => n5683, ZN => n5622);
   U2773 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n5654, B1 => 
                           REGISTERS_22_2_port, B2 => n5681, ZN => n5621);
   U2774 : AOI22_X1 port map( A1 => REGISTERS_26_2_port, A2 => n5688, B1 => 
                           REGISTERS_29_2_port, B2 => n5685, ZN => n5620);
   U2775 : NAND4_X1 port map( A1 => n5623, A2 => n5622, A3 => n5621, A4 => 
                           n5620, ZN => n5632);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n5624, B1 => 
                           REGISTERS_28_2_port, B2 => n5682, ZN => n5630);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n5700, B1 => 
                           REGISTERS_18_2_port, B2 => n5684, ZN => n5629);
   U2778 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n5625, B1 => 
                           REGISTERS_24_2_port, B2 => n5699, ZN => n5628);
   U2779 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n5695, B1 => 
                           REGISTERS_19_2_port, B2 => n5626, ZN => n5627);
   U2780 : NAND4_X1 port map( A1 => n5630, A2 => n5629, A3 => n5628, A4 => 
                           n5627, ZN => n5631);
   U2781 : NOR2_X1 port map( A1 => n5632, A2 => n5631, ZN => n5644);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n5711, B1 => 
                           REGISTERS_0_2_port, B2 => n5668, ZN => n5636);
   U2783 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n5717, B1 => 
                           REGISTERS_6_2_port, B2 => n5716, ZN => n5635);
   U2784 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n5669, B1 => 
                           REGISTERS_1_2_port, B2 => n5719, ZN => n5634);
   U2785 : AOI22_X1 port map( A1 => REGISTERS_2_2_port, A2 => n5707, B1 => 
                           REGISTERS_5_2_port, B2 => n5718, ZN => n5633);
   U2786 : NAND4_X1 port map( A1 => n5636, A2 => n5635, A3 => n5634, A4 => 
                           n5633, ZN => n5642);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n5708, B1 => 
                           REGISTERS_12_2_port, B2 => n5721, ZN => n5640);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_14_2_port, A2 => n5716, B1 => 
                           REGISTERS_11_2_port, B2 => n5710, ZN => n5639);
   U2789 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n5711, B1 => 
                           REGISTERS_8_2_port, B2 => n5720, ZN => n5638);
   U2790 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n5672, B1 => 
                           REGISTERS_13_2_port, B2 => n5718, ZN => n5637);
   U2791 : NAND4_X1 port map( A1 => n5640, A2 => n5639, A3 => n5638, A4 => 
                           n5637, ZN => n5641);
   U2792 : AOI22_X1 port map( A1 => n5729, A2 => n5642, B1 => n5727, B2 => 
                           n5641, ZN => n5643);
   U2793 : OAI21_X1 port map( B1 => n5732, B2 => n5644, A => n5643, ZN => N387)
                           ;
   U2794 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n5645, B1 => 
                           REGISTERS_17_1_port, B2 => n5695, ZN => n5652);
   U2795 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n5693, B1 => 
                           REGISTERS_20_1_port, B2 => n5683, ZN => n5651);
   U2796 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n5686, B1 => 
                           REGISTERS_27_1_port, B2 => n5646, ZN => n5650);
   U2797 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n5648, B1 => 
                           REGISTERS_16_1_port, B2 => n5647, ZN => n5649);
   U2798 : NAND4_X1 port map( A1 => n5652, A2 => n5651, A3 => n5650, A4 => 
                           n5649, ZN => n5663);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n5654, B1 => 
                           REGISTERS_24_1_port, B2 => n5653, ZN => n5661);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_30_1_port, A2 => n5696, B1 => 
                           REGISTERS_22_1_port, B2 => n5681, ZN => n5660);
   U2801 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n5655, B1 => 
                           REGISTERS_31_1_port, B2 => n5698, ZN => n5659);
   U2802 : AOI22_X1 port map( A1 => REGISTERS_26_1_port, A2 => n5657, B1 => 
                           REGISTERS_23_1_port, B2 => n5656, ZN => n5658);
   U2803 : NAND4_X1 port map( A1 => n5661, A2 => n5660, A3 => n5659, A4 => 
                           n5658, ZN => n5662);
   U2804 : NOR2_X1 port map( A1 => n5663, A2 => n5662, ZN => n5680);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n5718, B1 => 
                           REGISTERS_2_1_port, B2 => n5707, ZN => n5667);
   U2806 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n5671, B1 => 
                           REGISTERS_4_1_port, B2 => n5721, ZN => n5666);
   U2807 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n5720, B1 => 
                           REGISTERS_3_1_port, B2 => n5717, ZN => n5665);
   U2808 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n5716, B1 => 
                           REGISTERS_1_1_port, B2 => n5708, ZN => n5664);
   U2809 : NAND4_X1 port map( A1 => n5667, A2 => n5666, A3 => n5665, A4 => 
                           n5664, ZN => n5678);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n5669, B1 => 
                           REGISTERS_8_1_port, B2 => n5668, ZN => n5676);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n5671, B1 => 
                           REGISTERS_14_1_port, B2 => n5670, ZN => n5675);
   U2812 : AOI22_X1 port map( A1 => REGISTERS_10_1_port, A2 => n5672, B1 => 
                           REGISTERS_11_1_port, B2 => n5710, ZN => n5674);
   U2813 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n5718, B1 => 
                           REGISTERS_9_1_port, B2 => n5708, ZN => n5673);
   U2814 : NAND4_X1 port map( A1 => n5676, A2 => n5675, A3 => n5674, A4 => 
                           n5673, ZN => n5677);
   U2815 : AOI22_X1 port map( A1 => n5729, A2 => n5678, B1 => n5727, B2 => 
                           n5677, ZN => n5679);
   U2816 : OAI21_X1 port map( B1 => n5732, B2 => n5680, A => n5679, ZN => N386)
                           ;
   U2817 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n5682, B1 => 
                           REGISTERS_22_0_port, B2 => n5681, ZN => n5692);
   U2818 : AOI22_X1 port map( A1 => REGISTERS_18_0_port, A2 => n5684, B1 => 
                           REGISTERS_20_0_port, B2 => n5683, ZN => n5691);
   U2819 : AOI22_X1 port map( A1 => REGISTERS_19_0_port, A2 => n5686, B1 => 
                           REGISTERS_29_0_port, B2 => n5685, ZN => n5690);
   U2820 : AOI22_X1 port map( A1 => REGISTERS_26_0_port, A2 => n5688, B1 => 
                           REGISTERS_21_0_port, B2 => n5687, ZN => n5689);
   U2821 : NAND4_X1 port map( A1 => n5692, A2 => n5691, A3 => n5690, A4 => 
                           n5689, ZN => n5706);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n5694, B1 => 
                           REGISTERS_25_0_port, B2 => n5693, ZN => n5704);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_30_0_port, A2 => n5696, B1 => 
                           REGISTERS_17_0_port, B2 => n5695, ZN => n5703);
   U2824 : AOI22_X1 port map( A1 => REGISTERS_31_0_port, A2 => n5698, B1 => 
                           REGISTERS_23_0_port, B2 => n5697, ZN => n5702);
   U2825 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n5700, B1 => 
                           REGISTERS_24_0_port, B2 => n5699, ZN => n5701);
   U2826 : NAND4_X1 port map( A1 => n5704, A2 => n5703, A3 => n5702, A4 => 
                           n5701, ZN => n5705);
   U2827 : NOR2_X1 port map( A1 => n5706, A2 => n5705, ZN => n5731);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n5707, B1 => 
                           REGISTERS_0_0_port, B2 => n5720, ZN => n5715);
   U2829 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n5718, B1 => 
                           REGISTERS_4_0_port, B2 => n5721, ZN => n5714);
   U2830 : AOI22_X1 port map( A1 => REGISTERS_6_0_port, A2 => n5709, B1 => 
                           REGISTERS_1_0_port, B2 => n5708, ZN => n5713);
   U2831 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n5711, B1 => 
                           REGISTERS_3_0_port, B2 => n5710, ZN => n5712);
   U2832 : NAND4_X1 port map( A1 => n5715, A2 => n5714, A3 => n5713, A4 => 
                           n5712, ZN => n5728);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n5717, B1 => 
                           REGISTERS_14_0_port, B2 => n5716, ZN => n5725);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n5718, B1 => 
                           REGISTERS_10_0_port, B2 => n5707, ZN => n5724);
   U2835 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n5720, B1 => 
                           REGISTERS_9_0_port, B2 => n5719, ZN => n5723);
   U2836 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n5721, B1 => 
                           REGISTERS_15_0_port, B2 => n5671, ZN => n5722);
   U2837 : NAND4_X1 port map( A1 => n5725, A2 => n5724, A3 => n5723, A4 => 
                           n5722, ZN => n5726);
   U2838 : AOI22_X1 port map( A1 => n5729, A2 => n5728, B1 => n5727, B2 => 
                           n5726, ZN => n5730);
   U2839 : OAI21_X1 port map( B1 => n5732, B2 => n5731, A => n5730, ZN => N385)
                           ;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, n778, IRAM_ADDRESS_29_port, n779, 
      IRAM_ADDRESS_27_port, n780, IRAM_ADDRESS_25_port, n781, 
      IRAM_ADDRESS_23_port, n782, IRAM_ADDRESS_21_port, n783, 
      IRAM_ADDRESS_19_port, n784, IRAM_ADDRESS_17_port, n785, 
      IRAM_ADDRESS_15_port, n786, IRAM_ADDRESS_13_port, n787, 
      IRAM_ADDRESS_11_port, n788, IRAM_ADDRESS_9_port, n789, 
      IRAM_ADDRESS_7_port, n790, IRAM_ADDRESS_5_port, n791, n792, n793, 
      DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      curr_instruction_to_cu_i_31_port, curr_instruction_to_cu_i_30_port, 
      curr_instruction_to_cu_i_29_port, curr_instruction_to_cu_i_28_port, 
      curr_instruction_to_cu_i_27_port, curr_instruction_to_cu_i_26_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_5_port, curr_instruction_to_cu_i_4_port, 
      curr_instruction_to_cu_i_3_port, curr_instruction_to_cu_i_2_port, 
      curr_instruction_to_cu_i_1_port, curr_instruction_to_cu_i_0_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n153, cu_i_n152, 
      cu_i_n151, cu_i_n135, cu_i_n133, cu_i_n132, cu_i_n128, cu_i_n127, cu_i_n4
      , cu_i_n3, cu_i_n2, cu_i_n210, cu_i_n209, cu_i_n145, cu_i_cw1_i_4_port, 
      cu_i_cw1_i_7_port, cu_i_cw1_i_8_port, cu_i_cw3_5_port, cu_i_cw3_6_port, 
      cu_i_cw2_4_port, cu_i_cw2_5_port, cu_i_cw2_6_port, cu_i_cw2_7_port, 
      cu_i_cw2_8_port, cu_i_cw1_0_port, cu_i_cw1_1_port, cu_i_cw1_2_port, 
      cu_i_cw1_3_port, cu_i_cw1_4_port, cu_i_cw1_5_port, cu_i_cw1_6_port, 
      cu_i_cw1_7_port, cu_i_cw1_8_port, cu_i_cw1_10_port, cu_i_cw1_11_port, 
      cu_i_cw1_12_port, cu_i_cw1_13_port, cu_i_cw1_14_port, cu_i_N279, 
      cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, 
      cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, 
      cu_i_cmd_word_4_port, cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, 
      cu_i_cmd_word_8_port, cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_immediate_i_26_port, 
      datapath_i_val_immediate_i_27_port, datapath_i_val_immediate_i_28_port, 
      datapath_i_val_immediate_i_29_port, datapath_i_val_immediate_i_30_port, 
      datapath_i_val_immediate_i_31_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n81, 
      datapath_i_decode_stage_dp_n80, datapath_i_decode_stage_dp_n79, 
      datapath_i_decode_stage_dp_n78, datapath_i_decode_stage_dp_n77, 
      datapath_i_decode_stage_dp_n44, datapath_i_decode_stage_dp_n43, 
      datapath_i_decode_stage_dp_n42, datapath_i_decode_stage_dp_n41, 
      datapath_i_decode_stage_dp_n40, datapath_i_decode_stage_dp_n39, 
      datapath_i_decode_stage_dp_n38, datapath_i_decode_stage_dp_n37, 
      datapath_i_decode_stage_dp_n36, datapath_i_decode_stage_dp_n35, 
      datapath_i_decode_stage_dp_n34, datapath_i_decode_stage_dp_n33, 
      datapath_i_decode_stage_dp_n32, datapath_i_decode_stage_dp_n31, 
      datapath_i_decode_stage_dp_n30, datapath_i_decode_stage_dp_n29, 
      datapath_i_decode_stage_dp_n28, datapath_i_decode_stage_dp_n27, 
      datapath_i_decode_stage_dp_n26, datapath_i_decode_stage_dp_n25, 
      datapath_i_decode_stage_dp_n24, datapath_i_decode_stage_dp_n23, 
      datapath_i_decode_stage_dp_n22, datapath_i_decode_stage_dp_n21, 
      datapath_i_decode_stage_dp_n20, datapath_i_decode_stage_dp_n19, 
      datapath_i_decode_stage_dp_n18, datapath_i_decode_stage_dp_n17, 
      datapath_i_decode_stage_dp_n16, datapath_i_decode_stage_dp_n15, 
      datapath_i_decode_stage_dp_n14, datapath_i_decode_stage_dp_n13, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_3_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n301, n302, n304, n305, n306,
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, DRAM_ENABLE_port, n326, 
      IRAM_ADDRESS_2_port, n328, IRAM_ADDRESS_3_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_26_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_20_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_14_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_8_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_4_port, IRAM_ENABLE_port, n345, n346, n347, n348, n349, n350
      , n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
      n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
      n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, 
      n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, 
      n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, 
      n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
      n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n_1592, n_1593, n_1594, n_1595,
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => cu_i_n151, QN => n_1592);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => cu_i_n2, QN => n769);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => cu_i_n4, QN => n771);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => cu_i_n152, QN => n721);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => cu_i_n153, QN => n725);
   cu_i_stall_reg : DFFR_X1 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n719, QN => n759);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n43, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n44, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1593, mul_exeception => 
                           n_1594, FUNC(0) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_3_port, 
                           FUNC(1) => datapath_i_execute_stage_dp_n7, FUNC(2) 
                           => datapath_i_execute_stage_dp_alu_op_type_i_1_port,
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1595, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n773, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n773, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n773, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n773, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n773, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n773, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n773, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n773, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n773, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n773, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n773, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n773, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n361, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n361, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n361, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n361, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n361, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n773, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n773, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n773, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n773, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n773, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n773, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n773, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n773, Z =>
                           DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n773, Z =>
                           DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n773, Z =>
                           DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n773, Z =>
                           DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n773, Z =>
                           DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n773, Z =>
                           DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n777, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n777, Z => 
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n777, Z => 
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n777, Z => 
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n777, Z => 
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n777, Z => 
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n777, Z => 
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n777, Z => 
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n777, Z => 
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n777, Z => 
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n777, Z => 
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n777, Z => 
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => n777, Z => 
                           DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => n777, Z => 
                           DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => n777, Z => 
                           DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => n777, Z => 
                           DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => n777, Z => 
                           DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => n777, Z => 
                           DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => n777, Z => 
                           DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => n777, Z => 
                           DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1596);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n301, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n301, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n301, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n301, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n301, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n772, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n301, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n776, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n775, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n774, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n775, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n774, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n775, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n774, D => datapath_i_n18, Q
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n774, D => datapath_i_n17, Q
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n775, D => datapath_i_n16, Q
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n774, D => datapath_i_n15, Q
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n775, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n774, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n775, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n774, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n775, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n774, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n776, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n776, D => 
                           curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n776, D => 
                           curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n776, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n776, D => 
                           curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n775, D => datapath_i_n12, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n11, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n10, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n776, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n133, CK => CLK, RN =>
                           RST, Q => cu_i_cw3_6_port, QN => n_1597);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n132, CK => CLK, RN =>
                           RST, Q => cu_i_cw3_5_port, QN => n768);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1598);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1599);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n128, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1600);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n_1601);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_4_port, QN => n_1602);
   cu_i_e_reg_D_I_14_Q_reg : DFFR_X1 port map( D => cu_i_n135, CK => CLK, RN =>
                           RST, Q => cu_i_cw1_14_port, QN => n_1603);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n772, CK => CLK, RN => RST,
                           Q => cu_i_cw1_13_port, QN => n_1604);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1605)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1606)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1607)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1608);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1609);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n302, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1610);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1611);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_n135, CK => CLK, RN => 
                           RST, Q => cu_i_cw1_4_port, QN => n_1612);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1613);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1614);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1615);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1616);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1617);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1618);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1619);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1620);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1621);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1622);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1623);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1624);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1625);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1626);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1627);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1628);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1629);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1630);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1631);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1632);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1633);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1634);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1635);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1636);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1637);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1638);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1639);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1640);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1641);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1642);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1643);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1644);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1645);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1646);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1647);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1648)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1649)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1650)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1651)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1652)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1653)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1654)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1655)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1656)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1657)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1658)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1659)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1660)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1661)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1662)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1663)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1664)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1665)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1666)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1667)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1668)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1669)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1670);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1671);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1672);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1673);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1674);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1675);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1676);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1677);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1678);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1679);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1680);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1681);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1682);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1683);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1684);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1685);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1686);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1687);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1688);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1689);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1690);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1691);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1692);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1693);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1694);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1695);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1696);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1697);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1698);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1699);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1700);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1701);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1702);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1703);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1704);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1705);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1706);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1707);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1708);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1709);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1710);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1711);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1712);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1713);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1714);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1715);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1716);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1717);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1718);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1719);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1720);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1721);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1722);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1723);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1724);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1725);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1726);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1727);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1728);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1729);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1730);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1731);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1732);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1733);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1734);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1735);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1736);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1737);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1738);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1739);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1740);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1741);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1742);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1743);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => n717, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1744, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1745, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1746, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1747, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1748, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1749, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1750, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1751, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1752, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1753, QN => n745);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1754, QN => n744);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1755, QN => n743);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1756, QN => n742);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1757, QN => n741);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1758, QN => n740);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1759, QN => n739);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1760, QN => n738);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1761, QN => n737);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1762, QN => n736);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1763, QN => n735);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1764, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1765, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1766, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1767, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1768, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1769, QN => n750);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1770, QN => n749);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1771, QN => n748);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1772, QN => n747);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1773, QN => n746);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1774, QN => n752);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1775, QN => n751);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1776);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1777);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1778);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1779);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1780);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1781);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1782);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1783);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1784);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1785);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1786);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1787);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1788);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1789);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1790);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1791);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1792);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1793);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1794);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1795);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1796);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1797);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1798);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1799);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1800);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1801);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1802);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1803);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1804);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1805);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1806);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1807);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1808);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n776, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1809);
   datapath_i_decode_stage_dp_reg_immediate_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_31_port, QN 
                           => n_1810);
   datapath_i_decode_stage_dp_reg_immediate_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_30_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_30_port, QN 
                           => n_1811);
   datapath_i_decode_stage_dp_reg_immediate_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_29_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_29_port, QN 
                           => n_1812);
   datapath_i_decode_stage_dp_reg_immediate_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_28_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_28_port, QN 
                           => n_1813);
   datapath_i_decode_stage_dp_reg_immediate_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_27_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_27_port, QN 
                           => n_1814);
   datapath_i_decode_stage_dp_reg_immediate_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_26_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_26_port, QN 
                           => n_1815);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_25_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1816);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1817);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1818);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1819);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1820);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1821);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1822);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1823);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1824);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1825);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1826);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1827);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1828);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1829);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1830);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1831);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1832);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1833);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1834);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1835);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1836);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1837);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1838);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1839);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1840);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1841);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n_1842);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n_1843);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n_1844);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n_1845);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n_1846);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n_1847);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n_1848);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1849);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1850);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1851);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1852);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1853);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1854);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1855);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1856);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1857);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1858);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1859);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1860);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1861);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1862);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1863);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1864);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1865);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1866);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1867);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1868);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1869);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1870);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1871);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1872);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1873);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1874);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1875);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1876);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1877);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1878);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1879);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1880);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1881);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1882);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1883);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1884);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1885);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1886);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1887);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1888);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1889);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1890);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1891);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1892);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1893);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1894);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1895);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1896);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1897);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1898);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1899);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1900);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1901);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1902);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1903);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1904);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1905);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1906);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1907);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1908);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1909);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1910);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1911);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1912);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1913);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1914);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1915);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n77, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1916);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1917);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n79, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1918);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n80, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1919);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n81, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1920);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n716);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n724);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_29_port, QN => 
                           n722);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n715);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n723);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n706);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1921);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1922);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1923);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1924);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1925);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1926);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1927);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n720);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1928);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1929);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1930);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n760);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1931);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1932);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1933);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1934);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1935);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1936);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1937);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n728);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n_1938);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n_1939);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n718);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n726);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n770);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1940
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1941
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1942
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1943
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1944
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1945
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1946
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1947
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1948
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1949
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1950
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1951
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1952
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1953
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1954
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1955
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1956
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1957
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1958
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1959
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1960
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1961
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1962)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1963)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1964)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1965)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1966)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1967)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1968)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1969)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1970)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1971)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1972);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => n778, QN => n_1973);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n767);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => n779, QN => n_1974);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n766);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => n780, QN => n_1975);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n765);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => n781, QN => n_1976);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n764);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => n782, QN => n_1977);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n763);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => n783, QN => n_1978);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n762);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => n784, QN => n_1979);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n761);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => n785, QN => n_1980);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n758);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => n786, QN => n_1981);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n757);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => n787, QN => n_1982);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n756);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => n788, QN => n_1983);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n755
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => n789, QN => n_1984);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n754
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => n790, QN => n_1985);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n753
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => n791, QN => n_1986);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => n792, QN => n_1987);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => n_1988, QN => n326);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1989);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1990);
   U308 : AND2_X1 port map( A1 => n306, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   U309 : AND2_X1 port map( A1 => n305, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U310 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U311 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U312 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U313 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U314 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U315 : AND2_X1 port map( A1 => n323, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U316 : AND2_X1 port map( A1 => n322, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U317 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U318 : AND2_X1 port map( A1 => n321, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U319 : AND2_X1 port map( A1 => n320, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U320 : AND2_X1 port map( A1 => n319, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U321 : AND2_X1 port map( A1 => n318, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U322 : AND2_X1 port map( A1 => n317, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U323 : AND2_X1 port map( A1 => n316, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U324 : AND2_X1 port map( A1 => n315, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U325 : AND2_X1 port map( A1 => n314, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U326 : AND2_X1 port map( A1 => n313, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U327 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U328 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U329 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U330 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U331 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U332 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U333 : AND2_X1 port map( A1 => n312, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U334 : AND2_X1 port map( A1 => n311, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U335 : AND2_X1 port map( A1 => n310, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U336 : AND2_X1 port map( A1 => n309, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U337 : AND2_X1 port map( A1 => n308, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U338 : AND2_X1 port map( A1 => n307, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U339 : AND2_X1 port map( A1 => n304, A2 => DRAM_READY, ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => cu_i_n3, QN => n_1991);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1992);
   U591 : BUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n777);
   U592 : CLKBUF_X1 port map( A => DRAM_DATA(0), Z => n304);
   U593 : CLKBUF_X1 port map( A => DRAM_DATA(8), Z => n305);
   U594 : CLKBUF_X1 port map( A => DRAM_DATA(9), Z => n306);
   U595 : CLKBUF_X1 port map( A => DRAM_DATA(10), Z => n307);
   U596 : CLKBUF_X1 port map( A => DRAM_DATA(11), Z => n308);
   U597 : CLKBUF_X1 port map( A => DRAM_DATA(12), Z => n309);
   U598 : CLKBUF_X1 port map( A => DRAM_DATA(13), Z => n310);
   U599 : CLKBUF_X1 port map( A => DRAM_DATA(14), Z => n311);
   U600 : CLKBUF_X1 port map( A => DRAM_DATA(15), Z => n312);
   U601 : CLKBUF_X1 port map( A => DRAM_DATA(21), Z => n313);
   U602 : CLKBUF_X1 port map( A => DRAM_DATA(22), Z => n314);
   U603 : CLKBUF_X1 port map( A => DRAM_DATA(23), Z => n315);
   U604 : CLKBUF_X1 port map( A => DRAM_DATA(24), Z => n316);
   U605 : CLKBUF_X1 port map( A => DRAM_DATA(25), Z => n317);
   U606 : CLKBUF_X1 port map( A => DRAM_DATA(26), Z => n318);
   U607 : CLKBUF_X1 port map( A => DRAM_DATA(27), Z => n319);
   U608 : CLKBUF_X1 port map( A => DRAM_DATA(28), Z => n320);
   U609 : CLKBUF_X1 port map( A => DRAM_DATA(29), Z => n321);
   U610 : CLKBUF_X1 port map( A => DRAM_DATA(30), Z => n322);
   U611 : CLKBUF_X1 port map( A => DRAM_DATA(31), Z => n323);
   U612 : INV_X1 port map( A => n362, ZN => n324);
   U613 : INV_X2 port map( A => n324, ZN => DRAM_ENABLE_port);
   U614 : INV_X2 port map( A => n375, ZN => n597);
   U615 : NAND2_X2 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n445, ZN => n705);
   U616 : INV_X2 port map( A => n445, ZN => n702);
   U617 : INV_X2 port map( A => n759, ZN => n669);
   U618 : INV_X2 port map( A => n326, ZN => IRAM_ADDRESS_2_port);
   U619 : OAI21_X2 port map( B1 => n732, B2 => n705, A => n679, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U620 : OAI21_X2 port map( B1 => n731, B2 => n705, A => n447, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U621 : OAI21_X2 port map( B1 => n738, B2 => n705, A => n446, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U622 : OAI21_X2 port map( B1 => n742, B2 => n705, A => n684, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U623 : OAI21_X2 port map( B1 => n739, B2 => n705, A => n682, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U624 : OAI21_X2 port map( B1 => n735, B2 => n705, A => n452, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U625 : OAI21_X2 port map( B1 => n748, B2 => n705, A => n450, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U626 : OAI21_X2 port map( B1 => n733, B2 => n705, A => n448, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U627 : OAI21_X2 port map( B1 => n710, B2 => n705, A => n691, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U628 : OAI21_X2 port map( B1 => n750, B2 => n705, A => n449, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);
   U629 : OAI21_X2 port map( B1 => n741, B2 => n705, A => n453, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U630 : OAI21_X2 port map( B1 => n734, B2 => n705, A => n451, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U631 : CLKBUF_X1 port map( A => IRAM_ADDRESS_31_port, Z => n328);
   U632 : CLKBUF_X1 port map( A => n792, Z => IRAM_ADDRESS_3_port);
   U633 : CLKBUF_X1 port map( A => n778, Z => IRAM_ADDRESS_30_port);
   U634 : CLKBUF_X1 port map( A => n779, Z => IRAM_ADDRESS_28_port);
   U635 : CLKBUF_X1 port map( A => n780, Z => IRAM_ADDRESS_26_port);
   U636 : CLKBUF_X1 port map( A => n781, Z => IRAM_ADDRESS_24_port);
   U637 : CLKBUF_X1 port map( A => n782, Z => IRAM_ADDRESS_22_port);
   U638 : CLKBUF_X1 port map( A => n783, Z => IRAM_ADDRESS_20_port);
   U639 : CLKBUF_X1 port map( A => n784, Z => IRAM_ADDRESS_18_port);
   U640 : CLKBUF_X1 port map( A => n785, Z => IRAM_ADDRESS_16_port);
   U641 : CLKBUF_X1 port map( A => n786, Z => IRAM_ADDRESS_14_port);
   U642 : CLKBUF_X1 port map( A => n787, Z => IRAM_ADDRESS_12_port);
   U643 : CLKBUF_X1 port map( A => n788, Z => IRAM_ADDRESS_10_port);
   U644 : CLKBUF_X1 port map( A => n789, Z => IRAM_ADDRESS_8_port);
   U645 : CLKBUF_X1 port map( A => n790, Z => IRAM_ADDRESS_6_port);
   U646 : CLKBUF_X1 port map( A => n791, Z => IRAM_ADDRESS_4_port);
   U647 : CLKBUF_X1 port map( A => n793, Z => IRAM_ENABLE_port);
   U648 : AOI21_X1 port map( B1 => n616, B2 => n615, A => cu_i_cw3_6_port, ZN 
                           => n617);
   U649 : CLKBUF_X1 port map( A => n637, Z => n652);
   U650 : OAI21_X1 port map( B1 => n490, B2 => n489, A => n768, ZN => 
                           write_rf_i);
   U651 : NOR2_X1 port map( A1 => n509, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n423);
   U652 : NOR2_X1 port map( A1 => n656, A2 => n443, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U653 : OAI21_X1 port map( B1 => cu_i_n2, B2 => cu_i_n4, A => cu_i_n151, ZN 
                           => n489);
   U654 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           curr_instruction_to_cu_i_28_port, A3 => n459, A4 => 
                           n352, ZN => n502);
   U655 : NOR2_X1 port map( A1 => cu_i_n3, A2 => n725, ZN => n408);
   U656 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n727, ZN => n513);
   U657 : CLKBUF_X1 port map( A => n513, Z => n458);
   U658 : AOI21_X1 port map( B1 => n373, B2 => n410, A => n495, ZN => n613);
   U659 : NOR3_X1 port map( A1 => n728, A2 => n718, A3 => n355, ZN => n410);
   U660 : OR3_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => 
                           curr_instruction_to_cu_i_29_port, A3 => n497, ZN => 
                           n611);
   U661 : NOR2_X1 port map( A1 => n609, A2 => n504, ZN => n411);
   U662 : NOR3_X1 port map( A1 => n716, A2 => n706, A3 => n497, ZN => 
                           cu_i_cmd_word_4_port);
   U663 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n716
                           , A3 => n724, ZN => n370);
   U664 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => n723
                           , ZN => n474);
   U665 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_29_port, A2 => n370,
                           A3 => n474, ZN => n351);
   U666 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => n722,
                           ZN => n491);
   U667 : NAND2_X1 port map( A1 => n706, A2 => n723, ZN => n459);
   U668 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           curr_instruction_to_cu_i_28_port, A3 => n459, ZN => 
                           n347);
   U669 : NAND2_X1 port map( A1 => n716, A2 => n722, ZN => n352);
   U670 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => n715,
                           A3 => n724, A4 => n352, ZN => n468);
   U671 : NOR2_X1 port map( A1 => n370, A2 => n722, ZN => n480);
   U672 : INV_X1 port map( A => n480, ZN => n345);
   U673 : NAND3_X1 port map( A1 => n724, A2 => n715, A3 => 
                           curr_instruction_to_cu_i_27_port, ZN => n349);
   U674 : INV_X1 port map( A => n349, ZN => n608);
   U675 : OAI221_X1 port map( B1 => n480, B2 => n608, C1 => n480, C2 => n491, A
                           => n706, ZN => n464);
   U676 : AND2_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => n491,
                           ZN => n475);
   U677 : OAI211_X1 port map( C1 => curr_instruction_to_cu_i_28_port, C2 => 
                           curr_instruction_to_cu_i_26_port, A => n475, B => 
                           n723, ZN => n485);
   U678 : OAI211_X1 port map( C1 => n345, C2 => n474, A => n464, B => n485, ZN 
                           => n346);
   U679 : AOI211_X1 port map( C1 => n491, C2 => n347, A => n468, B => n346, ZN 
                           => n499);
   U680 : INV_X1 port map( A => n370, ZN => n348);
   U681 : INV_X1 port map( A => n459, ZN => n473);
   U682 : NAND2_X1 port map( A1 => n348, A2 => n473, ZN => n371);
   U683 : NAND2_X1 port map( A1 => n499, A2 => n371, ZN => n407);
   U684 : AOI221_X1 port map( B1 => curr_instruction_to_cu_i_31_port, B2 => 
                           n706, C1 => n716, C2 => 
                           curr_instruction_to_cu_i_29_port, A => n349, ZN => 
                           n350);
   U685 : NOR3_X1 port map( A1 => n351, A2 => n407, A3 => n350, ZN => n505);
   U686 : INV_X1 port map( A => n408, ZN => n609);
   U687 : NOR2_X1 port map( A1 => n505, A2 => n609, ZN => n301);
   U688 : CLKBUF_X1 port map( A => n301, Z => n772);
   U689 : INV_X1 port map( A => n502, ZN => n504);
   U690 : OR2_X1 port map( A1 => n411, A2 => n772, ZN => cu_i_N278);
   U691 : OAI22_X1 port map( A1 => n759, A2 => cu_i_cw3_6_port, B1 => 
                           cu_i_cw2_6_port, B2 => n669, ZN => n353);
   U692 : INV_X1 port map( A => n353, ZN => cu_i_n133);
   U693 : OAI22_X1 port map( A1 => n759, A2 => cu_i_cw3_5_port, B1 => 
                           cu_i_cw2_5_port, B2 => n669, ZN => n354);
   U694 : INV_X1 port map( A => n354, ZN => cu_i_n132);
   U695 : NAND2_X1 port map( A1 => n408, A2 => n608, ZN => n497);
   U696 : AND2_X1 port map( A1 => n722, A2 => cu_i_cmd_word_4_port, ZN => 
                           cu_i_cmd_word_3_port);
   U697 : INV_X1 port map( A => n411, ZN => n495);
   U698 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => 
                           curr_instruction_to_cu_i_3_port, A3 => 
                           curr_instruction_to_cu_i_0_port, A4 => 
                           curr_instruction_to_cu_i_4_port, ZN => n355);
   U699 : OAI222_X1 port map( A1 => n611, A2 => n706, B1 => n495, B2 => n410, 
                           C1 => n609, C2 => n499, ZN => n302);
   U700 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n302, ZN => 
                           cu_i_cmd_word_1_port);
   U701 : INV_X1 port map( A => n611, ZN => n774);
   U702 : INV_X1 port map( A => n611, ZN => n775);
   U703 : OAI22_X1 port map( A1 => n759, A2 => cu_i_cmd_word_3_port, B1 => 
                           cu_i_cw2_7_port, B2 => n669, ZN => n365);
   U704 : INV_X1 port map( A => n365, ZN => DRAM_READNOTWRITE);
   U705 : NOR2_X1 port map( A1 => cu_i_n2, A2 => cu_i_n4, ZN => n356);
   U706 : NAND3_X1 port map( A1 => n356, A2 => cu_i_n151, A3 => cu_i_n152, ZN 
                           => cu_i_n145);
   U707 : INV_X1 port map( A => n611, ZN => n776);
   U708 : NAND2_X1 port map( A1 => n489, A2 => cu_i_n145, ZN => n373);
   U709 : INV_X1 port map( A => n613, ZN => n612);
   U710 : AOI221_X1 port map( B1 => n612, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n613, C2 => 
                           curr_instruction_to_cu_i_15_port, A => n776, ZN => 
                           n357);
   U711 : INV_X1 port map( A => n357, ZN => datapath_i_decode_stage_dp_n77);
   U712 : AOI221_X1 port map( B1 => n612, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n613, C2 => 
                           curr_instruction_to_cu_i_14_port, A => n776, ZN => 
                           n358);
   U713 : INV_X1 port map( A => n358, ZN => datapath_i_decode_stage_dp_n78);
   U714 : AOI221_X1 port map( B1 => n612, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n613, C2 => 
                           curr_instruction_to_cu_i_11_port, A => n776, ZN => 
                           n359);
   U715 : INV_X1 port map( A => n359, ZN => datapath_i_decode_stage_dp_n81);
   U716 : AOI221_X1 port map( B1 => n612, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n613, C2 => 
                           curr_instruction_to_cu_i_12_port, A => n776, ZN => 
                           n360);
   U717 : INV_X1 port map( A => n360, ZN => datapath_i_decode_stage_dp_n80);
   U718 : OAI22_X1 port map( A1 => n759, A2 => cu_i_cmd_word_4_port, B1 => 
                           cu_i_cw2_8_port, B2 => n669, ZN => n361);
   U719 : INV_X1 port map( A => n361, ZN => n362);
   U720 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n773);
   U721 : INV_X1 port map( A => n727, ZN => n509);
   U722 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_3_port, ZN => n363
                           );
   U723 : OAI21_X1 port map( B1 => n458, B2 => n747, A => n363, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U724 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_2_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_2_port, ZN => n364
                           );
   U725 : OAI21_X1 port map( B1 => n458, B2 => n746, A => n364, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U726 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n365, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U727 : CLKBUF_X1 port map( A => n423, Z => n511);
   U728 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_7_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_7_port, ZN => n366
                           );
   U729 : OAI21_X1 port map( B1 => n513, B2 => n730, A => n366, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U730 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_5_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_5_port, ZN => n367
                           );
   U731 : OAI21_X1 port map( B1 => n513, B2 => n749, A => n367, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U732 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_4_port, ZN => n368
                           );
   U733 : OAI21_X1 port map( B1 => n458, B2 => n748, A => n368, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U734 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_6_port, ZN => n369
                           );
   U735 : OAI21_X1 port map( B1 => n513, B2 => n750, A => n369, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U736 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_29_port, A2 => n370,
                           A3 => n609, A4 => n474, ZN => cu_i_cmd_word_7_port);
   U737 : OR2_X1 port map( A1 => n609, A2 => n371, ZN => n372);
   U738 : OAI21_X1 port map( B1 => n372, B2 => curr_instruction_to_cu_i_29_port
                           , A => n611, ZN => cu_i_cmd_word_6_port);
   U739 : OR2_X1 port map( A1 => cu_i_cmd_word_7_port, A2 => 
                           cu_i_cmd_word_6_port, ZN => cu_i_n135);
   U740 : NAND2_X1 port map( A1 => n502, A2 => n410, ZN => n477);
   U741 : AOI22_X1 port map( A1 => n408, A2 => n477, B1 => n411, B2 => n373, ZN
                           => n374);
   U742 : NAND2_X1 port map( A1 => cu_i_n3, A2 => n725, ZN => n506);
   U743 : AOI21_X1 port map( B1 => n374, B2 => n506, A => n669, ZN => n793);
   U744 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN 
                           => n376);
   U745 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN 
                           => n379);
   U746 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_2_port, ZN =>
                           n519);
   U747 : NOR2_X1 port map( A1 => n379, A2 => n519, ZN => n526);
   U748 : NAND2_X1 port map( A1 => n526, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n525);
   U749 : AOI221_X1 port map( B1 => cu_i_cw2_4_port, B2 => n759, C1 => 
                           cu_i_n135, C2 => n669, A => n717, ZN => n375);
   U750 : INV_X1 port map( A => n597, ZN => n599);
   U751 : NOR2_X1 port map( A1 => n376, A2 => n525, ZN => n532);
   U752 : AOI211_X1 port map( C1 => n376, C2 => n525, A => n599, B => n532, ZN 
                           => n378);
   U753 : NAND2_X1 port map( A1 => n793, A2 => IRAM_ADDRESS_2_port, ZN => n514)
                           ;
   U754 : INV_X1 port map( A => n514, ZN => n516);
   U755 : AND2_X1 port map( A1 => n516, A2 => n792, ZN => n522);
   U756 : NAND2_X1 port map( A1 => n522, A2 => n791, ZN => n521);
   U757 : NOR2_X1 port map( A1 => n521, A2 => n753, ZN => n528);
   U758 : NAND2_X1 port map( A1 => n528, A2 => n790, ZN => n527);
   U759 : NOR2_X1 port map( A1 => n527, A2 => n754, ZN => n534);
   U760 : AOI211_X1 port map( C1 => n527, C2 => n754, A => n534, B => n597, ZN 
                           => n377);
   U761 : OR2_X1 port map( A1 => n378, A2 => n377, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U762 : AOI211_X1 port map( C1 => n379, C2 => n519, A => n599, B => n526, ZN 
                           => n381);
   U763 : AOI211_X1 port map( C1 => n521, C2 => n753, A => n528, B => n597, ZN 
                           => n380);
   U764 : OR2_X1 port map( A1 => n381, A2 => n380, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U765 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_9_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_9_port, ZN => n382
                           );
   U766 : OAI21_X1 port map( B1 => n513, B2 => n732, A => n382, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U767 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_8_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_8_port, ZN => n383
                           );
   U768 : OAI21_X1 port map( B1 => n513, B2 => n731, A => n383, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U769 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN 
                           => n384);
   U770 : NAND2_X1 port map( A1 => n532, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n531);
   U771 : NOR2_X1 port map( A1 => n384, A2 => n531, ZN => n538);
   U772 : AOI211_X1 port map( C1 => n384, C2 => n531, A => n599, B => n538, ZN 
                           => n386);
   U773 : NAND2_X1 port map( A1 => n534, A2 => n789, ZN => n533);
   U774 : NOR2_X1 port map( A1 => n533, A2 => n755, ZN => n540);
   U775 : AOI211_X1 port map( C1 => n533, C2 => n755, A => n540, B => n597, ZN 
                           => n385);
   U776 : OR2_X1 port map( A1 => n386, A2 => n385, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U777 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_11_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_11_port, ZN => 
                           n387);
   U778 : OAI21_X1 port map( B1 => n513, B2 => n734, A => n387, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U779 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_10_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_10_port, ZN => 
                           n388);
   U780 : OAI21_X1 port map( B1 => n513, B2 => n733, A => n388, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U781 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, ZN
                           => n389);
   U782 : NAND2_X1 port map( A1 => n538, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n537);
   U783 : NOR2_X1 port map( A1 => n389, A2 => n537, ZN => n544);
   U784 : AOI211_X1 port map( C1 => n389, C2 => n537, A => n599, B => n544, ZN 
                           => n391);
   U785 : NAND2_X1 port map( A1 => n540, A2 => n788, ZN => n539);
   U786 : NOR2_X1 port map( A1 => n539, A2 => n756, ZN => n546);
   U787 : AOI211_X1 port map( C1 => n539, C2 => n756, A => n546, B => n597, ZN 
                           => n390);
   U788 : OR2_X1 port map( A1 => n391, A2 => n390, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U789 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_13_port, ZN => 
                           n392);
   U790 : OAI21_X1 port map( B1 => n513, B2 => n736, A => n392, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U791 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_12_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_12_port, ZN => 
                           n393);
   U792 : OAI21_X1 port map( B1 => n513, B2 => n735, A => n393, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U793 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, ZN
                           => n394);
   U794 : NAND2_X1 port map( A1 => n544, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n543);
   U795 : INV_X1 port map( A => n597, ZN => n607);
   U796 : NOR2_X1 port map( A1 => n394, A2 => n543, ZN => n550);
   U797 : AOI211_X1 port map( C1 => n394, C2 => n543, A => n607, B => n550, ZN 
                           => n396);
   U798 : NAND2_X1 port map( A1 => n546, A2 => n787, ZN => n545);
   U799 : NOR2_X1 port map( A1 => n545, A2 => n757, ZN => n552);
   U800 : AOI211_X1 port map( C1 => n545, C2 => n757, A => n552, B => n597, ZN 
                           => n395);
   U801 : OR2_X1 port map( A1 => n396, A2 => n395, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U802 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_15_port, ZN => 
                           n397);
   U803 : OAI21_X1 port map( B1 => n513, B2 => n738, A => n397, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U804 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_14_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_14_port, ZN => 
                           n398);
   U805 : OAI21_X1 port map( B1 => n513, B2 => n737, A => n398, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U806 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, ZN
                           => n399);
   U807 : NAND2_X1 port map( A1 => n550, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n549);
   U808 : NOR2_X1 port map( A1 => n399, A2 => n549, ZN => n556);
   U809 : AOI211_X1 port map( C1 => n399, C2 => n549, A => n599, B => n556, ZN 
                           => n401);
   U810 : NAND2_X1 port map( A1 => n552, A2 => n786, ZN => n551);
   U811 : NOR2_X1 port map( A1 => n551, A2 => n758, ZN => n558);
   U812 : AOI211_X1 port map( C1 => n551, C2 => n758, A => n558, B => n597, ZN 
                           => n400);
   U813 : OR2_X1 port map( A1 => n401, A2 => n400, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U814 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_17_port, ZN => 
                           n402);
   U815 : OAI21_X1 port map( B1 => n513, B2 => n740, A => n402, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U816 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_16_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_16_port, ZN => 
                           n403);
   U817 : OAI21_X1 port map( B1 => n513, B2 => n739, A => n403, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U818 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, ZN
                           => n404);
   U819 : NAND2_X1 port map( A1 => n556, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n555);
   U820 : NOR2_X1 port map( A1 => n404, A2 => n555, ZN => n562);
   U821 : AOI211_X1 port map( C1 => n404, C2 => n555, A => n607, B => n562, ZN 
                           => n406);
   U822 : NAND2_X1 port map( A1 => n558, A2 => n785, ZN => n557);
   U823 : NOR2_X1 port map( A1 => n557, A2 => n761, ZN => n564);
   U824 : AOI211_X1 port map( C1 => n557, C2 => n761, A => n564, B => n597, ZN 
                           => n405);
   U825 : OR2_X1 port map( A1 => n406, A2 => n405, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U826 : AOI211_X1 port map( C1 => n408, C2 => n407, A => cu_i_cmd_word_7_port
                           , B => cu_i_cmd_word_4_port, ZN => n409);
   U827 : NAND2_X1 port map( A1 => n409, A2 => n612, ZN => enable_rf_i);
   U828 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n490);
   U829 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U830 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_19_port, ZN => 
                           n412);
   U831 : OAI21_X1 port map( B1 => n513, B2 => n742, A => n412, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U832 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_18_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_18_port, ZN => 
                           n413);
   U833 : OAI21_X1 port map( B1 => n513, B2 => n741, A => n413, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U834 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, ZN
                           => n414);
   U835 : NAND2_X1 port map( A1 => n562, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n561);
   U836 : NOR2_X1 port map( A1 => n414, A2 => n561, ZN => n568);
   U837 : AOI211_X1 port map( C1 => n414, C2 => n561, A => n607, B => n568, ZN 
                           => n416);
   U838 : NAND2_X1 port map( A1 => n564, A2 => n784, ZN => n563);
   U839 : NOR2_X1 port map( A1 => n563, A2 => n762, ZN => n570);
   U840 : AOI211_X1 port map( C1 => n563, C2 => n762, A => n570, B => n597, ZN 
                           => n415);
   U841 : OR2_X1 port map( A1 => n416, A2 => n415, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U842 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_21_port, ZN => 
                           n417);
   U843 : OAI21_X1 port map( B1 => n513, B2 => n744, A => n417, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U844 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_20_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_20_port, ZN => 
                           n418);
   U845 : OAI21_X1 port map( B1 => n513, B2 => n743, A => n418, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U846 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, ZN
                           => n419);
   U847 : NAND2_X1 port map( A1 => n568, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n567);
   U848 : NOR2_X1 port map( A1 => n419, A2 => n567, ZN => n574);
   U849 : AOI211_X1 port map( C1 => n419, C2 => n567, A => n607, B => n574, ZN 
                           => n421);
   U850 : NAND2_X1 port map( A1 => n570, A2 => n783, ZN => n569);
   U851 : NOR2_X1 port map( A1 => n569, A2 => n763, ZN => n576);
   U852 : AOI211_X1 port map( C1 => n569, C2 => n763, A => n576, B => n597, ZN 
                           => n420);
   U853 : OR2_X1 port map( A1 => n421, A2 => n420, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U854 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_23_port, ZN => 
                           n422);
   U855 : OAI21_X1 port map( B1 => n513, B2 => n707, A => n422, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U856 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_22_port, B1 => n423, B2 
                           => datapath_i_new_pc_value_decode_22_port, ZN => 
                           n424);
   U857 : OAI21_X1 port map( B1 => n513, B2 => n745, A => n424, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U858 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, ZN
                           => n425);
   U859 : NAND2_X1 port map( A1 => n574, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n573);
   U860 : NOR2_X1 port map( A1 => n425, A2 => n573, ZN => n580);
   U861 : AOI211_X1 port map( C1 => n425, C2 => n573, A => n607, B => n580, ZN 
                           => n427);
   U862 : NAND2_X1 port map( A1 => n576, A2 => n782, ZN => n575);
   U863 : NOR2_X1 port map( A1 => n575, A2 => n764, ZN => n582);
   U864 : AOI211_X1 port map( C1 => n575, C2 => n764, A => n582, B => n597, ZN 
                           => n426);
   U865 : OR2_X1 port map( A1 => n427, A2 => n426, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U866 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_25_port, ZN => 
                           n428);
   U867 : OAI21_X1 port map( B1 => n513, B2 => n709, A => n428, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U868 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_24_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_24_port, ZN => 
                           n429);
   U869 : OAI21_X1 port map( B1 => n513, B2 => n708, A => n429, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U870 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, ZN
                           => n430);
   U871 : NAND2_X1 port map( A1 => n580, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n579);
   U872 : NOR2_X1 port map( A1 => n430, A2 => n579, ZN => n586);
   U873 : AOI211_X1 port map( C1 => n430, C2 => n579, A => n607, B => n586, ZN 
                           => n432);
   U874 : NAND2_X1 port map( A1 => n582, A2 => n781, ZN => n581);
   U875 : NOR2_X1 port map( A1 => n581, A2 => n765, ZN => n588);
   U876 : AOI211_X1 port map( C1 => n581, C2 => n765, A => n588, B => n597, ZN 
                           => n431);
   U877 : OR2_X1 port map( A1 => n432, A2 => n431, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U878 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_27_port, ZN => 
                           n433);
   U879 : OAI21_X1 port map( B1 => n458, B2 => n711, A => n433, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U880 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_26_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_26_port, ZN => 
                           n434);
   U881 : OAI21_X1 port map( B1 => n458, B2 => n710, A => n434, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U882 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, ZN
                           => n435);
   U883 : NAND2_X1 port map( A1 => n586, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n585);
   U884 : NOR2_X1 port map( A1 => n435, A2 => n585, ZN => n592);
   U885 : AOI211_X1 port map( C1 => n435, C2 => n585, A => n607, B => n592, ZN 
                           => n437);
   U886 : NAND2_X1 port map( A1 => n588, A2 => n780, ZN => n587);
   U887 : NOR2_X1 port map( A1 => n587, A2 => n766, ZN => n594);
   U888 : AOI211_X1 port map( C1 => n587, C2 => n766, A => n594, B => n597, ZN 
                           => n436);
   U889 : OR2_X1 port map( A1 => n437, A2 => n436, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U890 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_29_port, ZN => 
                           n438);
   U891 : OAI21_X1 port map( B1 => n458, B2 => n713, A => n438, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U892 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_28_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_28_port, ZN => 
                           n439);
   U893 : OAI21_X1 port map( B1 => n458, B2 => n712, A => n439, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U894 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, ZN
                           => n440);
   U895 : NAND2_X1 port map( A1 => n592, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n591);
   U896 : NOR2_X1 port map( A1 => n440, A2 => n591, ZN => n598);
   U897 : AOI211_X1 port map( C1 => n440, C2 => n591, A => n607, B => n598, ZN 
                           => n442);
   U898 : NAND2_X1 port map( A1 => n594, A2 => n779, ZN => n593);
   U899 : NOR2_X1 port map( A1 => n593, A2 => n767, ZN => n600);
   U900 : AOI211_X1 port map( C1 => n593, C2 => n767, A => n600, B => n597, ZN 
                           => n441);
   U901 : OR2_X1 port map( A1 => n442, A2 => n441, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U902 : AOI22_X1 port map( A1 => n669, A2 => cu_i_cmd_alu_op_type_0_port, B1 
                           => cu_i_cw1_0_port, B2 => n759, ZN => n656);
   U903 : AOI22_X1 port map( A1 => n669, A2 => cu_i_cmd_alu_op_type_1_port, B1 
                           => cu_i_cw1_1_port, B2 => n759, ZN => n658);
   U904 : AOI22_X1 port map( A1 => n669, A2 => cu_i_cmd_alu_op_type_2_port, B1 
                           => cu_i_cw1_2_port, B2 => n759, ZN => n675);
   U905 : AOI22_X1 port map( A1 => n669, A2 => cu_i_cmd_alu_op_type_3_port, B1 
                           => cu_i_cw1_3_port, B2 => n759, ZN => n655);
   U906 : AOI21_X1 port map( B1 => n658, B2 => n675, A => n655, ZN => n443);
   U907 : INV_X1 port map( A => n655, ZN => n674);
   U908 : OAI211_X1 port map( C1 => n656, C2 => n658, A => n674, B => n675, ZN 
                           => n444);
   U909 : INV_X1 port map( A => n444, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_3_port);
   U910 : AOI22_X1 port map( A1 => n669, A2 => n772, B1 => cu_i_cw1_13_port, B2
                           => n759, ZN => n676);
   U911 : CLKBUF_X1 port map( A => n676, Z => n677);
   U912 : MUX2_X1 port map( A => datapath_i_val_immediate_i_0_port, B => 
                           datapath_i_val_b_i_0_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U913 : MUX2_X1 port map( A => datapath_i_val_immediate_i_1_port, B => 
                           datapath_i_val_b_i_1_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U914 : MUX2_X1 port map( A => datapath_i_val_immediate_i_2_port, B => 
                           datapath_i_val_b_i_2_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U915 : MUX2_X1 port map( A => cu_i_cw1_14_port, B => cu_i_n135, S => n669, Z
                           => n445);
   U916 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port, 
                           A2 => n702, ZN => n703);
   U917 : CLKBUF_X1 port map( A => n703, Z => n698);
   U918 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n698, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n702, ZN => n446);
   U919 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 =>
                           n698, B1 => datapath_i_val_a_i_8_port, B2 => n702, 
                           ZN => n447);
   U920 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n698, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n702, ZN => n448);
   U921 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 =>
                           n698, B1 => datapath_i_val_a_i_6_port, B2 => n702, 
                           ZN => n449);
   U922 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 =>
                           n703, B1 => datapath_i_val_a_i_4_port, B2 => n702, 
                           ZN => n450);
   U923 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n698, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n702, ZN => n451);
   U924 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n698, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n702, ZN => n452);
   U925 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n698, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n702, ZN => n453);
   U926 : INV_X1 port map( A => n490, ZN => n616);
   U927 : NAND3_X1 port map( A1 => cu_i_n4, A2 => cu_i_n152, A3 => n616, ZN => 
                           n487);
   U928 : NOR2_X1 port map( A1 => n769, A2 => n487, ZN => n455);
   U929 : OAI21_X1 port map( B1 => n721, B2 => n771, A => n616, ZN => n488);
   U930 : OAI21_X1 port map( B1 => n490, B2 => cu_i_n2, A => n488, ZN => n454);
   U931 : MUX2_X1 port map( A => n455, B => n454, S => cu_i_n151, Z => 
                           cu_i_N277);
   U932 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_31_port, B1 => 
                           datapath_i_new_pc_value_decode_31_port, B2 => n511, 
                           ZN => n456);
   U933 : OAI21_X1 port map( B1 => n729, B2 => n458, A => n456, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U934 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_30_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_30_port, ZN => 
                           n457);
   U935 : OAI21_X1 port map( B1 => n458, B2 => n714, A => n457, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   datapath_i_execute_stage_dp_n9 <= '0';
   U937 : NOR2_X1 port map( A1 => n715, A2 => n459, ZN => n460);
   U938 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => n468
                           , B1 => n460, B2 => n475, ZN => n466);
   U939 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => n726, 
                           ZN => n493);
   U940 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => 
                           curr_instruction_to_cu_i_3_port, A3 => n504, A4 => 
                           n728, ZN => n479);
   U941 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => n718, 
                           ZN => n470);
   U942 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_4_port, ZN => n492);
   U943 : NAND2_X1 port map( A1 => n502, A2 => n492, ZN => n467);
   U944 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => 
                           curr_instruction_to_cu_i_1_port, A3 => n504, A4 => 
                           n728, ZN => n461);
   U945 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => n461,
                           ZN => n486);
   U946 : INV_X1 port map( A => n479, ZN => n462);
   U947 : OAI211_X1 port map( C1 => n726, C2 => n467, A => n486, B => n462, ZN 
                           => n463);
   U948 : AOI22_X1 port map( A1 => n493, A2 => n479, B1 => n470, B2 => n463, ZN
                           => n465);
   U949 : NAND3_X1 port map( A1 => n466, A2 => n465, A3 => n464, ZN => 
                           cu_i_N264);
   U950 : NOR2_X1 port map( A1 => n467, A2 => curr_instruction_to_cu_i_5_port, 
                           ZN => n469);
   U951 : AOI21_X1 port map( B1 => n469, B2 => n470, A => n468, ZN => n483);
   U952 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n770, 
                           A3 => n486, ZN => n472);
   U953 : AND3_X1 port map( A1 => n726, A2 => n479, A3 => n470, ZN => n471);
   U954 : AOI211_X1 port map( C1 => n480, C2 => n473, A => n472, B => n471, ZN 
                           => n478);
   U955 : INV_X1 port map( A => n474, ZN => n481);
   U956 : NAND3_X1 port map( A1 => n481, A2 => n475, A3 => n715, ZN => n476);
   U957 : NAND4_X1 port map( A1 => n483, A2 => n478, A3 => n477, A4 => n476, ZN
                           => cu_i_N265);
   U958 : OAI221_X1 port map( B1 => n493, B2 => curr_instruction_to_cu_i_0_port
                           , C1 => n493, C2 => n726, A => n479, ZN => n484);
   U959 : OAI221_X1 port map( B1 => n481, B2 => 
                           curr_instruction_to_cu_i_27_port, C1 => n481, C2 => 
                           n706, A => n480, ZN => n482);
   U960 : OAI211_X1 port map( C1 => n718, C2 => n484, A => n483, B => n482, ZN 
                           => cu_i_N266);
   U961 : OAI221_X1 port map( B1 => n486, B2 => n770, C1 => n486, C2 => n718, A
                           => n485, ZN => cu_i_N267);
   U962 : NAND2_X1 port map( A1 => n669, A2 => n490, ZN => cu_i_N274);
   U963 : AOI221_X1 port map( B1 => cu_i_n152, B2 => cu_i_n4, C1 => n721, C2 =>
                           n771, A => n490, ZN => cu_i_N275);
   U964 : NOR2_X1 port map( A1 => cu_i_n152, A2 => n490, ZN => cu_i_N273);
   U965 : AOI22_X1 port map( A1 => cu_i_n2, A2 => n488, B1 => n487, B2 => n769,
                           ZN => cu_i_N276);
   U966 : INV_X1 port map( A => n489, ZN => n615);
   U967 : AOI211_X1 port map( C1 => n669, C2 => cu_i_n145, A => n615, B => n490
                           , ZN => cu_i_N279);
   U968 : NAND2_X1 port map( A1 => n491, A2 => n706, ZN => n496);
   U969 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_5_port, A2 => n493,
                           A3 => n492, A4 => n718, ZN => n494);
   U970 : OAI22_X1 port map( A1 => n497, A2 => n496, B1 => n495, B2 => n494, ZN
                           => cu_i_cmd_word_8_port);
   U971 : MUX2_X1 port map( A => cu_i_cw1_12_port, B => cu_i_cmd_word_8_port, S
                           => n669, Z => alu_cin_i);
   U972 : MUX2_X1 port map( A => cu_i_cw1_4_port, B => cu_i_cw2_4_port, S => 
                           n669, Z => cu_i_cw1_i_4_port);
   U973 : MUX2_X1 port map( A => cu_i_cw1_7_port, B => cu_i_cw2_7_port, S => 
                           n669, Z => cu_i_cw1_i_7_port);
   U974 : MUX2_X1 port map( A => cu_i_cw1_8_port, B => cu_i_cw2_8_port, S => 
                           n719, Z => cu_i_cw1_i_8_port);
   U975 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_12_port, A2 => 
                           curr_instruction_to_cu_i_11_port, A3 => 
                           curr_instruction_to_cu_i_15_port, A4 => 
                           curr_instruction_to_cu_i_14_port, ZN => n498);
   U976 : NAND2_X1 port map( A1 => n498, A2 => n760, ZN => n503);
   U977 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_17_port, A2 => 
                           curr_instruction_to_cu_i_16_port, A3 => 
                           curr_instruction_to_cu_i_20_port, A4 => 
                           curr_instruction_to_cu_i_19_port, ZN => n500);
   U978 : AOI21_X1 port map( B1 => n500, B2 => n720, A => n499, ZN => n501);
   U979 : AOI221_X1 port map( B1 => n505, B2 => n504, C1 => n503, C2 => n502, A
                           => n501, ZN => n508);
   U980 : NOR2_X1 port map( A1 => cu_i_cmd_word_4_port, A2 => cu_i_n135, ZN => 
                           n507);
   U981 : OAI211_X1 port map( C1 => n508, C2 => n609, A => n507, B => n506, ZN 
                           => cu_i_n209);
   U982 : AND2_X1 port map( A1 => cu_i_n3, A2 => cu_i_n153, ZN => cu_i_n210);
   U983 : MUX2_X1 port map( A => cu_i_cw1_6_port, B => cu_i_cw2_6_port, S => 
                           n719, Z => cu_i_n128);
   U984 : MUX2_X1 port map( A => cu_i_cw1_5_port, B => cu_i_cw2_5_port, S => 
                           n719, Z => cu_i_n127);
   U985 : MUX2_X1 port map( A => IRAM_DATA(31), B => 
                           curr_instruction_to_cu_i_31_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U986 : MUX2_X1 port map( A => IRAM_DATA(30), B => 
                           curr_instruction_to_cu_i_30_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U987 : MUX2_X1 port map( A => IRAM_DATA(29), B => 
                           curr_instruction_to_cu_i_29_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U988 : MUX2_X1 port map( A => IRAM_DATA(28), B => 
                           curr_instruction_to_cu_i_28_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U989 : MUX2_X1 port map( A => IRAM_DATA(27), B => 
                           curr_instruction_to_cu_i_27_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U990 : MUX2_X1 port map( A => IRAM_DATA(26), B => 
                           curr_instruction_to_cu_i_26_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U991 : MUX2_X1 port map( A => IRAM_DATA(25), B => datapath_i_n9, S => n719, 
                           Z => datapath_i_fetch_stage_dp_n63);
   U992 : MUX2_X1 port map( A => IRAM_DATA(24), B => datapath_i_n10, S => n719,
                           Z => datapath_i_fetch_stage_dp_n62);
   U993 : MUX2_X1 port map( A => IRAM_DATA(23), B => datapath_i_n11, S => n669,
                           Z => datapath_i_fetch_stage_dp_n61);
   U994 : MUX2_X1 port map( A => IRAM_DATA(22), B => datapath_i_n12, S => n669,
                           Z => datapath_i_fetch_stage_dp_n60);
   U995 : MUX2_X1 port map( A => IRAM_DATA(21), B => datapath_i_n13, S => n669,
                           Z => datapath_i_fetch_stage_dp_n59);
   U996 : MUX2_X1 port map( A => IRAM_DATA(20), B => 
                           curr_instruction_to_cu_i_20_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U997 : MUX2_X1 port map( A => IRAM_DATA(19), B => 
                           curr_instruction_to_cu_i_19_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U998 : MUX2_X1 port map( A => IRAM_DATA(18), B => 
                           curr_instruction_to_cu_i_18_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n56);
   U999 : MUX2_X1 port map( A => IRAM_DATA(17), B => 
                           curr_instruction_to_cu_i_17_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U1000 : MUX2_X1 port map( A => IRAM_DATA(16), B => 
                           curr_instruction_to_cu_i_16_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U1001 : MUX2_X1 port map( A => IRAM_DATA(15), B => 
                           curr_instruction_to_cu_i_15_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U1002 : MUX2_X1 port map( A => IRAM_DATA(14), B => 
                           curr_instruction_to_cu_i_14_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U1003 : MUX2_X1 port map( A => IRAM_DATA(13), B => 
                           curr_instruction_to_cu_i_13_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n51);
   U1004 : MUX2_X1 port map( A => IRAM_DATA(12), B => 
                           curr_instruction_to_cu_i_12_port, S => n669, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U1005 : MUX2_X1 port map( A => IRAM_DATA(11), B => 
                           curr_instruction_to_cu_i_11_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U1006 : MUX2_X1 port map( A => IRAM_DATA(10), B => datapath_i_n14, S => n719
                           , Z => datapath_i_fetch_stage_dp_n48);
   U1007 : MUX2_X1 port map( A => IRAM_DATA(9), B => datapath_i_n15, S => n719,
                           Z => datapath_i_fetch_stage_dp_n47);
   U1008 : MUX2_X1 port map( A => IRAM_DATA(8), B => datapath_i_n16, S => n719,
                           Z => datapath_i_fetch_stage_dp_n46);
   U1009 : MUX2_X1 port map( A => IRAM_DATA(7), B => datapath_i_n17, S => n719,
                           Z => datapath_i_fetch_stage_dp_n45);
   U1010 : MUX2_X1 port map( A => IRAM_DATA(6), B => datapath_i_n18, S => n719,
                           Z => datapath_i_fetch_stage_dp_n44);
   U1011 : MUX2_X1 port map( A => IRAM_DATA(5), B => 
                           curr_instruction_to_cu_i_5_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U1012 : MUX2_X1 port map( A => IRAM_DATA(4), B => 
                           curr_instruction_to_cu_i_4_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U1013 : MUX2_X1 port map( A => IRAM_DATA(3), B => 
                           curr_instruction_to_cu_i_3_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U1014 : MUX2_X1 port map( A => IRAM_DATA(2), B => 
                           curr_instruction_to_cu_i_2_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U1015 : MUX2_X1 port map( A => IRAM_DATA(1), B => 
                           curr_instruction_to_cu_i_1_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U1016 : MUX2_X1 port map( A => IRAM_DATA(0), B => 
                           curr_instruction_to_cu_i_0_port, S => n719, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U1017 : AOI22_X1 port map( A1 => n509, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_0_port, ZN => n510
                           );
   U1018 : OAI21_X1 port map( B1 => n513, B2 => n751, A => n510, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U1019 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N5, B => 
                           datapath_i_fetch_stage_dp_N39_port, S => n607, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U1020 : AOI22_X1 port map( A1 => n717, A2 => 
                           datapath_i_alu_output_val_i_1_port, B1 => n511, B2 
                           => datapath_i_new_pc_value_decode_1_port, ZN => n512
                           );
   U1021 : OAI21_X1 port map( B1 => n513, B2 => n752, A => n512, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U1022 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N6, B => 
                           datapath_i_fetch_stage_dp_N40_port, S => n607, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U1023 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n514, ZN => n515);
   U1024 : AOI22_X1 port map( A1 => n607, A2 => n515, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n597, ZN => datapath_i_fetch_stage_dp_n35);
   U1025 : OAI21_X1 port map( B1 => n516, B2 => IRAM_ADDRESS_3_port, A => n607,
                           ZN => n518);
   U1026 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_3_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, ZN
                           => n520);
   U1027 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_3_port,
                           B2 => datapath_i_new_pc_value_mem_stage_i_2_port, A 
                           => n597, ZN => n517);
   U1028 : OAI22_X1 port map( A1 => n522, A2 => n518, B1 => n520, B2 => n517, 
                           ZN => datapath_i_fetch_stage_dp_n34);
   U1029 : OAI211_X1 port map( C1 => n520, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n597, B => n519, ZN => n524);
   U1030 : OAI211_X1 port map( C1 => n522, C2 => IRAM_ADDRESS_4_port, A => n607
                           , B => n521, ZN => n523);
   U1031 : NAND2_X1 port map( A1 => n524, A2 => n523, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U1032 : OAI211_X1 port map( C1 => n526, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n597, B => n525, ZN => n530);
   U1033 : OAI211_X1 port map( C1 => n528, C2 => IRAM_ADDRESS_6_port, A => n599
                           , B => n527, ZN => n529);
   U1034 : NAND2_X1 port map( A1 => n530, A2 => n529, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U1035 : OAI211_X1 port map( C1 => n532, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n597, B => n531, ZN => n536);
   U1036 : OAI211_X1 port map( C1 => n534, C2 => IRAM_ADDRESS_8_port, A => n599
                           , B => n533, ZN => n535);
   U1037 : NAND2_X1 port map( A1 => n536, A2 => n535, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U1038 : OAI211_X1 port map( C1 => n538, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n597, B => n537, ZN => n542);
   U1039 : OAI211_X1 port map( C1 => n540, C2 => IRAM_ADDRESS_10_port, A => 
                           n599, B => n539, ZN => n541);
   U1040 : NAND2_X1 port map( A1 => n542, A2 => n541, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U1041 : OAI211_X1 port map( C1 => n544, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n597, B => n543, ZN => n548);
   U1042 : OAI211_X1 port map( C1 => n546, C2 => IRAM_ADDRESS_12_port, A => 
                           n599, B => n545, ZN => n547);
   U1043 : NAND2_X1 port map( A1 => n548, A2 => n547, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U1044 : OAI211_X1 port map( C1 => n550, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n597, B => n549, ZN => n554);
   U1045 : OAI211_X1 port map( C1 => n552, C2 => IRAM_ADDRESS_14_port, A => 
                           n599, B => n551, ZN => n553);
   U1046 : NAND2_X1 port map( A1 => n554, A2 => n553, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U1047 : OAI211_X1 port map( C1 => n556, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n597, B => n555, ZN => n560);
   U1048 : OAI211_X1 port map( C1 => n558, C2 => IRAM_ADDRESS_16_port, A => 
                           n599, B => n557, ZN => n559);
   U1049 : NAND2_X1 port map( A1 => n560, A2 => n559, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U1050 : OAI211_X1 port map( C1 => n562, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n597, B => n561, ZN => n566);
   U1051 : OAI211_X1 port map( C1 => n564, C2 => IRAM_ADDRESS_18_port, A => 
                           n599, B => n563, ZN => n565);
   U1052 : NAND2_X1 port map( A1 => n566, A2 => n565, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U1053 : OAI211_X1 port map( C1 => n568, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n597, B => n567, ZN => n572);
   U1054 : OAI211_X1 port map( C1 => n570, C2 => IRAM_ADDRESS_20_port, A => 
                           n599, B => n569, ZN => n571);
   U1055 : NAND2_X1 port map( A1 => n572, A2 => n571, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U1056 : OAI211_X1 port map( C1 => n574, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n597, B => n573, ZN => n578);
   U1057 : OAI211_X1 port map( C1 => n576, C2 => IRAM_ADDRESS_22_port, A => 
                           n607, B => n575, ZN => n577);
   U1058 : NAND2_X1 port map( A1 => n578, A2 => n577, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U1059 : OAI211_X1 port map( C1 => n580, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n597, B => n579, ZN => n584);
   U1060 : OAI211_X1 port map( C1 => n582, C2 => IRAM_ADDRESS_24_port, A => 
                           n599, B => n581, ZN => n583);
   U1061 : NAND2_X1 port map( A1 => n584, A2 => n583, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U1062 : OAI211_X1 port map( C1 => n586, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n597, B => n585, ZN => n590);
   U1063 : OAI211_X1 port map( C1 => n588, C2 => IRAM_ADDRESS_26_port, A => 
                           n599, B => n587, ZN => n589);
   U1064 : NAND2_X1 port map( A1 => n590, A2 => n589, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U1065 : OAI211_X1 port map( C1 => n592, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n597, B => n591, ZN => n596);
   U1066 : OAI211_X1 port map( C1 => n594, C2 => IRAM_ADDRESS_28_port, A => 
                           n607, B => n593, ZN => n595);
   U1067 : NAND2_X1 port map( A1 => n596, A2 => n595, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U1068 : NAND2_X1 port map( A1 => n598, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n604);
   U1069 : OAI211_X1 port map( C1 => n598, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n597, B => n604, ZN => n602);
   U1070 : NAND2_X1 port map( A1 => n600, A2 => n778, ZN => n603);
   U1071 : OAI211_X1 port map( C1 => n600, C2 => IRAM_ADDRESS_30_port, A => 
                           n599, B => n603, ZN => n601);
   U1072 : NAND2_X1 port map( A1 => n602, A2 => n601, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U1073 : XOR2_X1 port map( A => n328, B => n603, Z => n606);
   U1074 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n604, Z => n605);
   U1075 : AOI22_X1 port map( A1 => n607, A2 => n606, B1 => n605, B2 => n597, 
                           ZN => datapath_i_fetch_stage_dp_n2);
   U1076 : AND2_X1 port map( A1 => n772, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U1077 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => 
                           curr_instruction_to_cu_i_26_port, A3 => 
                           curr_instruction_to_cu_i_29_port, A4 => n608, ZN => 
                           n610);
   U1078 : OAI21_X1 port map( B1 => n610, B2 => n609, A => n612, ZN => 
                           read_rf_p2_i);
   U1079 : OAI221_X1 port map( B1 => n613, B2 => n720, C1 => n612, C2 => n760, 
                           A => n611, ZN => datapath_i_decode_stage_dp_n79);
   U1080 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ZN => n614);
   U1081 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n614, ZN => n618);
   U1082 : INV_X2 port map( A => n618, ZN => n654);
   U1083 : AND2_X2 port map( A1 => n654, A2 => n617, ZN => n644);
   U1084 : NOR2_X1 port map( A1 => n618, A2 => n617, ZN => n637);
   U1085 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_0_port, ZN => n619);
   U1086 : OAI21_X1 port map( B1 => n751, B2 => n654, A => n619, ZN => 
                           datapath_i_decode_stage_dp_n44);
   U1087 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_1_port, ZN => n620);
   U1088 : OAI21_X1 port map( B1 => n752, B2 => n654, A => n620, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U1089 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_2_port, ZN => n621);
   U1090 : OAI21_X1 port map( B1 => n746, B2 => n654, A => n621, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U1091 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_3_port, ZN => n622);
   U1092 : OAI21_X1 port map( B1 => n747, B2 => n654, A => n622, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U1093 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_4_port, ZN => n623);
   U1094 : OAI21_X1 port map( B1 => n748, B2 => n654, A => n623, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U1095 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n637, B2
                           => datapath_i_data_from_alu_i_5_port, ZN => n624);
   U1096 : OAI21_X1 port map( B1 => n749, B2 => n654, A => n624, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U1097 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n637, B2
                           => datapath_i_data_from_alu_i_6_port, ZN => n625);
   U1098 : OAI21_X1 port map( B1 => n750, B2 => n654, A => n625, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U1099 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_7_port, ZN => n626);
   U1100 : OAI21_X1 port map( B1 => n730, B2 => n654, A => n626, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U1101 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n652, B2
                           => datapath_i_data_from_alu_i_8_port, ZN => n627);
   U1102 : OAI21_X1 port map( B1 => n731, B2 => n654, A => n627, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U1103 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n637, B2
                           => datapath_i_data_from_alu_i_9_port, ZN => n628);
   U1104 : OAI21_X1 port map( B1 => n732, B2 => n654, A => n628, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U1105 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => n629
                           );
   U1106 : OAI21_X1 port map( B1 => n733, B2 => n654, A => n629, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U1107 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => n630
                           );
   U1108 : OAI21_X1 port map( B1 => n734, B2 => n654, A => n630, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U1109 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => n631
                           );
   U1110 : OAI21_X1 port map( B1 => n735, B2 => n654, A => n631, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U1111 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => n632
                           );
   U1112 : OAI21_X1 port map( B1 => n736, B2 => n654, A => n632, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U1113 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => n633
                           );
   U1114 : OAI21_X1 port map( B1 => n737, B2 => n654, A => n633, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U1115 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => n634
                           );
   U1116 : OAI21_X1 port map( B1 => n738, B2 => n654, A => n634, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U1117 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => n635
                           );
   U1118 : OAI21_X1 port map( B1 => n739, B2 => n654, A => n635, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U1119 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => n636
                           );
   U1120 : OAI21_X1 port map( B1 => n740, B2 => n654, A => n636, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U1121 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n637, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => n638
                           );
   U1122 : OAI21_X1 port map( B1 => n741, B2 => n654, A => n638, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U1123 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => n639
                           );
   U1124 : OAI21_X1 port map( B1 => n742, B2 => n654, A => n639, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U1125 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => n640
                           );
   U1126 : OAI21_X1 port map( B1 => n743, B2 => n654, A => n640, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U1127 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => n641
                           );
   U1128 : OAI21_X1 port map( B1 => n744, B2 => n654, A => n641, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U1129 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => n642
                           );
   U1130 : OAI21_X1 port map( B1 => n745, B2 => n654, A => n642, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U1131 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => n643
                           );
   U1132 : OAI21_X1 port map( B1 => n707, B2 => n654, A => n643, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U1133 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => n645
                           );
   U1134 : OAI21_X1 port map( B1 => n708, B2 => n654, A => n645, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U1135 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => n646
                           );
   U1136 : OAI21_X1 port map( B1 => n709, B2 => n654, A => n646, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U1137 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => n647
                           );
   U1138 : OAI21_X1 port map( B1 => n710, B2 => n654, A => n647, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U1139 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => n648
                           );
   U1140 : OAI21_X1 port map( B1 => n711, B2 => n654, A => n648, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U1141 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => n649
                           );
   U1142 : OAI21_X1 port map( B1 => n712, B2 => n654, A => n649, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U1143 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => n650
                           );
   U1144 : OAI21_X1 port map( B1 => n713, B2 => n654, A => n650, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U1145 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => n651
                           );
   U1146 : OAI21_X1 port map( B1 => n714, B2 => n654, A => n651, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U1147 : AOI22_X1 port map( A1 => n644, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n652, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => n653
                           );
   U1148 : OAI21_X1 port map( B1 => n729, B2 => n654, A => n653, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U1149 : AOI21_X1 port map( B1 => n675, B2 => n656, A => n655, ZN => n657);
   U1150 : NOR2_X1 port map( A1 => n658, A2 => n657, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U1151 : AOI22_X1 port map( A1 => n669, A2 => cu_i_cmd_word_6_port, B1 => 
                           cu_i_cw1_10_port, B2 => n759, ZN => n673);
   U1152 : NOR4_X1 port map( A1 => datapath_i_val_a_i_15_port, A2 => 
                           datapath_i_val_a_i_16_port, A3 => 
                           datapath_i_val_a_i_17_port, A4 => 
                           datapath_i_val_a_i_18_port, ZN => n662);
   U1153 : NOR4_X1 port map( A1 => datapath_i_val_a_i_19_port, A2 => 
                           datapath_i_val_a_i_20_port, A3 => 
                           datapath_i_val_a_i_21_port, A4 => 
                           datapath_i_val_a_i_22_port, ZN => n661);
   U1154 : NOR4_X1 port map( A1 => datapath_i_val_a_i_7_port, A2 => 
                           datapath_i_val_a_i_8_port, A3 => 
                           datapath_i_val_a_i_9_port, A4 => 
                           datapath_i_val_a_i_10_port, ZN => n660);
   U1155 : NOR4_X1 port map( A1 => datapath_i_val_a_i_11_port, A2 => 
                           datapath_i_val_a_i_12_port, A3 => 
                           datapath_i_val_a_i_13_port, A4 => 
                           datapath_i_val_a_i_14_port, ZN => n659);
   U1156 : NAND4_X1 port map( A1 => n662, A2 => n661, A3 => n660, A4 => n659, 
                           ZN => n668);
   U1157 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n666);
   U1158 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n665);
   U1159 : NOR4_X1 port map( A1 => datapath_i_val_a_i_23_port, A2 => 
                           datapath_i_val_a_i_24_port, A3 => 
                           datapath_i_val_a_i_25_port, A4 => 
                           datapath_i_val_a_i_26_port, ZN => n664);
   U1160 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n663);
   U1161 : NAND4_X1 port map( A1 => n666, A2 => n665, A3 => n664, A4 => n663, 
                           ZN => n667);
   U1162 : NOR2_X1 port map( A1 => n668, A2 => n667, ZN => n671);
   U1163 : AOI22_X1 port map( A1 => n669, A2 => cu_i_cmd_word_7_port, B1 => 
                           cu_i_cw1_11_port, B2 => n759, ZN => n670);
   U1164 : NAND2_X1 port map( A1 => n671, A2 => n670, ZN => n672);
   U1165 : OAI22_X1 port map( A1 => n673, A2 => n672, B1 => n671, B2 => n670, 
                           ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U1166 : NOR2_X1 port map( A1 => n675, A2 => n674, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U1167 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U1168 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U1169 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U1170 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U1171 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U1172 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U1173 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U1174 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n776, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U1175 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U1176 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U1177 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U1178 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U1179 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U1180 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U1181 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U1182 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U1183 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U1184 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U1185 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_25_port
                           );
   U1186 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, S 
                           => n775, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_26_port
                           );
   U1187 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U1188 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_27_port
                           );
   U1189 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_28_port
                           );
   U1190 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_29_port
                           );
   U1191 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_30_port
                           );
   U1192 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U1193 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U1194 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U1195 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U1196 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U1197 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U1198 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n774, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U1199 : MUX2_X1 port map( A => datapath_i_val_immediate_i_7_port, B => 
                           datapath_i_val_b_i_7_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U1200 : MUX2_X1 port map( A => datapath_i_val_immediate_i_8_port, B => 
                           datapath_i_val_b_i_8_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U1201 : MUX2_X1 port map( A => datapath_i_val_immediate_i_9_port, B => 
                           datapath_i_val_b_i_9_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U1202 : MUX2_X1 port map( A => datapath_i_val_immediate_i_10_port, B => 
                           datapath_i_val_b_i_10_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U1203 : MUX2_X1 port map( A => datapath_i_val_immediate_i_11_port, B => 
                           datapath_i_val_b_i_11_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U1204 : MUX2_X1 port map( A => datapath_i_val_immediate_i_12_port, B => 
                           datapath_i_val_b_i_12_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U1205 : MUX2_X1 port map( A => datapath_i_val_immediate_i_13_port, B => 
                           datapath_i_val_b_i_13_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U1206 : MUX2_X1 port map( A => datapath_i_val_immediate_i_14_port, B => 
                           datapath_i_val_b_i_14_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U1207 : MUX2_X1 port map( A => datapath_i_val_immediate_i_15_port, B => 
                           datapath_i_val_b_i_15_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U1208 : MUX2_X1 port map( A => datapath_i_val_immediate_i_16_port, B => 
                           datapath_i_val_b_i_16_port, S => n676, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U1209 : MUX2_X1 port map( A => datapath_i_val_immediate_i_17_port, B => 
                           datapath_i_val_b_i_17_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U1210 : MUX2_X1 port map( A => datapath_i_val_immediate_i_18_port, B => 
                           datapath_i_val_b_i_18_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U1211 : MUX2_X1 port map( A => datapath_i_val_immediate_i_19_port, B => 
                           datapath_i_val_b_i_19_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U1212 : MUX2_X1 port map( A => datapath_i_val_immediate_i_20_port, B => 
                           datapath_i_val_b_i_20_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U1213 : MUX2_X1 port map( A => datapath_i_val_immediate_i_21_port, B => 
                           datapath_i_val_b_i_21_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U1214 : MUX2_X1 port map( A => datapath_i_val_immediate_i_22_port, B => 
                           datapath_i_val_b_i_22_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U1215 : MUX2_X1 port map( A => datapath_i_val_immediate_i_23_port, B => 
                           datapath_i_val_b_i_23_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U1216 : MUX2_X1 port map( A => datapath_i_val_immediate_i_24_port, B => 
                           datapath_i_val_b_i_24_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U1217 : MUX2_X1 port map( A => datapath_i_val_immediate_i_25_port, B => 
                           datapath_i_val_b_i_25_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U1218 : MUX2_X1 port map( A => datapath_i_val_immediate_i_26_port, B => 
                           datapath_i_val_b_i_26_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U1219 : MUX2_X1 port map( A => datapath_i_val_immediate_i_27_port, B => 
                           datapath_i_val_b_i_27_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U1220 : MUX2_X1 port map( A => datapath_i_val_immediate_i_28_port, B => 
                           datapath_i_val_b_i_28_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U1221 : MUX2_X1 port map( A => datapath_i_val_immediate_i_29_port, B => 
                           datapath_i_val_b_i_29_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U1222 : MUX2_X1 port map( A => datapath_i_val_immediate_i_30_port, B => 
                           datapath_i_val_b_i_30_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U1223 : MUX2_X1 port map( A => datapath_i_val_immediate_i_31_port, B => 
                           datapath_i_val_b_i_31_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U1224 : MUX2_X1 port map( A => datapath_i_val_immediate_i_3_port, B => 
                           datapath_i_val_b_i_3_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U1225 : MUX2_X1 port map( A => datapath_i_val_immediate_i_4_port, B => 
                           datapath_i_val_b_i_4_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U1226 : MUX2_X1 port map( A => datapath_i_val_immediate_i_5_port, B => 
                           datapath_i_val_b_i_5_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U1227 : MUX2_X1 port map( A => datapath_i_val_immediate_i_6_port, B => 
                           datapath_i_val_b_i_6_port, S => n677, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U1228 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n698, B1 => datapath_i_val_a_i_7_port, B2 => n702
                           , ZN => n678);
   U1229 : OAI21_X1 port map( B1 => n730, B2 => n705, A => n678, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U1230 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n698, B1 => datapath_i_val_a_i_9_port, B2 => n702
                           , ZN => n679);
   U1231 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n698, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n702, ZN => n680);
   U1232 : OAI21_X1 port map( B1 => n736, B2 => n705, A => n680, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U1233 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n698, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n702, ZN => n681);
   U1234 : OAI21_X1 port map( B1 => n737, B2 => n705, A => n681, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U1235 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n698, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n702, ZN => n682);
   U1236 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n698, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n702, ZN => n683);
   U1237 : OAI21_X1 port map( B1 => n740, B2 => n705, A => n683, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U1238 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n703, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n702, ZN => n684);
   U1239 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n703, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n702, ZN => n685);
   U1240 : OAI21_X1 port map( B1 => n743, B2 => n705, A => n685, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U1241 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n703, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n702, ZN => n686);
   U1242 : OAI21_X1 port map( B1 => n744, B2 => n705, A => n686, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U1243 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n703, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n702, ZN => n687);
   U1244 : OAI21_X1 port map( B1 => n745, B2 => n705, A => n687, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U1245 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n703, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n702, ZN => n688);
   U1246 : OAI21_X1 port map( B1 => n707, B2 => n705, A => n688, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U1247 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n703, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n702, ZN => n689);
   U1248 : OAI21_X1 port map( B1 => n708, B2 => n705, A => n689, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U1249 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n698, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n702, ZN => n690);
   U1250 : OAI21_X1 port map( B1 => n709, B2 => n705, A => n690, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U1251 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n698, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n702, ZN => n691);
   U1252 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n698, B1 => datapath_i_val_a_i_0_port, B2 => n702
                           , ZN => n692);
   U1253 : OAI21_X1 port map( B1 => n705, B2 => n751, A => n692, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U1254 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n698, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n702, ZN => n693);
   U1255 : OAI21_X1 port map( B1 => n711, B2 => n705, A => n693, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U1256 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n698, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n702, ZN => n694);
   U1257 : OAI21_X1 port map( B1 => n712, B2 => n705, A => n694, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U1258 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n703, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n702, ZN => n695);
   U1259 : OAI21_X1 port map( B1 => n713, B2 => n705, A => n695, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U1260 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n698, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n702, ZN => n696);
   U1261 : OAI21_X1 port map( B1 => n714, B2 => n705, A => n696, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U1262 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n698, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n702, ZN => n697);
   U1263 : OAI21_X1 port map( B1 => n729, B2 => n705, A => n697, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U1264 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n698, B1 => datapath_i_val_a_i_1_port, B2 => n702
                           , ZN => n699);
   U1265 : OAI21_X1 port map( B1 => n705, B2 => n752, A => n699, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U1266 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n703, B1 => datapath_i_val_a_i_2_port, B2 => n702
                           , ZN => n700);
   U1267 : OAI21_X1 port map( B1 => n746, B2 => n705, A => n700, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U1268 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n703, B1 => datapath_i_val_a_i_3_port, B2 => n702
                           , ZN => n701);
   U1269 : OAI21_X1 port map( B1 => n747, B2 => n705, A => n701, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U1270 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n703, B1 => datapath_i_val_a_i_5_port, B2 => n702
                           , ZN => n704);
   U1271 : OAI21_X1 port map( B1 => n749, B2 => n705, A => n704, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);

end SYN_dlx_rtl;
