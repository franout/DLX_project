
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal DATA2_I_30_port, DATA2_I_28_port, DATA2_I_27_port, DATA2_I_26_port, 
      DATA2_I_25_port, DATA2_I_24_port, DATA2_I_23_port, DATA2_I_22_port, 
      DATA2_I_21_port, DATA2_I_20_port, DATA2_I_19_port, DATA2_I_18_port, 
      DATA2_I_17_port, DATA2_I_16_port, DATA2_I_15_port, DATA2_I_14_port, 
      DATA2_I_13_port, DATA2_I_12_port, DATA2_I_11_port, DATA2_I_10_port, 
      DATA2_I_9_port, DATA2_I_8_port, DATA2_I_7_port, DATA2_I_6_port, 
      DATA2_I_5_port, DATA2_I_4_port, DATA2_I_3_port, DATA2_I_2_port, 
      DATA2_I_1_port, DATA2_I_0_port, data1_mul_15_port, data1_mul_0_port, 
      data2_mul_2_port, data2_mul_1_port, N2517, N2518, N2519, N2520, N2521, 
      N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n554, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1429, 
      n2808, n3020, n3026, n3027, n3028, n3029, n3030, n3036, n3940, n3957, 
      n3958, n3973, n3974, n3990, n3991, n3992, n3993, n3994, n3995, n4007, 
      n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4293, n4295, n4302, 
      n4395, n7769, n7822, n8626, n8732, n8733, n8734, n8735, n8736, n8737, 
      n8738, n8739, n8740, n8748, n8749, n8751, n8752, n8753, n8754, n8755, 
      n8764, n8928, n8978, n9045, n9048, n9051, n9054, n9057, n9060, n9063, 
      n9066, n9069, n9072, n9075, n9078, n9081, n9084, n11966, n12313, n12526, 
      n13963, n14004, n14058, n14059, n14060, n14061, n14062, n14063, n14064, 
      n14065, n14066, n14067, n14068, n14074, n14075, n14094, n14102, n14145, 
      n14286, n14287, n1809, n1894, n1896, n17503, n17932, n18839, n18845, 
      n18846, n18847, n18848, n18850, n18851, n18852, n18853, n18854, n18855, 
      n18856, n18860, n18861, n18867, n18872, n18877, n18878, n18882, n18892, 
      n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18902, n18903, 
      n18904, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, 
      n18917, n18918, n18920, n18921, n18922, n18923, n18925, n18926, n18927, 
      n18929, n18930, n18933, n18934, n18935, n18945, n18946, n18948, n18949, 
      n18950, n18952, n18954, n18964, n18965, n18967, n18968, n18969, n18972, 
      n18973, n18974, n18976, n18977, n18980, n18981, n18982, n18988, n18989, 
      n18992, n18993, n18999, n19000, n19001, n19003, n19004, n19005, n19010, 
      n19018, n19021, n19024, n19027, n19030, n19033, n19037, n19038, n19042, 
      n19047, n19051, n19055, n19059, n19063, n19067, n19071, n19075, n19079, 
      n19083, n19084, n19085, n19089, n19090, n19091, n19092, n19097, n19098, 
      n19099, n19100, n19105, n19106, n19107, n19108, n19113, n19114, n19115, 
      n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, 
      n19130, n19131, n19132, n19133, n19134, n19135, n19147, n19148, n19149, 
      n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, 
      n19160, n19161, n19162, n19163, n19164, n19165, n19168, n19169, n19170, 
      n19171, n19172, n19174, n19175, n19176, n19178, n19179, n19180, n19181, 
      n19182, n19183, n19184, n19185, n19186, n19187, n19194, n19200, n19202, 
      n19213, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, 
      n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, 
      n19248, n19250, n19251, n19252, n19253, n19259, n19261, n19262, n19264, 
      n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19277, 
      n19278, n19280, n19283, n19291, n19292, n19293, n19294, n19399, n19419, 
      n19433, n1806, n1816, n1826, n1836, n1841, n1843, n21296, n21378, n21379,
      n21484, n21485, n21490, n21491, n21556, n21603, n21604, n21607, n21633, 
      n21634, n21635, n21745, n21746, n21841, n21842, n21843, n21845, n22091, 
      n22276, n22281, n22313, n22526, n22532, n22765, n22797, n22800, n22802, 
      n22975, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, 
      n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, 
      n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, 
      n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, 
      n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, 
      n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, 
      n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, 
      n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, 
      n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, 
      n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, 
      n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23689, 
      n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, 
      n23699, n23700, n23701, n23702, n23703, n23705, n23706, n23707, n23708, 
      n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, 
      n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, 
      n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, 
      n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, 
      n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, 
      n23755, n23756, n23757, n23759, n23760, n23762, n23763, n23764, n23765, 
      n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, 
      n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, 
      n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, 
      n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, 
      n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, 
      n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, 
      n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, 
      n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, 
      n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, 
      n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, 
      n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, 
      n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, 
      n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, 
      n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, 
      n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, 
      n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, 
      n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, 
      n23919, n23920, n23922, n23923, n23924, n23925, n23926, n23927, n23928, 
      n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, 
      n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, 
      n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, 
      n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, 
      n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, 
      n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, 
      n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, 
      n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, 
      n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, 
      n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, 
      n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, 
      n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, 
      n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24046, 
      n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, 
      n24056, n24057, n24058, n24060, n24061, n24062, n24063, n24064, n24065, 
      n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, 
      n24075, n24076, n24077, n24079, n24080, n24081, n24082, n24083, n24084, 
      n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, 
      n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, 
      n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, 
      n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, 
      n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, 
      n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, 
      n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, 
      n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, 
      n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, 
      n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, 
      n24175, n24176, n24177, n24178, n24179, n24181, n25858, n25859, n25861, 
      n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, 
      n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, 
      n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1807, 
      n1808, n1810, n1811, n1812, n1813, n1814, n1815, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1827, n1828, n1829, n1830, 
      n1831, n1832, n1833, n1834, n1835, n1837, n1838, n1839, n1840, n1842, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
      n1864, n1865, n1866, n1868, n1869, n1870, n1871, n25889, n25890, n25891, 
      n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, 
      n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, 
      n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, 
      n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, 
      n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, 
      n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, 
      n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, 
      n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, 
      n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, 
      n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, 
      n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, 
      n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, 
      n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, 
      n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, 
      n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, 
      n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, 
      n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, 
      n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, 
      n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, 
      n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, 
      n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, 
      n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, 
      n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, 
      n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, 
      n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, 
      n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, 
      n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, 
      n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, 
      n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, 
      n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, 
      n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, 
      n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, 
      n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, 
      n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, 
      n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, 
      n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, 
      n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, 
      n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, 
      n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, 
      n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, 
      n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, 
      n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, 
      n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, 
      n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, 
      n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, 
      n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, 
      n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, 
      n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, 
      n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, 
      n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, 
      n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, 
      n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, 
      n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, 
      n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, 
      n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, 
      n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, 
      n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, 
      n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, 
      n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, 
      n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, 
      n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, 
      n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, 
      n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, 
      n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, 
      n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, 
      n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, 
      n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, 
      n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, 
      n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, 
      n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, 
      n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, 
      n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, 
      n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, 
      n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, 
      n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, 
      n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, 
      n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, 
      n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, 
      n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, 
      n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, 
      n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, 
      n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, 
      n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, 
      n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, 
      n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, 
      n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, 
      n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, 
      n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, 
      n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, 
      n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, 
      n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, 
      n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, 
      n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, 
      n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, 
      n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, 
      n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, 
      n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, 
      n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, 
      n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, 
      n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, 
      n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, 
      n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, 
      n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, 
      n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, 
      n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, 
      n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, 
      n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, 
      n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, 
      n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, 
      n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, 
      n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, 
      n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, 
      n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, 
      n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, 
      n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, 
      n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, 
      n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, 
      n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, 
      n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, 
      n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, 
      n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, 
      n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, 
      n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, 
      n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, 
      n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, 
      n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, 
      n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, 
      n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, 
      n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, 
      n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, 
      n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, 
      n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, 
      n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, 
      n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, 
      n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, 
      n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, 
      n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, 
      n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, 
      n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, 
      n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, 
      n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, 
      n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, 
      n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, 
      n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, 
      n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, 
      n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, 
      n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, 
      n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, 
      n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, 
      n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, 
      n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, 
      n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, 
      n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, 
      n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, 
      n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, 
      n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, 
      n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, 
      n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, 
      n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, 
      n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, 
      n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, 
      n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, 
      n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, 
      n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, 
      n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, 
      n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, 
      n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, 
      n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, 
      n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, 
      n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, 
      n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, 
      n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, 
      n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, 
      n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, 
      n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, 
      n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, 
      n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, 
      n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, 
      n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, 
      n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, 
      n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, 
      n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, 
      n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, 
      n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, 
      n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, 
      n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, 
      n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, 
      n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, 
      n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, 
      n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, 
      n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, 
      n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, 
      n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, 
      n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, 
      n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, 
      n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, 
      n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, 
      n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, 
      n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, 
      n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, 
      n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, 
      n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, 
      n27710, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, 
      n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, 
      n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, 
      n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, 
      n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, 
      n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, 
      n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, 
      n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, 
      n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, 
      n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, 
      n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, 
      n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, 
      n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, 
      n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, 
      n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, 
      n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, 
      n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, 
      n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, 
      n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, 
      n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, 
      n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, 
      n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, 
      n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, 
      n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, 
      n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, 
      n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, 
      n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, 
      n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, 
      n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, 
      n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, 
      n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, 
      n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, 
      n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, 
      n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, 
      n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, 
      n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, 
      n_1552, n_1553 : std_logic;

begin
   
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n554, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n554, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n554, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n27710, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n554, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n554, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n27710, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n554, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n554, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n27710, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n27710, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n554, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n554, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n554, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n554, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n554, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n554, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n554, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n554, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n554, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n554, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n554, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n554, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n554, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n554, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n27710, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n7822, Q => 
                           n9045);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n7822, Q => 
                           n9048);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n7822, Q => 
                           n9051);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n7822, Q => 
                           n9054);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n7822, Q => 
                           n9057);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n7822, Q => 
                           n9060);
   data1_mul_reg_8_inst : DLL_X1 port map( D => n24181, GN => n7822, Q => n9063
                           );
   data1_mul_reg_7_inst : DLL_X1 port map( D => n24179, GN => n7822, Q => n9066
                           );
   data1_mul_reg_6_inst : DLL_X1 port map( D => n24178, GN => n7822, Q => n9069
                           );
   data1_mul_reg_5_inst : DLL_X1 port map( D => n24177, GN => n7822, Q => n9072
                           );
   data1_mul_reg_4_inst : DLL_X1 port map( D => n24176, GN => n7822, Q => n9075
                           );
   data1_mul_reg_3_inst : DLL_X1 port map( D => n24048, GN => n7822, Q => n9078
                           );
   data1_mul_reg_2_inst : DLL_X1 port map( D => n24049, GN => n7822, Q => n9081
                           );
   data1_mul_reg_1_inst : DLL_X1 port map( D => n24175, GN => n7822, Q => n9084
                           );
   data1_mul_reg_0_inst : DLL_X1 port map( D => n24173, GN => n7822, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n7822, Q => 
                           n22975);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n7822, Q => 
                           n19294);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n7822, Q => 
                           n19293);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n7822, Q => 
                           n19292);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n7822, Q => 
                           n14287);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n7822, Q => 
                           n14286);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n7822, Q => 
                           n4302);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n7822, Q => 
                           n8978);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n7822, Q => 
                           n7769);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n7822, Q => 
                           n4295);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n7822, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n7822, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n27710, Q => n4293)
                           ;
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1805, B => n1807, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1804, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1803, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1802, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1800, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1799, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1798, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1797, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1796, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1795, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1794, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1793, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1792, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1791, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1790, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3036,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => n19135);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => n19134);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => n19133);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => n19132);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => n19131);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => n19130);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => n19129);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => n19128);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => n19127);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => n19126);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => n19125);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => n19124);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => n19123);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => n19122);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1004, S => n19121);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => n23879, 
                           CI => n3026, CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => n19115);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => n23878, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => n23877, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => n23876, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => n23875, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => n23874,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => n23873,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => n23872,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => n23871,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => n23870,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => n23869,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => n23868,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => n23867,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => n23866,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => n14102);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => n23866,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => n19114, S => n19113);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n18847, B => n23866, CI => n19114, CO => n_1005, S 
                           => boothmul_pipelined_i_sum_B_in_3_22_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3030,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => n19108);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => n4018);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => n4017);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => n4016);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => n4015);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => n4014);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => n4013);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => n4012);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => n8764);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => n14094, S => n19107);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n14145, B => n14102, CI => n14094, CO => n19106, S 
                           => n19105);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n23911, B => n23860, CI => n23852, CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n23910, B => n23859, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n23909, B => n23859, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n23598, B => n23859, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1006, S => n4007);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => n4018, 
                           CI => n3029, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => n19100);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => n4017, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => n4016, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => n8755);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => n4015, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => n8754);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => n4014, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => n8753);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => n4013, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => n8752);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => n4012, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => n8751, S => n19099);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n8928, B => n8764, CI => n8751, CO => n19098, S => 
                           n19097);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n23659, B => n23853, CI => n23844, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => n3995);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n23658, B => n23851, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => n3994);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n23657, B => boothmul_pipelined_i_sum_B_in_4_19_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => n3993);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n23656, B => boothmul_pipelined_i_sum_B_in_4_20_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => n3992);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n23655, B => boothmul_pipelined_i_sum_B_in_4_21_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => n3991, S => n3990);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n23654, B => n4007, CI => n3991, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n23653, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => n8749);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n23604, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1007, S => n8748);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => n8755, 
                           CI => n3028, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => n19092);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => n8754, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => n8753, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => n19091);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => n8752, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => n19090, S => n19089);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           n23908, B => n23845, CI => n23837, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => n8740);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n23907, B => n23843, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => n8739);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n23906, B => n3995, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => n8738);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n23905, B => n3994, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => n8737);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n23904, B => n3993, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => n8736);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n23903, B => n3992, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => n8735);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n23902, B => n3990, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => n8734);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n23901, B => boothmul_pipelined_i_sum_B_in_5_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => n8733, S => n8732);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n23900, B => n8749, CI => n8733, CO => n3974, S => 
                           n3973);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n23899, B => n8748, CI => n3974, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n23898, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => n14075);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n23597, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1008, S => n14074);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           n18851, B => n19091, CI => n3027, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => n19085);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           n23652, B => n23836, CI => n23835, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           n23651, B => n8740, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => n14068);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n23650, B => n8739, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => n14067);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n23649, B => n8738, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => n14066);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n23648, B => n8737, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => n14065);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n23647, B => n8736, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => n14064);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n23646, B => n8735, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => n14063);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n23645, B => n8734, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => n14062);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n23644, B => n8732, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => n14061);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n23643, B => n3973, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => n14060);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n23642, B => boothmul_pipelined_i_sum_B_in_6_24_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => n14059, S => n14058);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n23641, B => n14075, CI => n14059, CO => n3958, S =>
                           n3957);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n23640, B => n14074, CI => n3958, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n23639, B => n14074, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => n19084);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n23603, B => n14074, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1009, S => n19083);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           n23602, B => n14068, CI => n3020, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => n19079);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n23997, B => n14067, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => n19075);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n23996, B => n14066, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => n19071);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n23995, B => n14065, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => n19067);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n23994, B => n14064, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => n19063);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n23993, B => n14063, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => n19059);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n23992, B => n14062, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => n19055);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n23991, B => n14061, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => n19051);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n23990, B => n14060, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => n19047);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n23989, B => n14058, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => n19042);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n23988, B => n3957, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => n19038);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n23987, B => boothmul_pipelined_i_sum_B_in_7_26_port
                           , CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => n19037, S => n19033);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n23986, B => n19084, CI => n19037, CO => n3940, S =>
                           n19030);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n23985, B => n19083, CI => n3940, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => n19027);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           n23983, B => n23829, CI => n23776, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => n19024);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           n23981, B => n23829, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => n19021);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           n23981, B => n23829, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1010, S => n19018);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n7822, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n554, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n554, Q => n4395);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n554, Q => 
                           DATA2_I_28_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n554, Q => 
                           DATA2_I_27_port);
   clk_r_REG14058_S3 : DFFS_X1 port map( D => n1849, CK => clk, SN => rst_BAR, 
                           Q => n_1011, QN => n24181);
   clk_r_REG14094_S3 : DFFS_X1 port map( D => n1850, CK => clk, SN => rst_BAR, 
                           Q => n_1012, QN => n24179);
   clk_r_REG14439_S6 : DFFS_X1 port map( D => n1851, CK => clk, SN => rst_BAR, 
                           Q => n_1013, QN => n24178);
   clk_r_REG13655_S6 : DFFS_X1 port map( D => n1852, CK => clk, SN => rst_BAR, 
                           Q => n_1014, QN => n24177);
   clk_r_REG14338_S3 : DFFS_X1 port map( D => n1853, CK => clk, SN => rst_BAR, 
                           Q => n_1015, QN => n24176);
   clk_r_REG14978_S3 : DFFS_X1 port map( D => n1854, CK => clk, SN => rst_BAR, 
                           Q => n_1016, QN => n24175);
   clk_r_REG14980_S4 : DFFS_X1 port map( D => n24175, CK => clk, SN => rst_BAR,
                           Q => n24174, QN => n_1017);
   clk_r_REG16594_S5 : DFFS_X1 port map( D => n1855, CK => clk, SN => rst_BAR, 
                           Q => n_1018, QN => n24173);
   clk_r_REG16737_S2 : DFFS_X1 port map( D => n1871, CK => clk, SN => rst_BAR, 
                           Q => n_1019, QN => n24172);
   clk_r_REG14303_S3 : DFFR_X1 port map( D => n25892, CK => clk, RN => rst_BAR,
                           Q => n24171, QN => n_1020);
   clk_r_REG14344_S5 : DFFS_X1 port map( D => n1801, CK => clk, SN => rst_BAR, 
                           Q => n24170, QN => n_1021);
   clk_r_REG14320_S3 : DFFR_X1 port map( D => n1841, CK => clk, RN => rst_BAR, 
                           Q => n27680, QN => n24168);
   clk_r_REG16961_S7 : DFFR_X1 port map( D => n1832, CK => clk, RN => rst_BAR, 
                           Q => n24167, QN => n_1022);
   clk_r_REG13830_S4 : DFFR_X1 port map( D => n1788, CK => clk, RN => rst_BAR, 
                           Q => n24166, QN => n_1023);
   clk_r_REG14837_S3 : DFFR_X1 port map( D => DATA1(2), CK => clk, RN => 
                           rst_BAR, Q => n_1024, QN => n24165);
   clk_r_REG14697_S3 : DFFR_X1 port map( D => DATA1(3), CK => clk, RN => 
                           rst_BAR, Q => n_1025, QN => n24164);
   clk_r_REG14556_S8 : DFFS_X1 port map( D => n1840, CK => clk, SN => rst_BAR, 
                           Q => n24163, QN => n_1026);
   clk_r_REG14505_S4 : DFFR_X1 port map( D => n1786, CK => clk, RN => rst_BAR, 
                           Q => n24162, QN => n_1027);
   clk_r_REG16597_S7 : DFFS_X1 port map( D => n1807, CK => clk, SN => rst_BAR, 
                           Q => n24161, QN => n_1028);
   clk_r_REG16584_S7 : DFFR_X1 port map( D => n22313, CK => clk, RN => rst_BAR,
                           Q => n24160, QN => n_1029);
   clk_r_REG14524_S5 : DFFR_X1 port map( D => n1814, CK => clk, RN => rst_BAR, 
                           Q => n24159, QN => n_1030);
   clk_r_REG14329_S3 : DFFS_X1 port map( D => n1843, CK => clk, SN => rst_BAR, 
                           Q => n_1031, QN => n24157);
   clk_r_REG14309_S3 : DFFS_X1 port map( D => n27709, CK => clk, SN => rst_BAR,
                           Q => n24155, QN => n_1032);
   clk_r_REG14326_S3 : DFFS_X1 port map( D => n1857, CK => clk, SN => rst_BAR, 
                           Q => n24154, QN => n_1033);
   clk_r_REG14243_S3 : DFFR_X1 port map( D => n1836, CK => clk, RN => rst_BAR, 
                           Q => n_1034, QN => n24153);
   clk_r_REG14242_S3 : DFFS_X1 port map( D => n1836, CK => clk, SN => n25890, Q
                           => n_1035, QN => n24152);
   clk_r_REG14249_S3 : DFFR_X1 port map( D => n1894, CK => clk, RN => rst_BAR, 
                           Q => n27668, QN => n24151);
   clk_r_REG14233_S3 : DFFS_X1 port map( D => n1896, CK => clk, SN => rst_BAR, 
                           Q => n27692, QN => n24150);
   clk_r_REG14332_S3 : DFFR_X1 port map( D => n1858, CK => clk, RN => rst_BAR, 
                           Q => n24149, QN => n_1036);
   clk_r_REG14287_S4 : DFFS_X1 port map( D => n1839, CK => clk, SN => rst_BAR, 
                           Q => n24148, QN => n_1037);
   clk_r_REG14618_S3 : DFFS_X1 port map( D => n1831, CK => clk, SN => rst_BAR, 
                           Q => n24147, QN => n_1038);
   clk_r_REG14270_S4 : DFFR_X1 port map( D => n1834, CK => clk, RN => rst_BAR, 
                           Q => n24146, QN => n_1039);
   clk_r_REG14269_S4 : DFFS_X1 port map( D => n1834, CK => clk, SN => n25890, Q
                           => n24145, QN => n_1040);
   clk_r_REG14262_S4 : DFFS_X1 port map( D => n1845, CK => clk, SN => rst_BAR, 
                           Q => n24144, QN => n_1041);
   clk_r_REG14266_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => n25890, Q
                           => n24143, QN => n_1042);
   clk_r_REG14296_S3 : DFFS_X1 port map( D => n1819, CK => clk, SN => rst_BAR, 
                           Q => n24142, QN => n_1043);
   clk_r_REG14293_S4 : DFFS_X1 port map( D => n1827, CK => clk, SN => n25890, Q
                           => n24141, QN => n_1044);
   clk_r_REG14116_S4 : DFFS_X1 port map( D => n1817, CK => clk, SN => rst_BAR, 
                           Q => n24140, QN => n_1045);
   clk_r_REG14272_S3 : DFFS_X1 port map( D => n1818, CK => clk, SN => rst_BAR, 
                           Q => n24139, QN => n_1046);
   clk_r_REG14291_S3 : DFFS_X1 port map( D => n1838, CK => clk, SN => n25890, Q
                           => n24138, QN => n_1047);
   clk_r_REG14264_S3 : DFFS_X1 port map( D => n1847, CK => clk, SN => n25890, Q
                           => n24137, QN => n_1048);
   clk_r_REG14263_S3 : DFFS_X1 port map( D => n1823, CK => clk, SN => rst_BAR, 
                           Q => n24136, QN => n_1049);
   clk_r_REG14103_S4 : DFFR_X1 port map( D => n1820, CK => clk, RN => rst_BAR, 
                           Q => n24135, QN => n_1050);
   clk_r_REG14285_S3 : DFFS_X1 port map( D => n1835, CK => clk, SN => rst_BAR, 
                           Q => n24134, QN => n_1051);
   clk_r_REG15112_S4 : DFFS_X1 port map( D => n25882, CK => clk, SN => rst_BAR,
                           Q => n24132, QN => n_1052);
   clk_r_REG14008_S4 : DFFS_X1 port map( D => n1829, CK => clk, SN => n25890, Q
                           => n24131, QN => n_1053);
   clk_r_REG13792_S4 : DFFR_X1 port map( D => n1833, CK => clk, RN => rst_BAR, 
                           Q => n24126, QN => n_1054);
   clk_r_REG14273_S3 : DFFS_X1 port map( D => n1818, CK => clk, SN => rst_BAR, 
                           Q => n24125, QN => n_1055);
   clk_r_REG14267_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => rst_BAR, 
                           Q => n24124, QN => n_1056);
   clk_r_REG14226_S3 : DFFR_X1 port map( D => n25870, CK => clk, RN => rst_BAR,
                           Q => n24123, QN => n27676);
   clk_r_REG14166_S3 : DFFR_X1 port map( D => n25865, CK => clk, RN => rst_BAR,
                           Q => n24122, QN => n27706);
   clk_r_REG14167_S3 : DFFS_X1 port map( D => n25865, CK => clk, SN => rst_BAR,
                           Q => n24121, QN => n_1057);
   clk_r_REG13866_S10 : DFFR_X1 port map( D => n1824, CK => clk, RN => rst_BAR,
                           Q => n24120, QN => n_1058);
   clk_r_REG14276_S3 : DFFR_X1 port map( D => n1828, CK => clk, RN => rst_BAR, 
                           Q => n24119, QN => n_1059);
   clk_r_REG14297_S3 : DFFR_X1 port map( D => n1819, CK => clk, RN => rst_BAR, 
                           Q => n24118, QN => n_1060);
   clk_r_REG14098_S4 : DFFR_X1 port map( D => n1822, CK => clk, RN => rst_BAR, 
                           Q => n24117, QN => n_1061);
   clk_r_REG14110_S4 : DFFR_X1 port map( D => n1821, CK => clk, RN => rst_BAR, 
                           Q => n24116, QN => n_1062);
   clk_r_REG14294_S4 : DFFR_X1 port map( D => n1827, CK => clk, RN => rst_BAR, 
                           Q => n24115, QN => n_1063);
   clk_r_REG13784_S5 : DFFS_X1 port map( D => n1787, CK => clk, SN => rst_BAR, 
                           Q => n24114, QN => n_1064);
   clk_r_REG14222_S3 : DFFR_X1 port map( D => n1868, CK => clk, RN => rst_BAR, 
                           Q => n24113, QN => n_1065);
   clk_r_REG14190_S3 : DFFS_X1 port map( D => n1864, CK => clk, SN => rst_BAR, 
                           Q => n24112, QN => n_1066);
   clk_r_REG14194_S3 : DFFS_X1 port map( D => n1870, CK => clk, SN => rst_BAR, 
                           Q => n24111, QN => n_1067);
   clk_r_REG14201_S3 : DFFS_X1 port map( D => n25866, CK => clk, SN => rst_BAR,
                           Q => n24110, QN => n_1068);
   clk_r_REG14146_S4 : DFFR_X1 port map( D => n25886, CK => clk, RN => rst_BAR,
                           Q => n24109, QN => n_1069);
   clk_r_REG14180_S3 : DFFS_X1 port map( D => n25859, CK => clk, SN => rst_BAR,
                           Q => n24108, QN => n27683);
   clk_r_REG14250_S3 : DFFR_X1 port map( D => n1894, CK => clk, RN => rst_BAR, 
                           Q => n24107, QN => n27691);
   clk_r_REG14253_S3 : DFFS_X1 port map( D => n1860, CK => clk, SN => rst_BAR, 
                           Q => n24106, QN => n_1070);
   clk_r_REG14324_S3 : DFFR_X1 port map( D => n1862, CK => clk, RN => rst_BAR, 
                           Q => n24105, QN => n27673);
   clk_r_REG14176_S3 : DFFR_X1 port map( D => n25873, CK => clk, RN => rst_BAR,
                           Q => n24104, QN => n27678);
   clk_r_REG14204_S3 : DFFR_X1 port map( D => n25875, CK => clk, RN => rst_BAR,
                           Q => n24103, QN => n_1071);
   clk_r_REG14046_S5 : DFFR_X1 port map( D => n1811, CK => clk, RN => rst_BAR, 
                           Q => n24102, QN => n_1072);
   clk_r_REG14334_S3 : DFFR_X1 port map( D => n1858, CK => clk, RN => rst_BAR, 
                           Q => n24101, QN => n_1073);
   clk_r_REG14037_S5 : DFFS_X1 port map( D => n25881, CK => clk, SN => rst_BAR,
                           Q => n24100, QN => n_1074);
   clk_r_REG14197_S3 : DFFR_X1 port map( D => n25874, CK => clk, RN => rst_BAR,
                           Q => n24099, QN => n_1075);
   clk_r_REG14216_S3 : DFFR_X1 port map( D => n25868, CK => clk, RN => rst_BAR,
                           Q => n24098, QN => n_1076);
   clk_r_REG14322_S3 : DFFR_X1 port map( D => n25879, CK => clk, RN => n25889, 
                           Q => n24097, QN => n27671);
   clk_r_REG14218_S3 : DFFS_X1 port map( D => n25876, CK => clk, SN => rst_BAR,
                           Q => n24096, QN => n_1077);
   clk_r_REG14183_S3 : DFFR_X1 port map( D => n25871, CK => clk, RN => rst_BAR,
                           Q => n24095, QN => n_1078);
   clk_r_REG14184_S3 : DFFS_X1 port map( D => n25871, CK => clk, SN => rst_BAR,
                           Q => n24094, QN => n_1079);
   clk_r_REG14173_S3 : DFFR_X1 port map( D => n25867, CK => clk, RN => rst_BAR,
                           Q => n24093, QN => n_1080);
   clk_r_REG14172_S3 : DFFS_X1 port map( D => n25867, CK => clk, SN => rst_BAR,
                           Q => n24092, QN => n_1081);
   clk_r_REG14206_S3 : DFFR_X1 port map( D => n25869, CK => clk, RN => rst_BAR,
                           Q => n24091, QN => n27702);
   clk_r_REG14188_S3 : DFFR_X1 port map( D => n1866, CK => clk, RN => rst_BAR, 
                           Q => n24090, QN => n_1082);
   clk_r_REG14187_S3 : DFFS_X1 port map( D => n1866, CK => clk, SN => rst_BAR, 
                           Q => n24089, QN => n27677);
   clk_r_REG15180_S5 : DFFR_X1 port map( D => n25888, CK => clk, RN => rst_BAR,
                           Q => n24088, QN => n_1083);
   clk_r_REG14090_S4 : DFFR_X1 port map( D => n21556, CK => clk, RN => rst_BAR,
                           Q => n24087, QN => n_1084);
   clk_r_REG14619_S3 : DFFR_X1 port map( D => n1831, CK => clk, RN => n25890, Q
                           => n24086, QN => n_1085);
   clk_r_REG14621_S3 : DFFR_X1 port map( D => n1830, CK => clk, RN => rst_BAR, 
                           Q => n24085, QN => n_1086);
   clk_r_REG14210_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, 
                           Q => n24084, QN => n_1087);
   clk_r_REG14211_S3 : DFFS_X1 port map( D => n1869, CK => clk, SN => rst_BAR, 
                           Q => n24083, QN => n_1088);
   clk_r_REG14316_S3 : DFFR_X1 port map( D => n1865, CK => clk, RN => rst_BAR, 
                           Q => n24082, QN => n27681);
   clk_r_REG14335_S3 : DFFR_X1 port map( D => n1863, CK => clk, RN => rst_BAR, 
                           Q => n24081, QN => n27670);
   clk_r_REG14336_S3 : DFFS_X1 port map( D => n1863, CK => clk, SN => rst_BAR, 
                           Q => n24080, QN => n27663);
   clk_r_REG14126_S4 : DFFS_X1 port map( D => n25884, CK => clk, SN => rst_BAR,
                           Q => n24079, QN => n_1089);
   clk_r_REG16455_S4 : DFFS_X1 port map( D => n1808, CK => clk, SN => rst_BAR, 
                           Q => n_1090, QN => n25872);
   clk_r_REG14440_S6 : DFFS_X1 port map( D => n1851, CK => clk, SN => rst_BAR, 
                           Q => n24077, QN => n_1091);
   clk_r_REG16595_S5 : DFFS_X1 port map( D => n1855, CK => clk, SN => rst_BAR, 
                           Q => n24076, QN => n_1092);
   clk_r_REG14317_S3 : DFFR_X1 port map( D => n1865, CK => clk, RN => rst_BAR, 
                           Q => n24075, QN => n_1093);
   clk_r_REG14195_S3 : DFFS_X1 port map( D => n1870, CK => clk, SN => rst_BAR, 
                           Q => n24074, QN => n_1094);
   clk_r_REG14212_S3 : DFFS_X1 port map( D => n1869, CK => clk, SN => rst_BAR, 
                           Q => n24073, QN => n_1095);
   clk_r_REG14223_S3 : DFFR_X1 port map( D => n1868, CK => clk, RN => rst_BAR, 
                           Q => n24072, QN => n_1096);
   clk_r_REG14202_S3 : DFFR_X1 port map( D => n25866, CK => clk, RN => rst_BAR,
                           Q => n24071, QN => n_1097);
   clk_r_REG14200_S3 : DFFS_X1 port map( D => n25866, CK => clk, SN => n25890, 
                           Q => n24070, QN => n_1098);
   clk_r_REG14177_S3 : DFFR_X1 port map( D => n25873, CK => clk, RN => rst_BAR,
                           Q => n24069, QN => n_1099);
   clk_r_REG14215_S3 : DFFR_X1 port map( D => n25868, CK => clk, RN => rst_BAR,
                           Q => n24068, QN => n_1100);
   clk_r_REG14325_S3 : DFFR_X1 port map( D => n1862, CK => clk, RN => rst_BAR, 
                           Q => n24067, QN => n_1101);
   clk_r_REG14171_S3 : DFFR_X1 port map( D => n25867, CK => clk, RN => rst_BAR,
                           Q => n24066, QN => n27686);
   clk_r_REG14213_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, 
                           Q => n24065, QN => n_1102);
   clk_r_REG14192_S3 : DFFS_X1 port map( D => n1864, CK => clk, SN => rst_BAR, 
                           Q => n24064, QN => n_1103);
   clk_r_REG14168_S3 : DFFS_X1 port map( D => n25865, CK => clk, SN => n25890, 
                           Q => n24063, QN => n27708);
   clk_r_REG14179_S3 : DFFS_X1 port map( D => n25859, CK => clk, SN => rst_BAR,
                           Q => n24062, QN => n_1104);
   clk_r_REG14225_S3 : DFFR_X1 port map( D => n25870, CK => clk, RN => rst_BAR,
                           Q => n24061, QN => n_1105);
   clk_r_REG14331_S3 : DFFR_X1 port map( D => n1843, CK => clk, RN => rst_BAR, 
                           Q => n24060, QN => n27689);
   clk_r_REG14251_S3 : DFFR_X1 port map( D => n1859, CK => clk, RN => rst_BAR, 
                           Q => n_1106, QN => n27699);
   clk_r_REG14241_S3 : DFFR_X1 port map( D => n1861, CK => clk, RN => rst_BAR, 
                           Q => n24058, QN => n_1107);
   clk_r_REG14252_S3 : DFFR_X1 port map( D => n1836, CK => clk, RN => rst_BAR, 
                           Q => n24057, QN => n_1108);
   clk_r_REG16585_S6 : DFFS_X1 port map( D => n1852, CK => clk, SN => rst_BAR, 
                           Q => n24056, QN => n_1109);
   clk_r_REG14441_S6 : DFFS_X1 port map( D => n1851, CK => clk, SN => rst_BAR, 
                           Q => n24055, QN => n_1110);
   clk_r_REG14339_S3 : DFFS_X1 port map( D => n1853, CK => clk, SN => rst_BAR, 
                           Q => n24054, QN => n_1111);
   clk_r_REG16596_S5 : DFFS_X1 port map( D => n1855, CK => clk, SN => rst_BAR, 
                           Q => n24053, QN => n_1112);
   clk_r_REG14979_S3 : DFFS_X1 port map( D => n1854, CK => clk, SN => rst_BAR, 
                           Q => n24052, QN => n_1113);
   clk_r_REG14323_S3 : DFFR_X1 port map( D => n1841, CK => clk, RN => rst_BAR, 
                           Q => n24051, QN => n_1114);
   clk_r_REG16738_S2 : DFFS_X1 port map( D => n1871, CK => clk, SN => rst_BAR, 
                           Q => n24050, QN => n_1115);
   clk_r_REG14838_S3 : DFFR_X1 port map( D => DATA1(2), CK => clk, RN => 
                           rst_BAR, Q => n24049, QN => n_1116);
   clk_r_REG14698_S3 : DFFR_X1 port map( D => DATA1(3), CK => clk, RN => 
                           rst_BAR, Q => n24048, QN => n27682);
   clk_r_REG14095_S3 : DFFS_X1 port map( D => n1850, CK => clk, SN => rst_BAR, 
                           Q => n24047, QN => n27704);
   clk_r_REG14059_S3 : DFFS_X1 port map( D => n1849, CK => clk, SN => rst_BAR, 
                           Q => n24046, QN => n_1117);
   clk_r_REG13922_S4 : DFFR_X1 port map( D => n22975, CK => clk, RN => rst_BAR,
                           Q => n27700, QN => n25858);
   clk_r_REG13692_S4 : DFFR_X1 port map( D => n19294, CK => clk, RN => rst_BAR,
                           Q => n24044, QN => n_1118);
   clk_r_REG14328_S3 : DFFS_X1 port map( D => n1856, CK => clk, SN => rst_BAR, 
                           Q => n_1119, QN => n24041);
   clk_r_REG14327_S3 : DFFR_X1 port map( D => n1856, CK => clk, RN => rst_BAR, 
                           Q => n_1120, QN => n24040);
   clk_r_REG14220_S3 : DFFR_X1 port map( D => n1863, CK => clk, RN => rst_BAR, 
                           Q => n_1121, QN => n24039);
   clk_r_REG14219_S3 : DFFS_X1 port map( D => n1863, CK => clk, SN => rst_BAR, 
                           Q => n27696, QN => n24038);
   clk_r_REG14620_S3 : DFFR_X1 port map( D => n1830, CK => clk, RN => rst_BAR, 
                           Q => n27703, QN => n24036);
   clk_r_REG14209_S3 : DFFS_X1 port map( D => n19271, CK => clk, SN => rst_BAR,
                           Q => n24035, QN => n_1122);
   clk_r_REG14315_S3 : DFFR_X1 port map( D => n1865, CK => clk, RN => rst_BAR, 
                           Q => n27665, QN => n24034);
   clk_r_REG14191_S3 : DFFR_X1 port map( D => n19261, CK => clk, RN => rst_BAR,
                           Q => n24033, QN => n_1123);
   clk_r_REG16739_S3 : DFFR_X1 port map( D => n1825, CK => clk, RN => rst_BAR, 
                           Q => n_1124, QN => n24032);
   clk_r_REG14151_S4 : DFFS_X1 port map( D => n19270, CK => clk, SN => rst_BAR,
                           Q => n24031, QN => n_1125);
   clk_r_REG14564_S4 : DFFS_X1 port map( D => n1809, CK => clk, SN => rst_BAR, 
                           Q => n24030, QN => n_1126);
   clk_r_REG14156_S3 : DFFR_X1 port map( D => n1831, CK => clk, RN => rst_BAR, 
                           Q => n27701, QN => n24029);
   clk_r_REG13769_S5 : DFFS_X1 port map( D => n19283, CK => clk, SN => rst_BAR,
                           Q => n24028, QN => n_1127);
   clk_r_REG14087_S4 : DFFS_X1 port map( D => n19278, CK => clk, SN => rst_BAR,
                           Q => n24026, QN => n_1128);
   clk_r_REG13800_S4 : DFFR_X1 port map( D => n19277, CK => clk, RN => n25889, 
                           Q => n24025, QN => n_1129);
   clk_r_REG14024_S5 : DFFR_X1 port map( D => n19272, CK => clk, RN => rst_BAR,
                           Q => n24024, QN => n_1130);
   clk_r_REG14025_S6 : DFFR_X1 port map( D => n24024, CK => clk, RN => rst_BAR,
                           Q => n24023, QN => n_1131);
   clk_r_REG14026_S7 : DFFR_X1 port map( D => n24023, CK => clk, RN => rst_BAR,
                           Q => n24022, QN => n_1132);
   clk_r_REG14027_S8 : DFFR_X1 port map( D => n24022, CK => clk, RN => rst_BAR,
                           Q => n24021, QN => n_1133);
   clk_r_REG14028_S9 : DFFR_X1 port map( D => n24021, CK => clk, RN => rst_BAR,
                           Q => n24020, QN => n_1134);
   clk_r_REG14092_S4 : DFFS_X1 port map( D => n1789, CK => clk, SN => rst_BAR, 
                           Q => n_1135, QN => n24019);
   clk_r_REG14693_S4 : DFFS_X1 port map( D => n19269, CK => clk, SN => rst_BAR,
                           Q => n24018, QN => n_1136);
   clk_r_REG14308_S4 : DFFS_X1 port map( D => n19267, CK => clk, SN => rst_BAR,
                           Q => n24017, QN => n_1137);
   clk_r_REG13746_S4 : DFFS_X1 port map( D => n19266, CK => clk, SN => rst_BAR,
                           Q => n24016, QN => n_1138);
   clk_r_REG13943_S10 : DFFS_X1 port map( D => n19265, CK => clk, SN => rst_BAR
                           , Q => n24015, QN => n_1139);
   clk_r_REG14051_S5 : DFFS_X1 port map( D => n17503, CK => clk, SN => rst_BAR,
                           Q => n24014, QN => n_1140);
   clk_r_REG14319_S3 : DFFS_X1 port map( D => n19262, CK => clk, SN => rst_BAR,
                           Q => n24013, QN => n_1141);
   clk_r_REG14154_S3 : DFFS_X1 port map( D => n8626, CK => clk, SN => n25890, Q
                           => n24012, QN => n_1142);
   clk_r_REG14155_S3 : DFFS_X1 port map( D => n19259, CK => clk, SN => rst_BAR,
                           Q => n24011, QN => n_1143);
   clk_r_REG13640_S4 : DFFR_X1 port map( D => n19253, CK => clk, RN => rst_BAR,
                           Q => n24010, QN => n_1144);
   clk_r_REG13641_S5 : DFFR_X1 port map( D => n24010, CK => clk, RN => rst_BAR,
                           Q => n24009, QN => n_1145);
   clk_r_REG13642_S6 : DFFR_X1 port map( D => n24009, CK => clk, RN => rst_BAR,
                           Q => n24008, QN => n_1146);
   clk_r_REG13643_S7 : DFFR_X1 port map( D => n24008, CK => clk, RN => rst_BAR,
                           Q => n24007, QN => n_1147);
   clk_r_REG13644_S8 : DFFR_X1 port map( D => n24007, CK => clk, RN => rst_BAR,
                           Q => n24006, QN => n_1148);
   clk_r_REG13645_S9 : DFFR_X1 port map( D => n24006, CK => clk, RN => rst_BAR,
                           Q => n24005, QN => n_1149);
   clk_r_REG14147_S4 : DFFS_X1 port map( D => n19252, CK => clk, SN => rst_BAR,
                           Q => n24004, QN => n_1150);
   clk_r_REG13874_S5 : DFFS_X1 port map( D => n19248, CK => clk, SN => n25890, 
                           Q => n23999, QN => n_1151);
   clk_r_REG13678_S4 : DFFR_X1 port map( D => n25883, CK => clk, RN => rst_BAR,
                           Q => n_1152, QN => n23998);
   clk_r_REG13978_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_16_port, CK => clk, 
                           RN => rst_BAR, Q => n23997, QN => n_1153);
   clk_r_REG13972_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_17_port, CK => clk, 
                           RN => rst_BAR, Q => n23996, QN => n_1154);
   clk_r_REG13967_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_18_port, CK => clk, 
                           RN => rst_BAR, Q => n23995, QN => n_1155);
   clk_r_REG13961_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_19_port, CK => clk, 
                           RN => rst_BAR, Q => n23994, QN => n_1156);
   clk_r_REG13956_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_20_port, CK => clk, 
                           RN => rst_BAR, Q => n23993, QN => n_1157);
   clk_r_REG13950_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_21_port, CK => clk, 
                           RN => rst_BAR, Q => n23992, QN => n_1158);
   clk_r_REG13944_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_22_port, CK => clk, 
                           RN => n25889, Q => n23991, QN => n_1159);
   clk_r_REG13938_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_23_port, CK => clk, 
                           RN => rst_BAR, Q => n23990, QN => n_1160);
   clk_r_REG13933_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_24_port, CK => clk, 
                           RN => rst_BAR, Q => n23989, QN => n_1161);
   clk_r_REG13928_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_25_port, CK => clk, 
                           RN => rst_BAR, Q => n23988, QN => n_1162);
   clk_r_REG13927_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_26_port, CK => clk, 
                           RN => rst_BAR, Q => n23987, QN => n_1163);
   clk_r_REG13926_S5 : DFFR_X1 port map( D => n19234, CK => clk, RN => rst_BAR,
                           Q => n23986, QN => n_1164);
   clk_r_REG13925_S5 : DFFR_X1 port map( D => n19233, CK => clk, RN => rst_BAR,
                           Q => n23985, QN => n_1165);
   clk_r_REG13923_S5 : DFFR_X1 port map( D => n19232, CK => clk, RN => rst_BAR,
                           Q => n23984, QN => n_1166);
   clk_r_REG13924_S6 : DFFR_X1 port map( D => n23984, CK => clk, RN => rst_BAR,
                           Q => n23983, QN => n_1167);
   clk_r_REG13694_S5 : DFFR_X1 port map( D => n19231, CK => clk, RN => n25889, 
                           Q => n23982, QN => n_1168);
   clk_r_REG13695_S6 : DFFR_X1 port map( D => n23982, CK => clk, RN => rst_BAR,
                           Q => n23981, QN => n_1169);
   clk_r_REG14692_S4 : DFFR_X1 port map( D => n19147, CK => clk, RN => rst_BAR,
                           Q => n23980, QN => n_1170);
   clk_r_REG13854_S5 : DFFR_X1 port map( D => n25887, CK => clk, RN => rst_BAR,
                           Q => n_1171, QN => n23978);
   clk_r_REG14217_S3 : DFFS_X1 port map( D => n25876, CK => clk, SN => n25890, 
                           Q => n_1172, QN => n23977);
   clk_r_REG14214_S3 : DFFR_X1 port map( D => n25868, CK => clk, RN => rst_BAR,
                           Q => n27707, QN => n23976);
   clk_r_REG14203_S3 : DFFR_X1 port map( D => n25875, CK => clk, RN => rst_BAR,
                           Q => n_1173, QN => n23975);
   clk_r_REG14145_S4 : DFFR_X1 port map( D => n25886, CK => clk, RN => rst_BAR,
                           Q => n_1174, QN => n23974);
   clk_r_REG14083_S4 : DFFR_X1 port map( D => n25885, CK => clk, RN => n25889, 
                           Q => n_1175, QN => n23973);
   clk_r_REG14199_S3 : DFFR_X1 port map( D => n25866, CK => clk, RN => rst_BAR,
                           Q => n_1176, QN => n23971);
   clk_r_REG14198_S3 : DFFS_X1 port map( D => n25866, CK => clk, SN => rst_BAR,
                           Q => n_1177, QN => n23970);
   clk_r_REG14150_S4 : DFFR_X1 port map( D => n1813, CK => clk, RN => rst_BAR, 
                           Q => n_1178, QN => n23969);
   clk_r_REG15245_S5 : DFFS_X1 port map( D => n17932, CK => clk, SN => rst_BAR,
                           Q => n23968, QN => n_1179);
   clk_r_REG14318_S3 : DFFR_X1 port map( D => n1862, CK => clk, RN => n25889, Q
                           => n_1180, QN => n23967);
   clk_r_REG14208_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, 
                           Q => n_1181, QN => n23966);
   clk_r_REG14207_S3 : DFFS_X1 port map( D => n1869, CK => clk, SN => rst_BAR, 
                           Q => n_1182, QN => n23965);
   clk_r_REG14186_S3 : DFFR_X1 port map( D => n1866, CK => clk, RN => rst_BAR, 
                           Q => n_1183, QN => n23964);
   clk_r_REG14185_S3 : DFFS_X1 port map( D => n1866, CK => clk, SN => rst_BAR, 
                           Q => n27664, QN => n23963);
   clk_r_REG14189_S3 : DFFS_X1 port map( D => n1864, CK => clk, SN => rst_BAR, 
                           Q => n27674, QN => n23962);
   clk_r_REG14174_S4 : DFFS_X1 port map( D => n1429, CK => clk, SN => rst_BAR, 
                           Q => n23961, QN => n_1184);
   clk_r_REG14048_S5 : DFFS_X1 port map( D => n21635, CK => clk, SN => rst_BAR,
                           Q => n23960, QN => n_1185);
   clk_r_REG13783_S5 : DFFR_X1 port map( D => n1815, CK => clk, RN => rst_BAR, 
                           Q => n_1186, QN => n23959);
   clk_r_REG14228_S3 : DFFR_X1 port map( D => n1860, CK => clk, RN => rst_BAR, 
                           Q => n_1187, QN => n23958);
   clk_r_REG14227_S3 : DFFS_X1 port map( D => n1860, CK => clk, SN => rst_BAR, 
                           Q => n27687, QN => n23957);
   clk_r_REG14246_S3 : DFFR_X1 port map( D => n1859, CK => clk, RN => rst_BAR, 
                           Q => n_1188, QN => n23956);
   clk_r_REG14245_S3 : DFFS_X1 port map( D => n1859, CK => clk, SN => n25890, Q
                           => n27688, QN => n23955);
   clk_r_REG14231_S3 : DFFS_X1 port map( D => n1861, CK => clk, SN => rst_BAR, 
                           Q => n27693, QN => n23953);
   clk_r_REG14044_S5 : DFFR_X1 port map( D => n1811, CK => clk, RN => rst_BAR, 
                           Q => n_1189, QN => n23952);
   clk_r_REG14498_S8 : DFFR_X1 port map( D => n19202, CK => clk, RN => rst_BAR,
                           Q => n23951, QN => n_1190);
   clk_r_REG14148_S4 : DFFS_X1 port map( D => n2808, CK => clk, SN => n25890, Q
                           => n23950, QN => n_1191);
   clk_r_REG15110_S4 : DFFS_X1 port map( D => n22765, CK => clk, SN => rst_BAR,
                           Q => n23948, QN => n_1192);
   clk_r_REG13897_S5 : DFFR_X1 port map( D => n18861, CK => clk, RN => rst_BAR,
                           Q => n23947, QN => n_1193);
   clk_r_REG13898_S6 : DFFR_X1 port map( D => n23947, CK => clk, RN => rst_BAR,
                           Q => n23946, QN => n_1194);
   clk_r_REG13899_S7 : DFFR_X1 port map( D => n23946, CK => clk, RN => rst_BAR,
                           Q => n23945, QN => n_1195);
   clk_r_REG13900_S8 : DFFR_X1 port map( D => n23945, CK => clk, RN => rst_BAR,
                           Q => n23944, QN => n_1196);
   clk_r_REG13901_S9 : DFFR_X1 port map( D => n23944, CK => clk, RN => rst_BAR,
                           Q => n23943, QN => n_1197);
   clk_r_REG13902_S10 : DFFS_X1 port map( D => n23943, CK => clk, SN => rst_BAR
                           , Q => n23942, QN => n_1198);
   clk_r_REG14829_S4 : DFFR_X1 port map( D => n19187, CK => clk, RN => rst_BAR,
                           Q => n23941, QN => n_1199);
   clk_r_REG14830_S5 : DFFR_X1 port map( D => n23941, CK => clk, RN => rst_BAR,
                           Q => n23940, QN => n_1200);
   clk_r_REG14831_S6 : DFFR_X1 port map( D => n23940, CK => clk, RN => rst_BAR,
                           Q => n23939, QN => n_1201);
   clk_r_REG14832_S7 : DFFR_X1 port map( D => n23939, CK => clk, RN => rst_BAR,
                           Q => n23938, QN => n_1202);
   clk_r_REG14833_S8 : DFFR_X1 port map( D => n23938, CK => clk, RN => rst_BAR,
                           Q => n23937, QN => n_1203);
   clk_r_REG14834_S9 : DFFR_X1 port map( D => n23937, CK => clk, RN => rst_BAR,
                           Q => n23936, QN => n_1204);
   clk_r_REG14099_S4 : DFFS_X1 port map( D => n19186, CK => clk, SN => rst_BAR,
                           Q => n23935, QN => n_1205);
   clk_r_REG14056_S4 : DFFR_X1 port map( D => n21634, CK => clk, RN => rst_BAR,
                           Q => n23934, QN => n_1206);
   clk_r_REG14091_S3 : DFFS_X1 port map( D => n18976, CK => clk, SN => n25890, 
                           Q => n23933, QN => n_1207);
   clk_r_REG14076_S10 : DFFS_X1 port map( D => n19184, CK => clk, SN => rst_BAR
                           , Q => n23932, QN => n_1208);
   clk_r_REG14114_S4 : DFFR_X1 port map( D => n22526, CK => clk, RN => rst_BAR,
                           Q => n23931, QN => n_1209);
   clk_r_REG14256_S3 : DFFR_X1 port map( D => n19183, CK => clk, RN => rst_BAR,
                           Q => n23930, QN => n_1210);
   clk_r_REG13786_S5 : DFFR_X1 port map( D => n19182, CK => clk, RN => rst_BAR,
                           Q => n23929, QN => n_1211);
   clk_r_REG13785_S5 : DFFS_X1 port map( D => n19268, CK => clk, SN => rst_BAR,
                           Q => n23928, QN => n_1212);
   clk_r_REG13776_S4 : DFFR_X1 port map( D => n19181, CK => clk, RN => n25889, 
                           Q => n23927, QN => n_1213);
   clk_r_REG14254_S4 : DFFS_X1 port map( D => n19180, CK => clk, SN => rst_BAR,
                           Q => n23926, QN => n_1214);
   clk_r_REG13747_S5 : DFFS_X1 port map( D => n19178, CK => clk, SN => rst_BAR,
                           Q => n23925, QN => n_1215);
   clk_r_REG16072_S3 : DFFS_X1 port map( D => n19176, CK => clk, SN => rst_BAR,
                           Q => n23924, QN => n_1216);
   clk_r_REG13725_S4 : DFFR_X1 port map( D => n19175, CK => clk, RN => rst_BAR,
                           Q => n23923, QN => n_1217);
   clk_r_REG14278_S4 : DFFR_X1 port map( D => n19174, CK => clk, RN => rst_BAR,
                           Q => n23922, QN => n_1218);
   clk_r_REG13718_S4 : DFFS_X1 port map( D => n12313, CK => clk, SN => rst_BAR,
                           Q => n_1219, QN => n25880);
   clk_r_REG14314_S3 : DFFR_X1 port map( D => n19171, CK => clk, RN => rst_BAR,
                           Q => n23920, QN => n_1220);
   clk_r_REG14312_S3 : DFFS_X1 port map( D => n19170, CK => clk, SN => rst_BAR,
                           Q => n23919, QN => n_1221);
   clk_r_REG13815_S4 : DFFR_X1 port map( D => n18917, CK => clk, RN => rst_BAR,
                           Q => n23918, QN => n_1222);
   clk_r_REG13966_S10 : DFFR_X1 port map( D => n19264, CK => clk, RN => n25889,
                           Q => n23917, QN => n_1223);
   clk_r_REG14579_S3 : DFFS_X1 port map( D => n19169, CK => clk, SN => rst_BAR,
                           Q => n23916, QN => n_1224);
   clk_r_REG14053_S5 : DFFR_X1 port map( D => n19168, CK => clk, RN => rst_BAR,
                           Q => n23915, QN => n_1225);
   clk_r_REG13693_S5 : DFFS_X1 port map( D => n22802, CK => clk, SN => rst_BAR,
                           Q => n23914, QN => n_1226);
   clk_r_REG13671_S11 : DFFS_X1 port map( D => n22281, CK => clk, SN => rst_BAR
                           , Q => n23913, QN => n_1227);
   clk_r_REG14050_S5 : DFFR_X1 port map( D => n19165, CK => clk, RN => rst_BAR,
                           Q => n23912, QN => n_1228);
   clk_r_REG14085_S5 : DFFR_X1 port map( D => n19163, CK => clk, RN => rst_BAR,
                           Q => n23911, QN => n_1229);
   clk_r_REG14086_S5 : DFFR_X1 port map( D => n19162, CK => clk, RN => rst_BAR,
                           Q => n23910, QN => n_1230);
   clk_r_REG14006_S5 : DFFR_X1 port map( D => n19161, CK => clk, RN => rst_BAR,
                           Q => n23909, QN => n_1231);
   clk_r_REG14350_S5 : DFFR_X1 port map( D => n19158, CK => clk, RN => n25890, 
                           Q => n23908, QN => n_1232);
   clk_r_REG14352_S6 : DFFR_X1 port map( D => n19157, CK => clk, RN => rst_BAR,
                           Q => n23907, QN => n_1233);
   clk_r_REG14354_S6 : DFFR_X1 port map( D => n19156, CK => clk, RN => rst_BAR,
                           Q => n23906, QN => n_1234);
   clk_r_REG14356_S6 : DFFR_X1 port map( D => n19155, CK => clk, RN => rst_BAR,
                           Q => n23905, QN => n_1235);
   clk_r_REG14358_S6 : DFFR_X1 port map( D => n19154, CK => clk, RN => rst_BAR,
                           Q => n23904, QN => n_1236);
   clk_r_REG14360_S6 : DFFR_X1 port map( D => n19153, CK => clk, RN => rst_BAR,
                           Q => n23903, QN => n_1237);
   clk_r_REG14362_S6 : DFFR_X1 port map( D => n19152, CK => clk, RN => rst_BAR,
                           Q => n23902, QN => n_1238);
   clk_r_REG14364_S6 : DFFR_X1 port map( D => n19151, CK => clk, RN => rst_BAR,
                           Q => n23901, QN => n_1239);
   clk_r_REG14366_S6 : DFFR_X1 port map( D => n19150, CK => clk, RN => rst_BAR,
                           Q => n23900, QN => n_1240);
   clk_r_REG14368_S6 : DFFR_X1 port map( D => n19149, CK => clk, RN => rst_BAR,
                           Q => n23899, QN => n_1241);
   clk_r_REG13989_S6 : DFFR_X1 port map( D => n19148, CK => clk, RN => rst_BAR,
                           Q => n23898, QN => n_1242);
   clk_r_REG14132_S10 : DFFS_X1 port map( D => n18882, CK => clk, SN => rst_BAR
                           , Q => n23896, QN => n_1243);
   clk_r_REG14182_S3 : DFFR_X1 port map( D => n25871, CK => clk, RN => rst_BAR,
                           Q => n27675, QN => n23895);
   clk_r_REG14181_S3 : DFFS_X1 port map( D => n25871, CK => clk, SN => rst_BAR,
                           Q => n27684, QN => n23894);
   clk_r_REG14196_S3 : DFFR_X1 port map( D => n25874, CK => clk, RN => n25890, 
                           Q => n_1244, QN => n23893);
   clk_r_REG14205_S3 : DFFR_X1 port map( D => n25869, CK => clk, RN => rst_BAR,
                           Q => n_1245, QN => n23892);
   clk_r_REG14175_S3 : DFFR_X1 port map( D => n25873, CK => clk, RN => rst_BAR,
                           Q => n27679, QN => n23891);
   clk_r_REG14124_S4 : DFFS_X1 port map( D => n19213, CK => clk, SN => rst_BAR,
                           Q => n23889, QN => n_1246);
   clk_r_REG14193_S3 : DFFS_X1 port map( D => n1870, CK => clk, SN => rst_BAR, 
                           Q => n27705, QN => n23888);
   clk_r_REG14221_S3 : DFFR_X1 port map( D => n1868, CK => clk, RN => rst_BAR, 
                           Q => n27661, QN => n23887);
   clk_r_REG13955_S10 : DFFR_X1 port map( D => n19433, CK => clk, RN => rst_BAR
                           , Q => n23886, QN => n_1247);
   clk_r_REG14685_S4 : DFFR_X1 port map( D => n19135, CK => clk, RN => rst_BAR,
                           Q => n23885, QN => n_1248);
   clk_r_REG14686_S5 : DFFR_X1 port map( D => n23885, CK => clk, RN => rst_BAR,
                           Q => n23884, QN => n_1249);
   clk_r_REG14687_S6 : DFFR_X1 port map( D => n23884, CK => clk, RN => rst_BAR,
                           Q => n23883, QN => n_1250);
   clk_r_REG14688_S7 : DFFR_X1 port map( D => n23883, CK => clk, RN => rst_BAR,
                           Q => n23882, QN => n_1251);
   clk_r_REG14689_S8 : DFFR_X1 port map( D => n23882, CK => clk, RN => rst_BAR,
                           Q => n23881, QN => n_1252);
   clk_r_REG14690_S9 : DFFR_X1 port map( D => n23881, CK => clk, RN => rst_BAR,
                           Q => n23880, QN => n_1253);
   clk_r_REG14343_S5 : DFFR_X1 port map( D => n19134, CK => clk, RN => rst_BAR,
                           Q => n23879, QN => n_1254);
   clk_r_REG14341_S4 : DFFR_X1 port map( D => n19133, CK => clk, RN => rst_BAR,
                           Q => n23878, QN => n_1255);
   clk_r_REG14070_S4 : DFFR_X1 port map( D => n19132, CK => clk, RN => rst_BAR,
                           Q => n23877, QN => n_1256);
   clk_r_REG14023_S4 : DFFR_X1 port map( D => n19131, CK => clk, RN => rst_BAR,
                           Q => n23876, QN => n_1257);
   clk_r_REG14022_S4 : DFFR_X1 port map( D => n19130, CK => clk, RN => rst_BAR,
                           Q => n23875, QN => n_1258);
   clk_r_REG14021_S4 : DFFR_X1 port map( D => n19129, CK => clk, RN => rst_BAR,
                           Q => n23874, QN => n_1259);
   clk_r_REG14020_S4 : DFFR_X1 port map( D => n19128, CK => clk, RN => rst_BAR,
                           Q => n23873, QN => n_1260);
   clk_r_REG14019_S4 : DFFR_X1 port map( D => n19127, CK => clk, RN => rst_BAR,
                           Q => n23872, QN => n_1261);
   clk_r_REG14018_S4 : DFFR_X1 port map( D => n19126, CK => clk, RN => rst_BAR,
                           Q => n23871, QN => n_1262);
   clk_r_REG14015_S4 : DFFR_X1 port map( D => n19125, CK => clk, RN => rst_BAR,
                           Q => n23870, QN => n_1263);
   clk_r_REG14004_S5 : DFFR_X1 port map( D => n19124, CK => clk, RN => rst_BAR,
                           Q => n23869, QN => n_1264);
   clk_r_REG13999_S5 : DFFR_X1 port map( D => n19123, CK => clk, RN => rst_BAR,
                           Q => n23868, QN => n_1265);
   clk_r_REG13996_S5 : DFFR_X1 port map( D => n19122, CK => clk, RN => rst_BAR,
                           Q => n23867, QN => n_1266);
   clk_r_REG13993_S5 : DFFR_X1 port map( D => n19121, CK => clk, RN => rst_BAR,
                           Q => n23866, QN => n_1267);
   clk_r_REG14133_S5 : DFFR_X1 port map( D => n19115, CK => clk, RN => rst_BAR,
                           Q => n23865, QN => n_1268);
   clk_r_REG14134_S6 : DFFR_X1 port map( D => n23865, CK => clk, RN => rst_BAR,
                           Q => n23864, QN => n_1269);
   clk_r_REG14135_S7 : DFFR_X1 port map( D => n23864, CK => clk, RN => rst_BAR,
                           Q => n23863, QN => n_1270);
   clk_r_REG14136_S8 : DFFR_X1 port map( D => n23863, CK => clk, RN => rst_BAR,
                           Q => n23862, QN => n_1271);
   clk_r_REG14137_S9 : DFFR_X1 port map( D => n23862, CK => clk, RN => n25889, 
                           Q => n23861, QN => n_1272);
   clk_r_REG13991_S5 : DFFR_X1 port map( D => n19113, CK => clk, RN => rst_BAR,
                           Q => n23860, QN => n_1273);
   clk_r_REG13992_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CK => clk, 
                           RN => rst_BAR, Q => n23859, QN => n_1274);
   clk_r_REG14071_S5 : DFFR_X1 port map( D => n19108, CK => clk, RN => rst_BAR,
                           Q => n23858, QN => n_1275);
   clk_r_REG14072_S6 : DFFR_X1 port map( D => n23858, CK => clk, RN => rst_BAR,
                           Q => n23857, QN => n_1276);
   clk_r_REG14073_S7 : DFFR_X1 port map( D => n23857, CK => clk, RN => rst_BAR,
                           Q => n23856, QN => n_1277);
   clk_r_REG14074_S8 : DFFR_X1 port map( D => n23856, CK => clk, RN => rst_BAR,
                           Q => n23855, QN => n_1278);
   clk_r_REG14075_S9 : DFFR_X1 port map( D => n23855, CK => clk, RN => rst_BAR,
                           Q => n23854, QN => n_1279);
   clk_r_REG13997_S6 : DFFR_X1 port map( D => n19107, CK => clk, RN => rst_BAR,
                           Q => n23853, QN => n_1280);
   clk_r_REG13994_S6 : DFFR_X1 port map( D => n19106, CK => clk, RN => rst_BAR,
                           Q => n23852, QN => n_1281);
   clk_r_REG13995_S6 : DFFR_X1 port map( D => n19105, CK => clk, RN => n25889, 
                           Q => n23851, QN => n_1282);
   clk_r_REG13842_S5 : DFFR_X1 port map( D => n19100, CK => clk, RN => rst_BAR,
                           Q => n23850, QN => n_1283);
   clk_r_REG13843_S6 : DFFR_X1 port map( D => n23850, CK => clk, RN => rst_BAR,
                           Q => n23849, QN => n_1284);
   clk_r_REG13844_S7 : DFFR_X1 port map( D => n23849, CK => clk, RN => rst_BAR,
                           Q => n23848, QN => n_1285);
   clk_r_REG13845_S8 : DFFR_X1 port map( D => n23848, CK => clk, RN => n25889, 
                           Q => n23847, QN => n_1286);
   clk_r_REG13846_S9 : DFFR_X1 port map( D => n23847, CK => clk, RN => rst_BAR,
                           Q => n23846, QN => n_1287);
   clk_r_REG14005_S6 : DFFR_X1 port map( D => n19099, CK => clk, RN => rst_BAR,
                           Q => n23845, QN => n_1288);
   clk_r_REG14000_S6 : DFFR_X1 port map( D => n19098, CK => clk, RN => rst_BAR,
                           Q => n23844, QN => n_1289);
   clk_r_REG14001_S6 : DFFR_X1 port map( D => n19097, CK => clk, RN => rst_BAR,
                           Q => n23843, QN => n_1290);
   clk_r_REG13861_S5 : DFFR_X1 port map( D => n19092, CK => clk, RN => rst_BAR,
                           Q => n23842, QN => n_1291);
   clk_r_REG13862_S6 : DFFR_X1 port map( D => n23842, CK => clk, RN => rst_BAR,
                           Q => n23841, QN => n_1292);
   clk_r_REG13863_S7 : DFFR_X1 port map( D => n23841, CK => clk, RN => rst_BAR,
                           Q => n23840, QN => n_1293);
   clk_r_REG13864_S8 : DFFR_X1 port map( D => n23840, CK => clk, RN => rst_BAR,
                           Q => n23839, QN => n_1294);
   clk_r_REG13865_S9 : DFFR_X1 port map( D => n23839, CK => clk, RN => rst_BAR,
                           Q => n23838, QN => n_1295);
   clk_r_REG14016_S6 : DFFR_X1 port map( D => n19090, CK => clk, RN => rst_BAR,
                           Q => n23837, QN => n_1296);
   clk_r_REG14017_S6 : DFFR_X1 port map( D => n19089, CK => clk, RN => rst_BAR,
                           Q => n23836, QN => n_1297);
   clk_r_REG13665_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CK => clk, RN => rst_BAR, Q => n23835, QN => n_1298)
                           ;
   clk_r_REG13666_S6 : DFFR_X1 port map( D => n19085, CK => clk, RN => rst_BAR,
                           Q => n23834, QN => n_1299);
   clk_r_REG13667_S7 : DFFR_X1 port map( D => n23834, CK => clk, RN => rst_BAR,
                           Q => n23833, QN => n_1300);
   clk_r_REG13668_S8 : DFFR_X1 port map( D => n23833, CK => clk, RN => rst_BAR,
                           Q => n23832, QN => n_1301);
   clk_r_REG13669_S9 : DFFR_X1 port map( D => n23832, CK => clk, RN => rst_BAR,
                           Q => n23831, QN => n_1302);
   clk_r_REG13670_S10 : DFFR_X1 port map( D => n23831, CK => clk, RN => rst_BAR
                           , Q => n23830, QN => n_1303);
   clk_r_REG13893_S7 : DFFR_X1 port map( D => n19083, CK => clk, RN => rst_BAR,
                           Q => n23829, QN => n_1304);
   clk_r_REG13911_S6 : DFFR_X1 port map( D => n19079, CK => clk, RN => rst_BAR,
                           Q => n23828, QN => n_1305);
   clk_r_REG13912_S7 : DFFR_X1 port map( D => n23828, CK => clk, RN => n25889, 
                           Q => n23827, QN => n_1306);
   clk_r_REG13913_S8 : DFFR_X1 port map( D => n23827, CK => clk, RN => rst_BAR,
                           Q => n23826, QN => n_1307);
   clk_r_REG13914_S9 : DFFR_X1 port map( D => n23826, CK => clk, RN => rst_BAR,
                           Q => n23825, QN => n_1308);
   clk_r_REG13979_S6 : DFFR_X1 port map( D => n19075, CK => clk, RN => rst_BAR,
                           Q => n23824, QN => n_1309);
   clk_r_REG13980_S7 : DFFR_X1 port map( D => n23824, CK => clk, RN => rst_BAR,
                           Q => n23823, QN => n_1310);
   clk_r_REG13981_S8 : DFFR_X1 port map( D => n23823, CK => clk, RN => rst_BAR,
                           Q => n23822, QN => n_1311);
   clk_r_REG13982_S9 : DFFR_X1 port map( D => n23822, CK => clk, RN => rst_BAR,
                           Q => n23821, QN => n_1312);
   clk_r_REG13973_S6 : DFFR_X1 port map( D => n19071, CK => clk, RN => rst_BAR,
                           Q => n23820, QN => n_1313);
   clk_r_REG13974_S7 : DFFR_X1 port map( D => n23820, CK => clk, RN => rst_BAR,
                           Q => n23819, QN => n_1314);
   clk_r_REG13975_S8 : DFFR_X1 port map( D => n23819, CK => clk, RN => rst_BAR,
                           Q => n23818, QN => n_1315);
   clk_r_REG13976_S9 : DFFR_X1 port map( D => n23818, CK => clk, RN => rst_BAR,
                           Q => n23817, QN => n_1316);
   clk_r_REG13968_S6 : DFFR_X1 port map( D => n19067, CK => clk, RN => rst_BAR,
                           Q => n23816, QN => n_1317);
   clk_r_REG13969_S7 : DFFR_X1 port map( D => n23816, CK => clk, RN => rst_BAR,
                           Q => n23815, QN => n_1318);
   clk_r_REG13970_S8 : DFFR_X1 port map( D => n23815, CK => clk, RN => rst_BAR,
                           Q => n23814, QN => n_1319);
   clk_r_REG13971_S9 : DFFR_X1 port map( D => n23814, CK => clk, RN => rst_BAR,
                           Q => n23813, QN => n_1320);
   clk_r_REG13962_S6 : DFFR_X1 port map( D => n19063, CK => clk, RN => rst_BAR,
                           Q => n23812, QN => n_1321);
   clk_r_REG13963_S7 : DFFR_X1 port map( D => n23812, CK => clk, RN => rst_BAR,
                           Q => n23811, QN => n_1322);
   clk_r_REG13964_S8 : DFFR_X1 port map( D => n23811, CK => clk, RN => rst_BAR,
                           Q => n23810, QN => n_1323);
   clk_r_REG13965_S9 : DFFR_X1 port map( D => n23810, CK => clk, RN => rst_BAR,
                           Q => n23809, QN => n_1324);
   clk_r_REG13957_S6 : DFFR_X1 port map( D => n19059, CK => clk, RN => rst_BAR,
                           Q => n23808, QN => n_1325);
   clk_r_REG13958_S7 : DFFR_X1 port map( D => n23808, CK => clk, RN => rst_BAR,
                           Q => n23807, QN => n_1326);
   clk_r_REG13959_S8 : DFFR_X1 port map( D => n23807, CK => clk, RN => n25889, 
                           Q => n23806, QN => n_1327);
   clk_r_REG13960_S9 : DFFR_X1 port map( D => n23806, CK => clk, RN => rst_BAR,
                           Q => n23805, QN => n_1328);
   clk_r_REG13951_S6 : DFFR_X1 port map( D => n19055, CK => clk, RN => n25890, 
                           Q => n23804, QN => n_1329);
   clk_r_REG13952_S7 : DFFR_X1 port map( D => n23804, CK => clk, RN => rst_BAR,
                           Q => n23803, QN => n_1330);
   clk_r_REG13953_S8 : DFFR_X1 port map( D => n23803, CK => clk, RN => rst_BAR,
                           Q => n23802, QN => n_1331);
   clk_r_REG13954_S9 : DFFR_X1 port map( D => n23802, CK => clk, RN => rst_BAR,
                           Q => n23801, QN => n_1332);
   clk_r_REG13945_S6 : DFFR_X1 port map( D => n19051, CK => clk, RN => rst_BAR,
                           Q => n23800, QN => n_1333);
   clk_r_REG13946_S7 : DFFR_X1 port map( D => n23800, CK => clk, RN => rst_BAR,
                           Q => n23799, QN => n_1334);
   clk_r_REG13947_S8 : DFFR_X1 port map( D => n23799, CK => clk, RN => rst_BAR,
                           Q => n23798, QN => n_1335);
   clk_r_REG13948_S9 : DFFR_X1 port map( D => n23798, CK => clk, RN => rst_BAR,
                           Q => n23797, QN => n_1336);
   clk_r_REG13939_S6 : DFFR_X1 port map( D => n19047, CK => clk, RN => rst_BAR,
                           Q => n23796, QN => n_1337);
   clk_r_REG13940_S7 : DFFR_X1 port map( D => n23796, CK => clk, RN => rst_BAR,
                           Q => n23795, QN => n_1338);
   clk_r_REG13941_S8 : DFFR_X1 port map( D => n23795, CK => clk, RN => rst_BAR,
                           Q => n23794, QN => n_1339);
   clk_r_REG13942_S9 : DFFR_X1 port map( D => n23794, CK => clk, RN => rst_BAR,
                           Q => n23793, QN => n_1340);
   clk_r_REG13934_S6 : DFFR_X1 port map( D => n19042, CK => clk, RN => rst_BAR,
                           Q => n23792, QN => n_1341);
   clk_r_REG13935_S7 : DFFR_X1 port map( D => n23792, CK => clk, RN => rst_BAR,
                           Q => n23791, QN => n_1342);
   clk_r_REG13936_S8 : DFFR_X1 port map( D => n23791, CK => clk, RN => rst_BAR,
                           Q => n23790, QN => n_1343);
   clk_r_REG13937_S9 : DFFR_X1 port map( D => n23790, CK => clk, RN => rst_BAR,
                           Q => n23789, QN => n_1344);
   clk_r_REG13929_S6 : DFFR_X1 port map( D => n19038, CK => clk, RN => rst_BAR,
                           Q => n23788, QN => n_1345);
   clk_r_REG13930_S7 : DFFR_X1 port map( D => n23788, CK => clk, RN => rst_BAR,
                           Q => n23787, QN => n_1346);
   clk_r_REG13931_S8 : DFFR_X1 port map( D => n23787, CK => clk, RN => rst_BAR,
                           Q => n23786, QN => n_1347);
   clk_r_REG13932_S9 : DFFR_X1 port map( D => n23786, CK => clk, RN => rst_BAR,
                           Q => n23785, QN => n_1348);
   clk_r_REG13876_S7 : DFFR_X1 port map( D => n19033, CK => clk, RN => rst_BAR,
                           Q => n23784, QN => n_1349);
   clk_r_REG13877_S8 : DFFR_X1 port map( D => n23784, CK => clk, RN => n25889, 
                           Q => n23783, QN => n_1350);
   clk_r_REG13878_S9 : DFFR_X1 port map( D => n23783, CK => clk, RN => rst_BAR,
                           Q => n23782, QN => n_1351);
   clk_r_REG13879_S10 : DFFR_X1 port map( D => n23782, CK => clk, RN => rst_BAR
                           , Q => n23781, QN => n_1352);
   clk_r_REG13880_S7 : DFFR_X1 port map( D => n19030, CK => clk, RN => rst_BAR,
                           Q => n23780, QN => n_1353);
   clk_r_REG13881_S8 : DFFR_X1 port map( D => n23780, CK => clk, RN => rst_BAR,
                           Q => n23779, QN => n_1354);
   clk_r_REG13882_S9 : DFFR_X1 port map( D => n23779, CK => clk, RN => rst_BAR,
                           Q => n23778, QN => n_1355);
   clk_r_REG13883_S10 : DFFR_X1 port map( D => n23778, CK => clk, RN => rst_BAR
                           , Q => n23777, QN => n_1356);
   clk_r_REG13884_S7 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CK => clk, RN => rst_BAR, Q => n23776, QN => n_1357)
                           ;
   clk_r_REG13885_S7 : DFFR_X1 port map( D => n19027, CK => clk, RN => rst_BAR,
                           Q => n23775, QN => n_1358);
   clk_r_REG13886_S8 : DFFR_X1 port map( D => n23775, CK => clk, RN => rst_BAR,
                           Q => n23774, QN => n_1359);
   clk_r_REG13887_S9 : DFFR_X1 port map( D => n23774, CK => clk, RN => rst_BAR,
                           Q => n23773, QN => n_1360);
   clk_r_REG13888_S10 : DFFR_X1 port map( D => n23773, CK => clk, RN => rst_BAR
                           , Q => n23772, QN => n_1361);
   clk_r_REG13890_S8 : DFFR_X1 port map( D => n19024, CK => clk, RN => rst_BAR,
                           Q => n23771, QN => n_1362);
   clk_r_REG13891_S9 : DFFR_X1 port map( D => n23771, CK => clk, RN => rst_BAR,
                           Q => n23770, QN => n_1363);
   clk_r_REG13892_S10 : DFFR_X1 port map( D => n23770, CK => clk, RN => rst_BAR
                           , Q => n23769, QN => n_1364);
   clk_r_REG13696_S7 : DFFR_X1 port map( D => n19021, CK => clk, RN => rst_BAR,
                           Q => n23768, QN => n_1365);
   clk_r_REG13697_S8 : DFFR_X1 port map( D => n23768, CK => clk, RN => rst_BAR,
                           Q => n23767, QN => n_1366);
   clk_r_REG13698_S9 : DFFR_X1 port map( D => n23767, CK => clk, RN => rst_BAR,
                           Q => n23766, QN => n_1367);
   clk_r_REG13894_S7 : DFFR_X1 port map( D => n19018, CK => clk, RN => rst_BAR,
                           Q => n23765, QN => n_1368);
   clk_r_REG13895_S8 : DFFR_X1 port map( D => n23765, CK => clk, RN => rst_BAR,
                           Q => n23764, QN => n_1369);
   clk_r_REG13896_S9 : DFFR_X1 port map( D => n23764, CK => clk, RN => rst_BAR,
                           Q => n23763, QN => n_1370);
   clk_r_REG13656_S6 : DFFR_X1 port map( D => n19010, CK => clk, RN => rst_BAR,
                           Q => n23762, QN => n_1371);
   clk_r_REG14109_S4 : DFFR_X1 port map( D => n21296, CK => clk, RN => rst_BAR,
                           Q => n_1372, QN => n25863);
   clk_r_REG14275_S3 : DFFR_X1 port map( D => n1828, CK => clk, RN => n25889, Q
                           => n_1373, QN => n23760);
   clk_r_REG14274_S3 : DFFS_X1 port map( D => n1842, CK => clk, SN => n25890, Q
                           => n_1374, QN => n23759);
   clk_r_REG14300_S3 : DFFR_X1 port map( D => n1816, CK => clk, RN => rst_BAR, 
                           Q => n_1375, QN => n25878);
   clk_r_REG14299_S3 : DFFR_X1 port map( D => n21379, CK => clk, RN => rst_BAR,
                           Q => n23757, QN => n_1376);
   clk_r_REG14302_S3 : DFFR_X1 port map( D => n21378, CK => clk, RN => rst_BAR,
                           Q => n23756, QN => n_1377);
   clk_r_REG14271_S3 : DFFS_X1 port map( D => n1818, CK => clk, SN => rst_BAR, 
                           Q => n_1378, QN => n23755);
   clk_r_REG14298_S4 : DFFR_X1 port map( D => n19399, CK => clk, RN => rst_BAR,
                           Q => n27690, QN => n25877);
   clk_r_REG14268_S4 : DFFR_X1 port map( D => n1834, CK => clk, RN => rst_BAR, 
                           Q => n_1379, QN => n23753);
   clk_r_REG14295_S3 : DFFR_X1 port map( D => n1819, CK => clk, RN => n25889, Q
                           => n_1380, QN => n23752);
   clk_r_REG14102_S4 : DFFR_X1 port map( D => n1820, CK => clk, RN => rst_BAR, 
                           Q => n_1381, QN => n23751);
   clk_r_REG14265_S3 : DFFS_X1 port map( D => n1826, CK => clk, SN => rst_BAR, 
                           Q => n23750, QN => n_1382);
   clk_r_REG14292_S4 : DFFR_X1 port map( D => n1827, CK => clk, RN => rst_BAR, 
                           Q => n27697, QN => n23749);
   clk_r_REG14290_S3 : DFFR_X1 port map( D => n1838, CK => clk, RN => rst_BAR, 
                           Q => n27695, QN => n23748);
   clk_r_REG14289_S3 : DFFR_X1 port map( D => n21485, CK => clk, RN => rst_BAR,
                           Q => n23747, QN => n_1383);
   clk_r_REG14307_S3 : DFFR_X1 port map( D => n21484, CK => clk, RN => rst_BAR,
                           Q => n23746, QN => n_1384);
   clk_r_REG14288_S3 : DFFR_X1 port map( D => n21491, CK => clk, RN => rst_BAR,
                           Q => n23745, QN => n_1385);
   clk_r_REG14301_S3 : DFFR_X1 port map( D => n21490, CK => clk, RN => rst_BAR,
                           Q => n23744, QN => n_1386);
   clk_r_REG14101_S4 : DFFS_X1 port map( D => n12526, CK => clk, SN => rst_BAR,
                           Q => n23743, QN => n_1387);
   clk_r_REG14100_S4 : DFFR_X1 port map( D => n12526, CK => clk, RN => rst_BAR,
                           Q => n23742, QN => n_1388);
   clk_r_REG14286_S4 : DFFR_X1 port map( D => n1839, CK => clk, RN => rst_BAR, 
                           Q => n27694, QN => n23741);
   clk_r_REG14284_S3 : DFFS_X1 port map( D => n1835, CK => clk, SN => rst_BAR, 
                           Q => n27698, QN => n23740);
   clk_r_REG14239_S3 : DFFS_X1 port map( D => n19005, CK => clk, SN => rst_BAR,
                           Q => n23739, QN => n_1389);
   clk_r_REG14113_S4 : DFFR_X1 port map( D => n19004, CK => clk, RN => rst_BAR,
                           Q => n23738, QN => n_1390);
   clk_r_REG14244_S3 : DFFR_X1 port map( D => n19003, CK => clk, RN => rst_BAR,
                           Q => n23737, QN => n_1391);
   clk_r_REG14283_S3 : DFFS_X1 port map( D => n13963, CK => clk, SN => rst_BAR,
                           Q => n23736, QN => n_1392);
   clk_r_REG14108_S4 : DFFR_X1 port map( D => n19001, CK => clk, RN => rst_BAR,
                           Q => n23735, QN => n_1393);
   clk_r_REG14107_S4 : DFFR_X1 port map( D => n19000, CK => clk, RN => rst_BAR,
                           Q => n23734, QN => n_1394);
   clk_r_REG14106_S4 : DFFR_X1 port map( D => n18999, CK => clk, RN => rst_BAR,
                           Q => n23733, QN => n_1395);
   clk_r_REG14282_S4 : DFFR_X1 port map( D => n14004, CK => clk, RN => rst_BAR,
                           Q => n23732, QN => n_1396);
   clk_r_REG14238_S3 : DFFS_X1 port map( D => n18993, CK => clk, SN => rst_BAR,
                           Q => n23731, QN => n_1397);
   clk_r_REG14280_S3 : DFFS_X1 port map( D => n18992, CK => clk, SN => n25890, 
                           Q => n23730, QN => n_1398);
   clk_r_REG14261_S4 : DFFR_X1 port map( D => n1845, CK => clk, RN => rst_BAR, 
                           Q => n_1399, QN => n23729);
   clk_r_REG14248_S3 : DFFS_X1 port map( D => n18989, CK => clk, SN => rst_BAR,
                           Q => n23728, QN => n_1400);
   clk_r_REG14237_S3 : DFFS_X1 port map( D => n18988, CK => clk, SN => rst_BAR,
                           Q => n23727, QN => n_1401);
   clk_r_REG14007_S4 : DFFR_X1 port map( D => n1829, CK => clk, RN => rst_BAR, 
                           Q => n_1402, QN => n23726);
   clk_r_REG14247_S3 : DFFS_X1 port map( D => n18982, CK => clk, SN => rst_BAR,
                           Q => n23725, QN => n_1403);
   clk_r_REG14236_S3 : DFFS_X1 port map( D => n18981, CK => clk, SN => rst_BAR,
                           Q => n23724, QN => n_1404);
   clk_r_REG13847_S10 : DFFS_X1 port map( D => n19185, CK => clk, SN => n25890,
                           Q => n23723, QN => n_1405);
   clk_r_REG14240_S3 : DFFR_X1 port map( D => n21603, CK => clk, RN => rst_BAR,
                           Q => n23722, QN => n_1406);
   clk_r_REG14281_S3 : DFFR_X1 port map( D => n21604, CK => clk, RN => n25889, 
                           Q => n23721, QN => n_1407);
   clk_r_REG13834_S4 : DFFR_X1 port map( D => n21607, CK => clk, RN => rst_BAR,
                           Q => n23720, QN => n_1408);
   clk_r_REG14029_S10 : DFFS_X1 port map( D => n18980, CK => clk, SN => rst_BAR
                           , Q => n23719, QN => n_1409);
   clk_r_REG14049_S5 : DFFR_X1 port map( D => n21633, CK => clk, RN => rst_BAR,
                           Q => n23718, QN => n_1410);
   clk_r_REG14230_S3 : DFFS_X1 port map( D => n18977, CK => clk, SN => n25890, 
                           Q => n23717, QN => n_1411);
   clk_r_REG14153_S3 : DFFS_X1 port map( D => n18974, CK => clk, SN => rst_BAR,
                           Q => n23716, QN => n_1412);
   clk_r_REG14138_S10 : DFFS_X1 port map( D => n18973, CK => clk, SN => rst_BAR
                           , Q => n23715, QN => n_1413);
   clk_r_REG14152_S4 : DFFS_X1 port map( D => n18972, CK => clk, SN => rst_BAR,
                           Q => n23714, QN => n_1414);
   clk_r_REG14695_S4 : DFFS_X1 port map( D => n18969, CK => clk, SN => rst_BAR,
                           Q => n23713, QN => n_1415);
   clk_r_REG14157_S3 : DFFS_X1 port map( D => n18968, CK => clk, SN => rst_BAR,
                           Q => n23712, QN => n_1416);
   clk_r_REG14694_S4 : DFFR_X1 port map( D => n18967, CK => clk, RN => rst_BAR,
                           Q => n23711, QN => n_1417);
   clk_r_REG14115_S4 : DFFR_X1 port map( D => n1817, CK => clk, RN => rst_BAR, 
                           Q => n_1418, QN => n23710);
   clk_r_REG14311_S3 : DFFS_X1 port map( D => n18965, CK => clk, SN => rst_BAR,
                           Q => n23709, QN => n_1419);
   clk_r_REG14691_S3 : DFFS_X1 port map( D => n18964, CK => clk, SN => n25890, 
                           Q => n23708, QN => n_1420);
   clk_r_REG14279_S4 : DFFR_X1 port map( D => n21746, CK => clk, RN => rst_BAR,
                           Q => n23707, QN => n_1421);
   clk_r_REG14304_S3 : DFFR_X1 port map( D => n21745, CK => clk, RN => rst_BAR,
                           Q => n23706, QN => n_1422);
   clk_r_REG14260_S3 : DFFR_X1 port map( D => n11966, CK => clk, RN => rst_BAR,
                           Q => n23705, QN => n_1423);
   clk_r_REG14259_S3 : DFFR_X1 port map( D => n21841, CK => clk, RN => rst_BAR,
                           Q => n27685, QN => n25861);
   clk_r_REG14258_S3 : DFFS_X1 port map( D => n21841, CK => clk, SN => rst_BAR,
                           Q => n23703, QN => n_1424);
   clk_r_REG14277_S3 : DFFS_X1 port map( D => n21843, CK => clk, SN => rst_BAR,
                           Q => n23702, QN => n_1425);
   clk_r_REG14257_S3 : DFFS_X1 port map( D => n18954, CK => clk, SN => rst_BAR,
                           Q => n23701, QN => n_1426);
   clk_r_REG14112_S4 : DFFS_X1 port map( D => n18952, CK => clk, SN => rst_BAR,
                           Q => n23700, QN => n_1427);
   clk_r_REG14111_S4 : DFFR_X1 port map( D => n18950, CK => clk, RN => rst_BAR,
                           Q => n23699, QN => n_1428);
   clk_r_REG14096_S4 : DFFR_X1 port map( D => n1822, CK => clk, RN => rst_BAR, 
                           Q => n_1429, QN => n23698);
   clk_r_REG14097_S4 : DFFR_X1 port map( D => n18949, CK => clk, RN => n25889, 
                           Q => n23697, QN => n_1430);
   clk_r_REG14105_S4 : DFFR_X1 port map( D => n18948, CK => clk, RN => rst_BAR,
                           Q => n23696, QN => n_1431);
   clk_r_REG14255_S3 : DFFR_X1 port map( D => n21842, CK => clk, RN => rst_BAR,
                           Q => n23695, QN => n_1432);
   clk_r_REG14235_S3 : DFFS_X1 port map( D => n18946, CK => clk, SN => rst_BAR,
                           Q => n23694, QN => n_1433);
   clk_r_REG13706_S5 : DFFS_X1 port map( D => n18945, CK => clk, SN => rst_BAR,
                           Q => n23693, QN => n_1434);
   clk_r_REG14234_S3 : DFFS_X1 port map( D => n21845, CK => clk, SN => rst_BAR,
                           Q => n23692, QN => n_1435);
   clk_r_REG13699_S7 : DFFR_X1 port map( D => n18935, CK => clk, RN => rst_BAR,
                           Q => n23691, QN => n_1436);
   clk_r_REG14310_S3 : DFFS_X1 port map( D => n18934, CK => clk, SN => rst_BAR,
                           Q => n23690, QN => n_1437);
   clk_r_REG14835_S10 : DFFS_X1 port map( D => n18933, CK => clk, SN => rst_BAR
                           , Q => n23689, QN => n_1438);
   clk_r_REG14063_S4 : DFFR_X1 port map( D => n1806, CK => clk, RN => rst_BAR, 
                           Q => n_1439, QN => n25864);
   clk_r_REG14062_S4 : DFFS_X1 port map( D => n1806, CK => clk, SN => rst_BAR, 
                           Q => n23687, QN => n_1440);
   clk_r_REG13788_S4 : DFFS_X1 port map( D => n18930, CK => clk, SN => rst_BAR,
                           Q => n23686, QN => n_1441);
   clk_r_REG13787_S4 : DFFS_X1 port map( D => n18929, CK => clk, SN => rst_BAR,
                           Q => n23685, QN => n_1442);
   clk_r_REG13889_S11 : DFFS_X1 port map( D => n18927, CK => clk, SN => rst_BAR
                           , Q => n23684, QN => n_1443);
   clk_r_REG13762_S4 : DFFS_X1 port map( D => n18926, CK => clk, SN => rst_BAR,
                           Q => n23683, QN => n_1444);
   clk_r_REG13755_S7 : DFFS_X1 port map( D => n18925, CK => clk, SN => rst_BAR,
                           Q => n23682, QN => n_1445);
   clk_r_REG13748_S4 : DFFS_X1 port map( D => n19179, CK => clk, SN => rst_BAR,
                           Q => n23681, QN => n_1446);
   clk_r_REG13739_S4 : DFFS_X1 port map( D => n22091, CK => clk, SN => rst_BAR,
                           Q => n23680, QN => n_1447);
   clk_r_REG13732_S4 : DFFR_X1 port map( D => n18923, CK => clk, RN => rst_BAR,
                           Q => n23679, QN => n_1448);
   clk_r_REG13949_S10 : DFFS_X1 port map( D => n18922, CK => clk, SN => rst_BAR
                           , Q => n23678, QN => n_1449);
   clk_r_REG13717_S4 : DFFS_X1 port map( D => n18921, CK => clk, SN => rst_BAR,
                           Q => n23677, QN => n_1450);
   clk_r_REG13822_S4 : DFFS_X1 port map( D => n19172, CK => clk, SN => rst_BAR,
                           Q => n23676, QN => n_1451);
   clk_r_REG14975_S10 : DFFS_X1 port map( D => n18920, CK => clk, SN => n25890,
                           Q => n23675, QN => n_1452);
   clk_r_REG14061_S4 : DFFS_X1 port map( D => n22532, CK => clk, SN => n25890, 
                           Q => n23674, QN => n_1453);
   clk_r_REG14117_S4 : DFFR_X1 port map( D => n18918, CK => clk, RN => rst_BAR,
                           Q => n23673, QN => n_1454);
   clk_r_REG13808_S4 : DFFS_X1 port map( D => n18916, CK => clk, SN => rst_BAR,
                           Q => n23672, QN => n_1455);
   clk_r_REG13977_S10 : DFFS_X1 port map( D => n18915, CK => clk, SN => rst_BAR
                           , Q => n23671, QN => n_1456);
   clk_r_REG13801_S4 : DFFR_X1 port map( D => n18914, CK => clk, RN => rst_BAR,
                           Q => n23670, QN => n_1457);
   clk_r_REG13985_S4 : DFFR_X1 port map( D => n18913, CK => clk, RN => rst_BAR,
                           Q => n23669, QN => n_1458);
   clk_r_REG13983_S10 : DFFS_X1 port map( D => n18912, CK => clk, SN => rst_BAR
                           , Q => n23668, QN => n_1459);
   clk_r_REG13799_S4 : DFFS_X1 port map( D => n18911, CK => clk, SN => rst_BAR,
                           Q => n23667, QN => n_1460);
   clk_r_REG13915_S10 : DFFS_X1 port map( D => n18910, CK => clk, SN => rst_BAR
                           , Q => n23666, QN => n_1461);
   clk_r_REG13685_S7 : DFFR_X1 port map( D => n18909, CK => clk, RN => rst_BAR,
                           Q => n23665, QN => n_1462);
   clk_r_REG14104_S4 : DFFR_X1 port map( D => n22276, CK => clk, RN => rst_BAR,
                           Q => n23664, QN => n_1463);
   clk_r_REG13657_S7 : DFFS_X1 port map( D => n19164, CK => clk, SN => rst_BAR,
                           Q => n23663, QN => n_1464);
   clk_r_REG13646_S10 : DFFS_X1 port map( D => n18904, CK => clk, SN => rst_BAR
                           , Q => n23662, QN => n_1465);
   clk_r_REG13714_S4 : DFFR_X1 port map( D => n18903, CK => clk, RN => rst_BAR,
                           Q => n23661, QN => n_1466);
   clk_r_REG14060_S4 : DFFS_X1 port map( D => n18902, CK => clk, SN => rst_BAR,
                           Q => n23660, QN => n_1467);
   clk_r_REG14038_S6 : DFFR_X1 port map( D => n18899, CK => clk, RN => rst_BAR,
                           Q => n23659, QN => n_1468);
   clk_r_REG14039_S6 : DFFR_X1 port map( D => n18898, CK => clk, RN => rst_BAR,
                           Q => n23658, QN => n_1469);
   clk_r_REG14040_S6 : DFFR_X1 port map( D => n18897, CK => clk, RN => rst_BAR,
                           Q => n23657, QN => n_1470);
   clk_r_REG14041_S6 : DFFR_X1 port map( D => n18896, CK => clk, RN => rst_BAR,
                           Q => n23656, QN => n_1471);
   clk_r_REG14042_S6 : DFFR_X1 port map( D => n18895, CK => clk, RN => rst_BAR,
                           Q => n23655, QN => n_1472);
   clk_r_REG14043_S6 : DFFR_X1 port map( D => n18894, CK => clk, RN => rst_BAR,
                           Q => n23654, QN => n_1473);
   clk_r_REG13990_S6 : DFFR_X1 port map( D => n18893, CK => clk, RN => rst_BAR,
                           Q => n23653, QN => n_1474);
   clk_r_REG13680_S5 : DFFR_X1 port map( D => n19247, CK => clk, RN => rst_BAR,
                           Q => n23652, QN => n_1475);
   clk_r_REG13910_S5 : DFFR_X1 port map( D => n19246, CK => clk, RN => n25889, 
                           Q => n23651, QN => n_1476);
   clk_r_REG14340_S5 : DFFR_X1 port map( D => n19245, CK => clk, RN => rst_BAR,
                           Q => n23650, QN => n_1477);
   clk_r_REG14342_S5 : DFFR_X1 port map( D => n19244, CK => clk, RN => rst_BAR,
                           Q => n23649, QN => n_1478);
   clk_r_REG14351_S5 : DFFR_X1 port map( D => n19243, CK => clk, RN => rst_BAR,
                           Q => n23648, QN => n_1479);
   clk_r_REG14353_S5 : DFFR_X1 port map( D => n19242, CK => clk, RN => rst_BAR,
                           Q => n23647, QN => n_1480);
   clk_r_REG14355_S5 : DFFR_X1 port map( D => n19241, CK => clk, RN => rst_BAR,
                           Q => n23646, QN => n_1481);
   clk_r_REG14357_S5 : DFFR_X1 port map( D => n19240, CK => clk, RN => n25889, 
                           Q => n23645, QN => n_1482);
   clk_r_REG14359_S5 : DFFR_X1 port map( D => n19239, CK => clk, RN => rst_BAR,
                           Q => n23644, QN => n_1483);
   clk_r_REG14361_S5 : DFFR_X1 port map( D => n19238, CK => clk, RN => rst_BAR,
                           Q => n23643, QN => n_1484);
   clk_r_REG14363_S5 : DFFR_X1 port map( D => n19237, CK => clk, RN => rst_BAR,
                           Q => n23642, QN => n_1485);
   clk_r_REG14365_S5 : DFFR_X1 port map( D => n19236, CK => clk, RN => rst_BAR,
                           Q => n23641, QN => n_1486);
   clk_r_REG14367_S5 : DFFR_X1 port map( D => n19235, CK => clk, RN => rst_BAR,
                           Q => n23640, QN => n_1487);
   clk_r_REG13988_S5 : DFFR_X1 port map( D => n18892, CK => clk, RN => rst_BAR,
                           Q => n23639, QN => n_1488);
   clk_r_REG13791_S4 : DFFR_X1 port map( D => n1833, CK => clk, RN => rst_BAR, 
                           Q => n_1489, QN => n23638);
   clk_r_REG14052_S5 : DFFS_X1 port map( D => n18878, CK => clk, SN => n25890, 
                           Q => n23637, QN => n_1490);
   clk_r_REG13829_S4 : DFFS_X1 port map( D => n18877, CK => clk, SN => rst_BAR,
                           Q => n23636, QN => n_1491);
   clk_r_REG14170_S3 : DFFR_X1 port map( D => n25867, CK => clk, RN => rst_BAR,
                           Q => n_1492, QN => n23635);
   clk_r_REG14169_S3 : DFFS_X1 port map( D => n25867, CK => clk, SN => rst_BAR,
                           Q => n_1493, QN => n23634);
   clk_r_REG14165_S3 : DFFR_X1 port map( D => n25865, CK => clk, RN => rst_BAR,
                           Q => n_1494, QN => n23632);
   clk_r_REG14164_S3 : DFFS_X1 port map( D => n25865, CK => clk, SN => rst_BAR,
                           Q => n_1495, QN => n23631);
   clk_r_REG14178_S3 : DFFS_X1 port map( D => n25859, CK => clk, SN => n25890, 
                           Q => n27672, QN => n23630);
   clk_r_REG13833_S4 : DFFS_X1 port map( D => n1837, CK => clk, SN => rst_BAR, 
                           Q => n_1496, QN => n23629);
   clk_r_REG14229_S3 : DFFS_X1 port map( D => n19419, CK => clk, SN => rst_BAR,
                           Q => n23628, QN => n_1497);
   clk_r_REG14345_S6 : DFFR_X1 port map( D => n18872, CK => clk, RN => rst_BAR,
                           Q => n23627, QN => n_1498);
   clk_r_REG14346_S7 : DFFR_X1 port map( D => n23627, CK => clk, RN => rst_BAR,
                           Q => n23626, QN => n_1499);
   clk_r_REG14347_S8 : DFFR_X1 port map( D => n23626, CK => clk, RN => n25889, 
                           Q => n23625, QN => n_1500);
   clk_r_REG14348_S9 : DFFR_X1 port map( D => n23625, CK => clk, RN => rst_BAR,
                           Q => n23624, QN => n_1501);
   clk_r_REG14349_S10 : DFFR_X1 port map( D => n23624, CK => clk, RN => rst_BAR
                           , Q => n23623, QN => n_1502);
   clk_r_REG14127_S5 : DFFR_X1 port map( D => n18867, CK => clk, RN => rst_BAR,
                           Q => n23622, QN => n_1503);
   clk_r_REG14128_S6 : DFFR_X1 port map( D => n23622, CK => clk, RN => rst_BAR,
                           Q => n23621, QN => n_1504);
   clk_r_REG14129_S7 : DFFR_X1 port map( D => n23621, CK => clk, RN => rst_BAR,
                           Q => n23620, QN => n_1505);
   clk_r_REG14130_S8 : DFFR_X1 port map( D => n23620, CK => clk, RN => rst_BAR,
                           Q => n23619, QN => n_1506);
   clk_r_REG14131_S9 : DFFR_X1 port map( D => n23619, CK => clk, RN => rst_BAR,
                           Q => n23618, QN => n_1507);
   clk_r_REG13856_S5 : DFFR_X1 port map( D => n19194, CK => clk, RN => rst_BAR,
                           Q => n23617, QN => n_1508);
   clk_r_REG13857_S6 : DFFR_X1 port map( D => n23617, CK => clk, RN => rst_BAR,
                           Q => n23616, QN => n_1509);
   clk_r_REG13858_S7 : DFFR_X1 port map( D => n23616, CK => clk, RN => rst_BAR,
                           Q => n23615, QN => n_1510);
   clk_r_REG13859_S8 : DFFR_X1 port map( D => n23615, CK => clk, RN => rst_BAR,
                           Q => n23614, QN => n_1511);
   clk_r_REG13860_S9 : DFFR_X1 port map( D => n23614, CK => clk, RN => rst_BAR,
                           Q => n23613, QN => n_1512);
   clk_r_REG14976_S4 : DFFS_X1 port map( D => n18860, CK => clk, SN => rst_BAR,
                           Q => n23612, QN => n_1513);
   clk_r_REG13681_S6 : DFFR_X1 port map( D => n18856, CK => clk, RN => rst_BAR,
                           Q => n23611, QN => n_1514);
   clk_r_REG13682_S7 : DFFR_X1 port map( D => n23611, CK => clk, RN => rst_BAR,
                           Q => n23610, QN => n_1515);
   clk_r_REG13683_S8 : DFFR_X1 port map( D => n23610, CK => clk, RN => rst_BAR,
                           Q => n23609, QN => n_1516);
   clk_r_REG13684_S9 : DFFR_X1 port map( D => n23609, CK => clk, RN => rst_BAR,
                           Q => n23608, QN => n_1517);
   clk_r_REG14055_S5 : DFFS_X1 port map( D => n18855, CK => clk, SN => rst_BAR,
                           Q => n23607, QN => n_1518);
   clk_r_REG14054_S5 : DFFR_X1 port map( D => n18854, CK => clk, RN => rst_BAR,
                           Q => n23606, QN => n_1519);
   clk_r_REG13713_S4 : DFFS_X1 port map( D => n18853, CK => clk, SN => rst_BAR,
                           Q => n23605, QN => n_1520);
   clk_r_REG14003_S5 : DFFR_X1 port map( D => n18852, CK => clk, RN => rst_BAR,
                           Q => n23604, QN => n_1521);
   clk_r_REG14002_S5 : DFFR_X1 port map( D => n18850, CK => clk, RN => n25889, 
                           Q => n23603, QN => n_1522);
   clk_r_REG13984_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_15_port, CK => clk, 
                           RN => rst_BAR, Q => n23602, QN => n_1523);
   clk_r_REG14306_S3 : DFFS_X1 port map( D => n1846, CK => clk, SN => rst_BAR, 
                           Q => n_1524, QN => n23601);
   clk_r_REG14305_S3 : DFFS_X1 port map( D => n1848, CK => clk, SN => rst_BAR, 
                           Q => n_1525, QN => n23600);
   clk_r_REG14313_S3 : DFFS_X1 port map( D => n18848, CK => clk, SN => rst_BAR,
                           Q => n23599, QN => n_1526);
   clk_r_REG13998_S5 : DFFR_X1 port map( D => n18846, CK => clk, RN => rst_BAR,
                           Q => n23598, QN => n_1527);
   clk_r_REG13875_S6 : DFFR_X1 port map( D => n18845, CK => clk, RN => rst_BAR,
                           Q => n23597, QN => n_1528);
   clk_r_REG14969_S4 : DFFR_X1 port map( D => n18839, CK => clk, RN => rst_BAR,
                           Q => n23596, QN => n_1529);
   clk_r_REG14970_S5 : DFFR_X1 port map( D => n23596, CK => clk, RN => rst_BAR,
                           Q => n23595, QN => n_1530);
   clk_r_REG14971_S6 : DFFR_X1 port map( D => n23595, CK => clk, RN => rst_BAR,
                           Q => n23594, QN => n_1531);
   clk_r_REG14972_S7 : DFFR_X1 port map( D => n23594, CK => clk, RN => rst_BAR,
                           Q => n23593, QN => n_1532);
   clk_r_REG14973_S8 : DFFR_X1 port map( D => n23593, CK => clk, RN => rst_BAR,
                           Q => n23592, QN => n_1533);
   clk_r_REG14974_S9 : DFFR_X1 port map( D => n23592, CK => clk, RN => rst_BAR,
                           Q => n23591, QN => n_1534);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n554, Q => 
                           DATA2_I_26_port);
   clk_r_REG14333_S3 : DFFR_X1 port map( D => n1858, CK => clk, RN => rst_BAR, 
                           Q => n27669, QN => n24156);
   clk_r_REG14330_S3 : DFFR_X1 port map( D => n1843, CK => clk, RN => rst_BAR, 
                           Q => n27667, QN => n24158);
   clk_r_REG14224_S3 : DFFR_X1 port map( D => n25870, CK => clk, RN => rst_BAR,
                           Q => n27666, QN => n23633);
   clk_r_REG14321_S3 : DFFR_X1 port map( D => n25879, CK => clk, RN => rst_BAR,
                           Q => n27662, QN => n23979);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n7822, Q => 
                           data1_mul_15_port);
   clk_r_REG15178_S5 : DFFS_X1 port map( D => n1810, CK => clk, SN => rst_BAR, 
                           Q => n24127, QN => n_1535);
   clk_r_REG13679_S4 : DFFR_X1 port map( D => n25883, CK => clk, RN => n25889, 
                           Q => n24133, QN => n_1536);
   clk_r_REG13873_S5 : DFFR_X1 port map( D => n19291, CK => clk, RN => n25889, 
                           Q => n24000, QN => n_1537);
   clk_r_REG13909_S4 : DFFS_X1 port map( D => n22800, CK => clk, SN => rst_BAR,
                           Q => n23897, QN => n_1538);
   clk_r_REG13664_S5 : DFFS_X1 port map( D => n19250, CK => clk, SN => rst_BAR,
                           Q => n24001, QN => n_1539);
   clk_r_REG15179_S5 : DFFR_X1 port map( D => n25888, CK => clk, RN => rst_BAR,
                           Q => n_1540, QN => n24037);
   clk_r_REG15113_S4 : DFFR_X1 port map( D => n22797, CK => clk, RN => rst_BAR,
                           Q => n24043, QN => n_1541);
   clk_r_REG15111_S4 : DFFS_X1 port map( D => n25882, CK => clk, SN => rst_BAR,
                           Q => n_1542, QN => n24042);
   clk_r_REG14232_S3 : DFFR_X1 port map( D => n1861, CK => clk, RN => rst_BAR, 
                           Q => n_1543, QN => n23954);
   clk_r_REG14088_S4 : DFFS_X1 port map( D => n1812, CK => clk, SN => rst_BAR, 
                           Q => n24129, QN => n_1544);
   clk_r_REG14089_S4 : DFFR_X1 port map( D => n21556, CK => clk, RN => rst_BAR,
                           Q => n_1545, QN => n24169);
   clk_r_REG14084_S4 : DFFR_X1 port map( D => n25885, CK => clk, RN => rst_BAR,
                           Q => n24130, QN => n_1546);
   clk_r_REG13855_S5 : DFFR_X1 port map( D => n25887, CK => clk, RN => rst_BAR,
                           Q => n24128, QN => n_1547);
   clk_r_REG14149_S4 : DFFR_X1 port map( D => n19200, CK => clk, RN => rst_BAR,
                           Q => n23949, QN => n_1548);
   clk_r_REG14047_S5 : DFFS_X1 port map( D => n19160, CK => clk, SN => rst_BAR,
                           Q => n24002, QN => n_1549);
   clk_r_REG14125_S4 : DFFS_X1 port map( D => n25884, CK => clk, SN => rst_BAR,
                           Q => n_1550, QN => n23972);
   clk_r_REG14036_S5 : DFFS_X1 port map( D => n25881, CK => clk, SN => rst_BAR,
                           Q => n_1551, QN => n23890);
   clk_r_REG14045_S5 : DFFR_X1 port map( D => n19280, CK => clk, RN => rst_BAR,
                           Q => n24027, QN => n_1552);
   clk_r_REG13841_S4 : DFFS_X1 port map( D => n19251, CK => clk, SN => rst_BAR,
                           Q => n24003, QN => n_1553);
   U3 : CLKBUF_X1 port map( A => rst_BAR, Z => n25889);
   U4 : CLKBUF_X1 port map( A => n25889, Z => n25890);
   U5 : OR2_X1 port map( A1 => n25968, A2 => n27624, ZN => n25891);
   U6 : INV_X1 port map( A => n25891, ZN => n25892);
   U7 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n25893);
   U8 : INV_X1 port map( A => n25893, ZN => n25894);
   U9 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n25895);
   U10 : INV_X1 port map( A => n25895, ZN => n25896);
   U11 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN => 
                           n25897);
   U12 : INV_X1 port map( A => n25897, ZN => n25898);
   U13 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n25899);
   U14 : INV_X1 port map( A => n25899, ZN => n25900);
   U15 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , A2 => n27281, ZN => n27310);
   U16 : NOR2_X2 port map( A1 => n25858, A2 => n22802, ZN => n27506);
   U17 : NOR2_X2 port map( A1 => n22802, A2 => n27700, ZN => n27505);
   U18 : OAI21_X2 port map( B1 => DATA2(1), B2 => n27583, A => n26013, ZN => 
                           n1836);
   U19 : NOR2_X2 port map( A1 => n26478, A2 => n27591, ZN => n26753);
   U20 : NOR2_X2 port map( A1 => n27281, A2 => n27314, ZN => n27316);
   U21 : INV_X2 port map( A => n26795, ZN => n27641);
   U22 : NOR3_X4 port map( A1 => n24044, A2 => n25872, A3 => n25858, ZN => 
                           n27507);
   U23 : INV_X1 port map( A => n26209, ZN => n26446);
   U24 : INV_X1 port map( A => n27570, ZN => n27557);
   U25 : INV_X1 port map( A => data1_mul_15_port, ZN => n1790);
   U26 : INV_X1 port map( A => n9045, ZN => n1791);
   U27 : INV_X1 port map( A => n9060, ZN => n1796);
   U28 : INV_X1 port map( A => n9075, ZN => n1802);
   U29 : INV_X1 port map( A => n554, ZN => n27249);
   U30 : OR3_X1 port map( A1 => n26166, A2 => n25977, A3 => n27645, ZN => 
                           n27638);
   U31 : NOR2_X1 port map( A1 => n27571, A2 => n27573, ZN => n27575);
   U32 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_2_4_port, ZN => 
                           n1801);
   U33 : INV_X1 port map( A => n7769, ZN => n27586);
   U34 : NAND3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4295, A3 => n27586, ZN => n1812);
   U35 : NOR2_X1 port map( A1 => n7769, A2 => n8978, ZN => n27584);
   U36 : AOI21_X1 port map( B1 => n8978, B2 => n7769, A => n27584, ZN => n1811)
                           ;
   U37 : INV_X1 port map( A => n14287, ZN => n27589);
   U38 : NAND3_X1 port map( A1 => n14286, A2 => n4302, A3 => n27589, ZN => 
                           n1810);
   U39 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n27320);
   U40 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n27320, ZN => n19213);
   U41 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_5_port, 
                           ZN => n27587);
   U42 : OR2_X1 port map( A1 => n27587, A2 => n19213, ZN => n25884);
   U43 : NOR2_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_2_5_port
                           , A2 => n4295, ZN => n27350);
   U44 : AOI21_X1 port map( B1 => n4295, B2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A =>
                           n27350, ZN => n1813);
   U45 : INV_X1 port map( A => cin, ZN => n1871);
   U46 : NOR2_X1 port map( A1 => DATA2(4), A2 => DATA2(5), ZN => n1863);
   U47 : INV_X1 port map( A => DATA2(1), ZN => n27571);
   U48 : INV_X1 port map( A => DATA2(0), ZN => n27573);
   U49 : INV_X1 port map( A => n1863, ZN => n27583);
   U50 : AOI21_X1 port map( B1 => DATA2(2), B2 => DATA2(3), A => n27583, ZN => 
                           n26014);
   U51 : INV_X1 port map( A => n26014, ZN => n26013);
   U52 : OAI21_X1 port map( B1 => n27575, B2 => n27583, A => n26013, ZN => 
                           n1841);
   U53 : INV_X1 port map( A => n1841, ZN => n1862);
   U54 : INV_X1 port map( A => DATA2(3), ZN => n27594);
   U55 : NOR2_X1 port map( A1 => n1863, A2 => n27594, ZN => n1865);
   U56 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n25942);
   U57 : INV_X1 port map( A => FUNC(2), ZN => n25941);
   U58 : NAND2_X1 port map( A1 => n25942, A2 => n25941, ZN => n554);
   U59 : INV_X1 port map( A => n27249, ZN => n27710);
   U60 : NAND2_X1 port map( A1 => n24176, A2 => DATA2_I_4_port, ZN => n25904);
   U61 : OAI21_X1 port map( B1 => n24176, B2 => DATA2_I_4_port, A => n25904, ZN
                           => n1429);
   U62 : NOR2_X1 port map( A1 => n24172, A2 => n27710, ZN => n27040);
   U63 : XNOR2_X1 port map( A => n24056, B => DATA2_I_5_port, ZN => n26360);
   U64 : INV_X1 port map( A => n26360, ZN => n26363);
   U65 : NAND2_X1 port map( A1 => n24048, A2 => DATA2_I_3_port, ZN => n25909);
   U66 : OAI21_X1 port map( B1 => n24048, B2 => DATA2_I_3_port, A => n25909, ZN
                           => n27532);
   U67 : INV_X1 port map( A => n27532, ZN => n25902);
   U68 : NAND2_X1 port map( A1 => n24049, A2 => DATA2_I_2_port, ZN => n25908);
   U69 : OAI21_X1 port map( B1 => n24049, B2 => DATA2_I_2_port, A => n25908, ZN
                           => n26670);
   U70 : INV_X1 port map( A => n26670, ZN => n26674);
   U71 : NAND2_X1 port map( A1 => n24173, A2 => DATA2_I_0_port, ZN => n26850);
   U72 : INV_X1 port map( A => n26850, ZN => n27035);
   U73 : AOI21_X1 port map( B1 => DATA2_I_1_port, B2 => n24175, A => n27035, ZN
                           => n25910);
   U74 : NOR2_X1 port map( A1 => n24175, A2 => DATA2_I_1_port, ZN => n25901);
   U75 : NOR2_X1 port map( A1 => n25910, A2 => n25901, ZN => n26673);
   U76 : NAND2_X1 port map( A1 => n26674, A2 => n26673, ZN => n26672);
   U77 : NAND2_X1 port map( A1 => n25908, A2 => n26672, ZN => n27531);
   U78 : NAND2_X1 port map( A1 => n25902, A2 => n27531, ZN => n25903);
   U79 : AND2_X1 port map( A1 => n25909, A2 => n25903, ZN => n26396);
   U80 : OAI21_X1 port map( B1 => n1429, B2 => n26396, A => n25904, ZN => 
                           n26358);
   U81 : INV_X1 port map( A => n26358, ZN => n26356);
   U82 : NAND2_X1 port map( A1 => n24177, A2 => DATA2_I_5_port, ZN => n25914);
   U83 : OAI21_X1 port map( B1 => n26363, B2 => n26356, A => n25914, ZN => 
                           n26325);
   U84 : NOR2_X1 port map( A1 => n24050, A2 => n27710, ZN => n26424);
   U85 : INV_X1 port map( A => n25904, ZN => n25913);
   U86 : INV_X1 port map( A => n25909, ZN => n25907);
   U87 : INV_X1 port map( A => n25908, ZN => n25906);
   U88 : NOR2_X1 port map( A1 => n24173, A2 => DATA2_I_0_port, ZN => n27034);
   U89 : NAND2_X1 port map( A1 => n24175, A2 => DATA2_I_1_port, ZN => n25905);
   U90 : OAI21_X1 port map( B1 => n24175, B2 => DATA2_I_1_port, A => n25905, ZN
                           => n26849);
   U91 : NOR2_X1 port map( A1 => n27034, A2 => n26849, ZN => n26844);
   U92 : AOI21_X1 port map( B1 => DATA2_I_1_port, B2 => n24175, A => n26844, ZN
                           => n26671);
   U93 : NOR2_X1 port map( A1 => n26671, A2 => n26670, ZN => n26669);
   U94 : NOR2_X1 port map( A1 => n25906, A2 => n26669, ZN => n26422);
   U95 : NOR2_X1 port map( A1 => n26422, A2 => n27532, ZN => n26421);
   U96 : NOR2_X1 port map( A1 => n25907, A2 => n26421, ZN => n26397);
   U97 : NOR2_X1 port map( A1 => n26397, A2 => n1429, ZN => n25912);
   U98 : NOR2_X1 port map( A1 => n25913, A2 => n25912, ZN => n26357);
   U99 : OAI21_X1 port map( B1 => n26363, B2 => n26357, A => n25914, ZN => 
                           n26326);
   U100 : AOI22_X1 port map( A1 => n27040, A2 => n26325, B1 => n26424, B2 => 
                           n26326, ZN => n26335);
   U101 : XNOR2_X1 port map( A => DATA2_I_6_port, B => n24077, ZN => n26329);
   U102 : OR2_X1 port map( A1 => n26335, A2 => n26329, ZN => n19270);
   U103 : XOR2_X1 port map( A => DATA1(21), B => DATA2_I_21_port, Z => n1809);
   U104 : XOR2_X1 port map( A => n24179, B => DATA2_I_7_port, Z => n26328);
   U105 : INV_X1 port map( A => n26329, ZN => n27539);
   U106 : NAND4_X1 port map( A1 => n25910, A2 => n24050, A3 => n25909, A4 => 
                           n25908, ZN => n25911);
   U107 : OAI221_X1 port map( B1 => n25913, B2 => n25912, C1 => n25913, C2 => 
                           n25911, A => n26360, ZN => n25915);
   U108 : NAND2_X1 port map( A1 => n24178, A2 => DATA2_I_6_port, ZN => n26333);
   U109 : OAI221_X1 port map( B1 => n27539, B2 => n25915, C1 => n27539, C2 => 
                           n25914, A => n26333, ZN => n25916);
   U110 : AOI22_X1 port map( A1 => n24179, A2 => DATA2_I_7_port, B1 => n26328, 
                           B2 => n25916, ZN => n26979);
   U111 : NAND2_X1 port map( A1 => n27249, A2 => n26979, ZN => n1789);
   U112 : NOR2_X1 port map( A1 => n24181, A2 => DATA2_I_8_port, ZN => n26266);
   U113 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => n24181, A => n26266, 
                           ZN => n21635);
   U114 : INV_X1 port map( A => DATA1(22), ZN => n27177);
   U115 : XNOR2_X1 port map( A => DATA2_I_22_port, B => n27177, ZN => n26808);
   U116 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n25950);
   U117 : INV_X1 port map( A => n25950, ZN => n25917);
   U118 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n25926);
   U119 : AND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n26899);
   U120 : INV_X1 port map( A => DATA1(17), ZN => n26915);
   U121 : XOR2_X1 port map( A => DATA2_I_17_port, B => n26915, Z => n26922);
   U122 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n26921);
   U123 : NOR2_X1 port map( A1 => n26922, A2 => n26921, ZN => n26920);
   U124 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => 
                           n25926, ZN => n25953);
   U125 : INV_X1 port map( A => n25953, ZN => n26900);
   U126 : OAI21_X1 port map( B1 => n26899, B2 => n26920, A => n26900, ZN => 
                           n26901);
   U127 : NAND2_X1 port map( A1 => n25926, A2 => n26901, ZN => n26884);
   U128 : AOI22_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, B1 => 
                           n25917, B2 => n26884, ZN => n26832);
   U129 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n25928);
   U130 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n25928, ZN => n26831);
   U131 : NOR2_X1 port map( A1 => n26832, A2 => n26831, ZN => n26830);
   U132 : AOI21_X1 port map( B1 => DATA2_I_20_port, B2 => DATA1(20), A => 
                           n26830, ZN => n27650);
   U133 : INV_X1 port map( A => n27650, ZN => n27558);
   U134 : AND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n25929);
   U135 : AOI21_X1 port map( B1 => n27558, B2 => n1809, A => n25929, ZN => 
                           n25930);
   U136 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n25948);
   U137 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n25948, ZN => n25922);
   U138 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n25947
                           );
   U139 : OAI21_X1 port map( B1 => DATA1(9), B2 => DATA2_I_9_port, A => n25947,
                           ZN => n26265);
   U140 : INV_X1 port map( A => DATA1(14), ZN => n26964);
   U141 : XOR2_X1 port map( A => DATA2_I_14_port, B => n26964, Z => n26968);
   U142 : INV_X1 port map( A => n21635, ZN => n25919);
   U143 : INV_X1 port map( A => DATA1(13), ZN => n26977);
   U144 : INV_X1 port map( A => DATA2_I_13_port, ZN => n25918);
   U145 : NOR2_X1 port map( A1 => n26977, A2 => n25918, ZN => n26962);
   U146 : AOI21_X1 port map( B1 => n26977, B2 => n25918, A => n26962, ZN => 
                           n26987);
   U147 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n26976);
   U148 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => 
                           n26976, ZN => n27552);
   U149 : INV_X1 port map( A => n27552, ZN => n26996);
   U150 : NAND2_X1 port map( A1 => n26987, A2 => n26996, ZN => n26946);
   U151 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n25921);
   U152 : AOI21_X1 port map( B1 => DATA2_I_11_port, B2 => DATA1(11), A => 
                           n25921, ZN => n27009);
   U153 : INV_X1 port map( A => n27009, ZN => n27011);
   U154 : OR4_X1 port map( A1 => n26968, A2 => n25919, A3 => n26946, A4 => 
                           n27011, ZN => n25920);
   U155 : NOR4_X1 port map( A1 => n26979, A2 => n25922, A3 => n26265, A4 => 
                           n25920, ZN => n25925);
   U156 : XOR2_X1 port map( A => DATA1(15), B => DATA2_I_15_port, Z => n26950);
   U157 : INV_X1 port map( A => n25921, ZN => n25923);
   U158 : INV_X1 port map( A => n25922, ZN => n27023);
   U159 : INV_X1 port map( A => n26265, ZN => n26269);
   U160 : NAND3_X1 port map( A1 => n24181, A2 => n26269, A3 => DATA2_I_8_port, 
                           ZN => n26267);
   U161 : NAND2_X1 port map( A1 => n25947, A2 => n26267, ZN => n27022);
   U162 : NAND2_X1 port map( A1 => n27023, A2 => n27022, ZN => n27020);
   U163 : NAND2_X1 port map( A1 => n25948, A2 => n27020, ZN => n27008);
   U164 : AOI22_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, B1 => 
                           n25923, B2 => n27008, ZN => n26994);
   U165 : NAND3_X1 port map( A1 => DATA1(12), A2 => n26987, A3 => 
                           DATA2_I_12_port, ZN => n26945);
   U166 : OAI21_X1 port map( B1 => n26994, B2 => n26946, A => n26945, ZN => 
                           n26960);
   U167 : NOR2_X1 port map( A1 => n26962, A2 => n26960, ZN => n26966);
   U168 : NAND2_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, ZN => 
                           n26947);
   U169 : OAI21_X1 port map( B1 => n26966, B2 => n26968, A => n26947, ZN => 
                           n26940);
   U170 : AND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n25924);
   U171 : AOI221_X1 port map( B1 => n25925, B2 => n26950, C1 => n26940, C2 => 
                           n26950, A => n25924, ZN => n25954);
   U172 : NAND2_X1 port map( A1 => n27249, A2 => n25954, ZN => n26919);
   U173 : INV_X1 port map( A => n26831, ZN => n26836);
   U174 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n26918);
   U175 : NOR2_X1 port map( A1 => n26918, A2 => n26922, ZN => n26917);
   U176 : OAI21_X1 port map( B1 => n26899, B2 => n26917, A => n26900, ZN => 
                           n26904);
   U177 : NAND2_X1 port map( A1 => n25926, A2 => n26904, ZN => n26885);
   U178 : INV_X1 port map( A => n26885, ZN => n26882);
   U179 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n25927);
   U180 : OAI21_X1 port map( B1 => n25950, B2 => n26882, A => n25927, ZN => 
                           n26835);
   U181 : NAND2_X1 port map( A1 => n26836, A2 => n26835, ZN => n26834);
   U182 : NAND2_X1 port map( A1 => n25928, A2 => n26834, ZN => n27646);
   U183 : AOI21_X1 port map( B1 => n1809, B2 => n27646, A => n25929, ZN => 
                           n25931);
   U184 : NOR2_X1 port map( A1 => n25954, A2 => n27710, ZN => n27648);
   U185 : INV_X1 port map( A => n27648, ZN => n26916);
   U186 : OAI22_X1 port map( A1 => n25930, A2 => n26919, B1 => n25931, B2 => 
                           n26916, ZN => n26806);
   U187 : INV_X1 port map( A => n25930, ZN => n25955);
   U188 : NAND2_X1 port map( A1 => n27648, A2 => n25931, ZN => n25932);
   U189 : OAI211_X1 port map( C1 => n25955, C2 => n26919, A => n26808, B => 
                           n25932, ZN => n26802);
   U190 : OAI21_X1 port map( B1 => n26808, B2 => n26806, A => n26802, ZN => 
                           n25933);
   U191 : INV_X1 port map( A => n25933, ZN => n19175);
   U192 : INV_X1 port map( A => FUNC(3), ZN => n1832);
   U193 : NAND3_X1 port map( A1 => FUNC(2), A2 => n25942, A3 => n1832, ZN => 
                           n7822);
   U194 : NOR4_X1 port map( A1 => DATA2(13), A2 => DATA2(12), A3 => DATA2(11), 
                           A4 => DATA2(6), ZN => n25940);
   U195 : NOR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n26166);
   U196 : NAND2_X1 port map( A1 => n1863, A2 => n27594, ZN => n25968);
   U197 : OR2_X1 port map( A1 => DATA2(2), A2 => n25968, ZN => n26478);
   U198 : INV_X1 port map( A => n26478, ZN => n26461);
   U199 : NAND2_X1 port map( A1 => n26166, A2 => n26461, ZN => n26666);
   U200 : INV_X1 port map( A => DATA2(15), ZN => n27266);
   U201 : INV_X1 port map( A => DATA2(14), ZN => n27267);
   U202 : INV_X1 port map( A => DATA2(10), ZN => n27270);
   U203 : INV_X1 port map( A => DATA2(8), ZN => n27272);
   U204 : NAND4_X1 port map( A1 => n27266, A2 => n27267, A3 => n27270, A4 => 
                           n27272, ZN => n25934);
   U205 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(7), A3 => n26666, A4 =>
                           n25934, ZN => n25939);
   U206 : INV_X1 port map( A => DATA1(12), ZN => n27547);
   U207 : INV_X1 port map( A => DATA1(9), ZN => n25975);
   U208 : NAND4_X1 port map( A1 => n26964, A2 => n26977, A3 => n27547, A4 => 
                           n25975, ZN => n25937);
   U209 : NOR4_X1 port map( A1 => DATA1(11), A2 => n24181, A3 => n24049, A4 => 
                           n24179, ZN => n25935);
   U210 : INV_X1 port map( A => DATA1(15), ZN => n26943);
   U211 : INV_X1 port map( A => DATA1(10), ZN => n27151);
   U212 : NAND4_X1 port map( A1 => n24052, A2 => n25935, A3 => n26943, A4 => 
                           n27151, ZN => n25936);
   U213 : NOR4_X1 port map( A1 => n24178, A2 => n23762, A3 => n25937, A4 => 
                           n25936, ZN => n25938);
   U214 : AOI211_X1 port map( C1 => n25940, C2 => n25939, A => n25938, B => 
                           n7822, ZN => n22313);
   U215 : INV_X1 port map( A => FUNC(0), ZN => n27077);
   U216 : NAND3_X1 port map( A1 => n25941, A2 => n27077, A3 => FUNC(1), ZN => 
                           n27570);
   U217 : INV_X1 port map( A => DATA2(11), ZN => n27269);
   U218 : NOR2_X1 port map( A1 => DATA1(11), A2 => n27269, ZN => n27150);
   U219 : INV_X1 port map( A => DATA1(11), ZN => n25995);
   U220 : NOR2_X1 port map( A1 => DATA2(11), A2 => n25995, ZN => n27096);
   U221 : CLKBUF_X1 port map( A => n22313, Z => n27542);
   U222 : NAND2_X1 port map( A1 => n27557, A2 => n1832, ZN => n27018);
   U223 : NAND3_X1 port map( A1 => FUNC(2), A2 => FUNC(3), A3 => n25942, ZN => 
                           n27033);
   U224 : NAND2_X1 port map( A1 => n27018, A2 => n27033, ZN => n26981);
   U225 : INV_X1 port map( A => n26981, ZN => n27549);
   U226 : NOR3_X1 port map( A1 => n27549, A2 => n27269, A3 => n25995, ZN => 
                           n25943);
   U227 : AOI21_X1 port map( B1 => n23838, B2 => n27542, A => n25943, ZN => 
                           n25944);
   U228 : INV_X1 port map( A => n25944, ZN => n25945);
   U229 : AOI221_X1 port map( B1 => n27557, B2 => n27150, C1 => n27557, C2 => 
                           n27096, A => n25945, ZN => n25946);
   U230 : INV_X1 port map( A => n25946, ZN => n1824);
   U231 : OAI21_X1 port map( B1 => n26266, B2 => n26265, A => n25947, ZN => 
                           n27017);
   U232 : NAND2_X1 port map( A1 => n27023, A2 => n27017, ZN => n27016);
   U233 : NAND2_X1 port map( A1 => n25948, A2 => n27016, ZN => n27010);
   U234 : NAND2_X1 port map( A1 => n27009, A2 => n27010, ZN => n17503);
   U235 : INV_X1 port map( A => DATA1(29), ZN => n26703);
   U236 : XOR2_X1 port map( A => n4395, B => n26703, Z => n26713);
   U237 : INV_X1 port map( A => n26713, ZN => n1815);
   U238 : INV_X1 port map( A => DATA1(28), ZN => n27198);
   U239 : XNOR2_X1 port map( A => DATA2_I_28_port, B => n27198, ZN => n25963);
   U240 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n26757);
   U241 : INV_X1 port map( A => DATA1(25), ZN => n26773);
   U242 : XNOR2_X1 port map( A => DATA2_I_25_port, B => n26773, ZN => n26776);
   U243 : NAND3_X1 port map( A1 => DATA1(24), A2 => n26776, A3 => 
                           DATA2_I_24_port, ZN => n26770);
   U244 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n25949);
   U245 : OAI21_X1 port map( B1 => DATA1(26), B2 => DATA2_I_26_port, A => 
                           n25949, ZN => n26756);
   U246 : AOI21_X1 port map( B1 => n26757, B2 => n26770, A => n26756, ZN => 
                           n26758);
   U247 : AOI21_X1 port map( B1 => DATA2_I_26_port, B2 => DATA1(26), A => 
                           n26758, ZN => n26736);
   U248 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n25960);
   U249 : OAI21_X1 port map( B1 => DATA1(27), B2 => DATA2_I_27_port, A => 
                           n25960, ZN => n26745);
   U250 : OAI21_X1 port map( B1 => n26736, B2 => n26745, A => n25960, ZN => 
                           n25959);
   U251 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n25957);
   U252 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => 
                           n25957, ZN => n26807);
   U253 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n26804);
   U254 : INV_X1 port map( A => n26922, ZN => n25951);
   U255 : AOI21_X1 port map( B1 => DATA2_I_19_port, B2 => DATA1(19), A => 
                           n25950, ZN => n26889);
   U256 : AOI21_X1 port map( B1 => DATA2_I_16_port, B2 => DATA1(16), A => 
                           n26918, ZN => n26932);
   U257 : NAND4_X1 port map( A1 => n25951, A2 => n1809, A3 => n26889, A4 => 
                           n26932, ZN => n25952);
   U258 : NOR4_X1 port map( A1 => n25954, A2 => n25953, A3 => n26831, A4 => 
                           n25952, ZN => n25956);
   U259 : OAI21_X1 port map( B1 => n25956, B2 => n25955, A => n26808, ZN => 
                           n25958);
   U260 : OAI221_X1 port map( B1 => n26807, B2 => n26804, C1 => n26807, C2 => 
                           n25958, A => n25957, ZN => n25961);
   U261 : NOR2_X1 port map( A1 => n27710, A2 => n25961, ZN => n26786);
   U262 : NAND2_X1 port map( A1 => n25963, A2 => n25959, ZN => n27659);
   U263 : OAI211_X1 port map( C1 => n25963, C2 => n25959, A => n26786, B => 
                           n27659, ZN => n25965);
   U264 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n26787);
   U265 : INV_X1 port map( A => n26787, ZN => n26784);
   U266 : NAND2_X1 port map( A1 => n26776, A2 => n26784, ZN => n26775);
   U267 : AOI21_X1 port map( B1 => n26757, B2 => n26775, A => n26756, ZN => 
                           n26759);
   U268 : AOI21_X1 port map( B1 => DATA2_I_26_port, B2 => DATA1(26), A => 
                           n26759, ZN => n26735);
   U269 : OAI21_X1 port map( B1 => n26735, B2 => n26745, A => n25960, ZN => 
                           n25962);
   U270 : NAND2_X1 port map( A1 => n25961, A2 => n27249, ZN => n27658);
   U271 : INV_X1 port map( A => n27658, ZN => n26788);
   U272 : NAND2_X1 port map( A1 => n25963, A2 => n25962, ZN => n27657);
   U273 : OAI211_X1 port map( C1 => n25963, C2 => n25962, A => n26788, B => 
                           n27657, ZN => n25964);
   U274 : AND2_X1 port map( A1 => n25965, A2 => n25964, ZN => n19283);
   U275 : INV_X1 port map( A => n27040, ZN => n1825);
   U276 : INV_X1 port map( A => DATA2(5), ZN => n27276);
   U277 : NAND4_X1 port map( A1 => n27077, A2 => n27276, A3 => FUNC(2), A4 => 
                           FUNC(1), ZN => n27041);
   U278 : INV_X1 port map( A => n27041, ZN => n25966);
   U279 : INV_X1 port map( A => DATA2(2), ZN => n27592);
   U280 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(4), ZN => n27590);
   U281 : NOR2_X1 port map( A1 => n27592, A2 => n27590, ZN => n27578);
   U282 : NAND2_X1 port map( A1 => n27575, A2 => n27578, ZN => n27042);
   U283 : NAND2_X1 port map( A1 => n25966, A2 => n27042, ZN => n26145);
   U284 : NOR2_X1 port map( A1 => FUNC(3), A2 => n26145, ZN => n1831);
   U285 : AOI21_X1 port map( B1 => DATA2(1), B2 => DATA2(2), A => n25968, ZN =>
                           n25967);
   U286 : INV_X1 port map( A => n25967, ZN => n26209);
   U287 : OAI21_X1 port map( B1 => DATA2(0), B2 => n25968, A => n26209, ZN => 
                           n26795);
   U288 : CLKBUF_X1 port map( A => n26795, Z => n27624);
   U289 : INV_X1 port map( A => n26166, ZN => n27593);
   U290 : NAND3_X1 port map( A1 => DATA2(3), A2 => n1863, A3 => n27592, ZN => 
                           n25989);
   U291 : NOR2_X1 port map( A1 => n27593, A2 => n25989, ZN => n1857);
   U292 : INV_X1 port map( A => n25968, ZN => n25977);
   U293 : OAI21_X1 port map( B1 => n27571, B2 => n27594, A => n26014, ZN => 
                           n25969);
   U294 : INV_X1 port map( A => n25969, ZN => n26425);
   U295 : INV_X1 port map( A => n26425, ZN => n27645);
   U296 : INV_X1 port map( A => n27638, ZN => n27709);
   U297 : NAND2_X1 port map( A1 => DATA2(0), A2 => n27571, ZN => n27579);
   U298 : OR2_X1 port map( A1 => n26478, A2 => n27579, ZN => n26415);
   U299 : INV_X1 port map( A => n26415, ZN => n26848);
   U300 : INV_X1 port map( A => n27575, ZN => n27591);
   U301 : INV_X1 port map( A => n26753, ZN => n26722);
   U302 : NOR2_X1 port map( A1 => n24047, A2 => n26722, ZN => n26021);
   U303 : INV_X1 port map( A => n26478, ZN => n26750);
   U304 : NOR2_X1 port map( A1 => n24055, A2 => n26750, ZN => n26036);
   U305 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(9), A => n26021, B => 
                           n26036, ZN => n25970);
   U306 : NAND3_X1 port map( A1 => DATA2(1), A2 => n26750, A3 => n27573, ZN => 
                           n26707);
   U307 : INV_X1 port map( A => n26707, ZN => n26724);
   U308 : NAND2_X1 port map( A1 => n24181, A2 => n26724, ZN => n26031);
   U309 : OAI211_X1 port map( C1 => n26666, C2 => n27151, A => n25970, B => 
                           n26031, ZN => n25971);
   U310 : INV_X1 port map( A => n25971, ZN => n25984);
   U311 : NOR2_X1 port map( A1 => n25975, A2 => n26722, ZN => n26034);
   U312 : NOR2_X1 port map( A1 => n24046, A2 => n26461, ZN => n26022);
   U313 : AOI211_X1 port map( C1 => n26724, C2 => DATA1(10), A => n26034, B => 
                           n26022, ZN => n25972);
   U314 : INV_X1 port map( A => n26415, ZN => n26704);
   U315 : NAND2_X1 port map( A1 => DATA1(11), A2 => n26704, ZN => n26079);
   U316 : OAI211_X1 port map( C1 => n26666, C2 => n27547, A => n25972, B => 
                           n26079, ZN => n25973);
   U317 : INV_X1 port map( A => n25973, ZN => n26008);
   U318 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(0), ZN => n26117);
   U319 : NAND2_X1 port map( A1 => n26446, A2 => n26117, ZN => n26794);
   U320 : INV_X1 port map( A => n26207, ZN => n26769);
   U321 : INV_X1 port map( A => n26666, ZN => n26847);
   U322 : NOR2_X1 port map( A1 => n24046, A2 => n26722, ZN => n26026);
   U323 : NOR2_X1 port map( A1 => n24047, A2 => n26750, ZN => n26046);
   U324 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(10), A => n26026, B => 
                           n26046, ZN => n25974);
   U325 : INV_X1 port map( A => n25974, ZN => n25976);
   U326 : NOR2_X1 port map( A1 => n25975, A2 => n26707, ZN => n26065);
   U327 : AOI211_X1 port map( C1 => n26847, C2 => DATA1(11), A => n25976, B => 
                           n26065, ZN => n26007);
   U328 : INV_X1 port map( A => n27579, ZN => n27580);
   U329 : AND3_X1 port map( A1 => DATA2(2), A2 => n25977, A3 => n27580, ZN => 
                           n26205);
   U330 : INV_X1 port map( A => n26205, ZN => n26754);
   U331 : OAI222_X1 port map( A1 => n25984, A2 => n26446, B1 => n26008, B2 => 
                           n26769, C1 => n26007, C2 => n26754, ZN => n26122);
   U332 : INV_X1 port map( A => n26122, ZN => n26167);
   U333 : INV_X1 port map( A => n26205, ZN => n26792);
   U334 : NOR2_X1 port map( A1 => n24047, A2 => n26707, ZN => n26027);
   U335 : CLKBUF_X1 port map( A => n26847, Z => n26719);
   U336 : NAND2_X1 port map( A1 => DATA1(9), A2 => n26719, ZN => n26069);
   U337 : NOR2_X1 port map( A1 => n26722, A2 => n24077, ZN => n26047);
   U338 : INV_X1 port map( A => n26047, ZN => n25978);
   U339 : OAI211_X1 port map( C1 => n24056, C2 => n26750, A => n26069, B => 
                           n25978, ZN => n25979);
   U340 : AOI211_X1 port map( C1 => n26704, C2 => n24181, A => n26027, B => 
                           n25979, ZN => n25986);
   U341 : OAI222_X1 port map( A1 => n26794, A2 => n26007, B1 => n26792, B2 => 
                           n25984, C1 => n26446, C2 => n25986, ZN => n26118);
   U342 : AND2_X1 port map( A1 => n24178, A2 => n26724, ZN => n26023);
   U343 : NOR2_X1 port map( A1 => n26666, A2 => n24046, ZN => n26060);
   U344 : INV_X1 port map( A => n26060, ZN => n25980);
   U345 : NAND2_X1 port map( A1 => n24177, A2 => n26753, ZN => n26035);
   U346 : OAI211_X1 port map( C1 => n24054, C2 => n26750, A => n25980, B => 
                           n26035, ZN => n25981);
   U347 : AOI211_X1 port map( C1 => n26848, C2 => n24179, A => n26023, B => 
                           n25981, ZN => n25985);
   U348 : NOR2_X1 port map( A1 => n24077, A2 => n26415, ZN => n26028);
   U349 : NOR2_X1 port map( A1 => n24054, A2 => n26722, ZN => n26042);
   U350 : NOR2_X1 port map( A1 => n24056, A2 => n26707, ZN => n26048);
   U351 : OAI22_X1 port map( A1 => n24047, A2 => n26666, B1 => n24164, B2 => 
                           n26750, ZN => n25982);
   U352 : NOR4_X1 port map( A1 => n26028, A2 => n26042, A3 => n26048, A4 => 
                           n25982, ZN => n26232);
   U353 : NOR2_X1 port map( A1 => n24055, A2 => n26666, ZN => n26029);
   U354 : NAND2_X1 port map( A1 => n24177, A2 => n26704, ZN => n26019);
   U355 : NAND2_X1 port map( A1 => n24048, A2 => n26753, ZN => n26039);
   U356 : OAI211_X1 port map( C1 => n24054, C2 => n26707, A => n26019, B => 
                           n26039, ZN => n25983);
   U357 : AOI211_X1 port map( C1 => n24049, C2 => n26478, A => n26029, B => 
                           n25983, ZN => n26231);
   U358 : OAI222_X1 port map( A1 => n26794, A2 => n25985, B1 => n26792, B2 => 
                           n26232, C1 => n26446, C2 => n26231, ZN => n26309);
   U359 : AOI22_X1 port map( A1 => n25892, A2 => n26118, B1 => n26309, B2 => 
                           n27645, ZN => n25988);
   U360 : OAI222_X1 port map( A1 => n26794, A2 => n25984, B1 => n26792, B2 => 
                           n25986, C1 => n26446, C2 => n25985, ZN => n26168);
   U361 : OAI222_X1 port map( A1 => n26769, A2 => n25986, B1 => n26792, B2 => 
                           n25985, C1 => n26446, C2 => n26232, ZN => n26493);
   U362 : AOI22_X1 port map( A1 => n1857, A2 => n26168, B1 => n27709, B2 => 
                           n26493, ZN => n25987);
   U363 : OAI211_X1 port map( C1 => n27641, C2 => n26167, A => n25988, B => 
                           n25987, ZN => n1822);
   U364 : NOR2_X1 port map( A1 => n27591, A2 => n25989, ZN => n1843);
   U365 : INV_X1 port map( A => n1843, ZN => n1856);
   U366 : NOR2_X1 port map( A1 => n26461, A2 => n26977, ZN => n26071);
   U367 : NOR2_X1 port map( A1 => n26964, A2 => n26722, ZN => n26086);
   U368 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(16), A => n26071, B => 
                           n26086, ZN => n25990);
   U369 : NAND2_X1 port map( A1 => DATA1(15), A2 => n26724, ZN => n26100);
   U370 : OAI211_X1 port map( C1 => n26666, C2 => n26915, A => n25990, B => 
                           n26100, ZN => n26001);
   U371 : INV_X1 port map( A => DATA1(18), ZN => n26903);
   U372 : NOR2_X1 port map( A1 => n26461, A2 => n26943, ZN => n26085);
   U373 : INV_X1 port map( A => DATA1(16), ZN => n26930);
   U374 : NOR2_X1 port map( A1 => n26930, A2 => n26722, ZN => n26098);
   U375 : AOI211_X1 port map( C1 => n26724, C2 => DATA1(17), A => n26085, B => 
                           n26098, ZN => n25991);
   U376 : NAND2_X1 port map( A1 => DATA1(19), A2 => n26719, ZN => n26140);
   U377 : OAI211_X1 port map( C1 => n26415, C2 => n26903, A => n25991, B => 
                           n26140, ZN => n26202);
   U378 : INV_X1 port map( A => n26794, ZN => n26207);
   U379 : NOR2_X1 port map( A1 => n26461, A2 => n26964, ZN => n26075);
   U380 : NOR2_X1 port map( A1 => n26943, A2 => n26722, ZN => n26096);
   U381 : AOI211_X1 port map( C1 => n26704, C2 => DATA1(17), A => n26075, B => 
                           n26096, ZN => n25992);
   U382 : NAND2_X1 port map( A1 => DATA1(16), A2 => n26724, ZN => n26103);
   U383 : OAI211_X1 port map( C1 => n26666, C2 => n26903, A => n25992, B => 
                           n26103, ZN => n26199);
   U384 : AOI222_X1 port map( A1 => n26001, A2 => n26209, B1 => n26202, B2 => 
                           n26207, C1 => n26199, C2 => n26205, ZN => n1846);
   U385 : NOR2_X1 port map( A1 => n26461, A2 => n27547, ZN => n26059);
   U386 : NOR2_X1 port map( A1 => n26977, A2 => n26722, ZN => n26076);
   U387 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(15), A => n26059, B => 
                           n26076, ZN => n25993);
   U388 : NAND2_X1 port map( A1 => DATA1(14), A2 => n26724, ZN => n26093);
   U389 : OAI211_X1 port map( C1 => n26666, C2 => n26930, A => n25993, B => 
                           n26093, ZN => n26000);
   U390 : AOI222_X1 port map( A1 => n26000, A2 => n26209, B1 => n26199, B2 => 
                           n26207, C1 => n26001, C2 => n26205, ZN => n1848);
   U391 : NOR2_X1 port map( A1 => n27547, A2 => n26707, ZN => n26077);
   U392 : NAND2_X1 port map( A1 => DATA1(11), A2 => n26753, ZN => n26061);
   U393 : NAND2_X1 port map( A1 => DATA1(10), A2 => n26478, ZN => n26030);
   U394 : OAI211_X1 port map( C1 => n26415, C2 => n26977, A => n26061, B => 
                           n26030, ZN => n25994);
   U395 : AOI211_X1 port map( C1 => n26719, C2 => DATA1(14), A => n26077, B => 
                           n25994, ZN => n26006);
   U396 : INV_X1 port map( A => n26006, ZN => n25997);
   U397 : NOR2_X1 port map( A1 => n27547, A2 => n26722, ZN => n26070);
   U398 : NOR2_X1 port map( A1 => n26461, A2 => n25995, ZN => n26064);
   U399 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(14), A => n26070, B => 
                           n26064, ZN => n25996);
   U400 : NAND2_X1 port map( A1 => DATA1(13), A2 => n26724, ZN => n26087);
   U401 : OAI211_X1 port map( C1 => n26666, C2 => n26943, A => n25996, B => 
                           n26087, ZN => n26002);
   U402 : AOI222_X1 port map( A1 => n25997, A2 => n26209, B1 => n26000, B2 => 
                           n26207, C1 => n26002, C2 => n26205, ZN => n26237);
   U403 : INV_X1 port map( A => n26237, ZN => n26005);
   U404 : NOR2_X1 port map( A1 => n27151, A2 => n26722, ZN => n26066);
   U405 : NAND2_X1 port map( A1 => DATA1(11), A2 => n26724, ZN => n26073);
   U406 : NAND2_X1 port map( A1 => DATA1(9), A2 => n26478, ZN => n26024);
   U407 : OAI211_X1 port map( C1 => n26415, C2 => n27547, A => n26073, B => 
                           n26024, ZN => n25998);
   U408 : AOI211_X1 port map( C1 => n26847, C2 => DATA1(13), A => n26066, B => 
                           n25998, ZN => n26009);
   U409 : OAI22_X1 port map( A1 => n26009, A2 => n26446, B1 => n26006, B2 => 
                           n26754, ZN => n25999);
   U410 : AOI21_X1 port map( B1 => n26207, B2 => n26002, A => n25999, ZN => 
                           n26236);
   U411 : AOI222_X1 port map( A1 => n26002, A2 => n26209, B1 => n26001, B2 => 
                           n26207, C1 => n26000, C2 => n26205, ZN => n26238);
   U412 : CLKBUF_X1 port map( A => n1857, Z => n27632);
   U413 : INV_X1 port map( A => n27632, ZN => n27636);
   U414 : OAI22_X1 port map( A1 => n26425, A2 => n26236, B1 => n26238, B2 => 
                           n27636, ZN => n26004);
   U415 : INV_X1 port map( A => n25892, ZN => n27607);
   U416 : OAI22_X1 port map( A1 => n27641, A2 => n1846, B1 => n1848, B2 => 
                           n27607, ZN => n26003);
   U417 : AOI211_X1 port map( C1 => n27709, C2 => n26005, A => n26004, B => 
                           n26003, ZN => n1847);
   U418 : OAI222_X1 port map( A1 => n26794, A2 => n26006, B1 => n26792, B2 => 
                           n26009, C1 => n26446, C2 => n26008, ZN => n26241);
   U419 : OAI222_X1 port map( A1 => n26794, A2 => n26009, B1 => n26792, B2 => 
                           n26008, C1 => n26446, C2 => n26007, ZN => n26114);
   U420 : INV_X1 port map( A => n26114, ZN => n26169);
   U421 : OAI22_X1 port map( A1 => n26169, A2 => n27638, B1 => n26236, B2 => 
                           n27607, ZN => n26011);
   U422 : OAI22_X1 port map( A1 => n27641, A2 => n26237, B1 => n26425, B2 => 
                           n26167, ZN => n26010);
   U423 : AOI211_X1 port map( C1 => n1857, C2 => n26241, A => n26011, B => 
                           n26010, ZN => n1823);
   U424 : OAI22_X1 port map( A1 => n1856, A2 => n1847, B1 => n1836, B2 => n1823
                           , ZN => n26012);
   U425 : INV_X1 port map( A => n26012, ZN => n19003);
   U426 : AOI21_X1 port map( B1 => DATA2(3), B2 => n27575, A => n26013, ZN => 
                           n1858);
   U427 : INV_X1 port map( A => n1836, ZN => n1860);
   U428 : INV_X1 port map( A => n26117, ZN => n26015);
   U429 : NOR3_X2 port map( A1 => n26015, A2 => n26014, A3 => n1860, ZN => 
                           n1861);
   U430 : INV_X1 port map( A => n1861, ZN => n1896);
   U431 : OAI22_X1 port map( A1 => n26236, A2 => n27636, B1 => n26237, B2 => 
                           n27607, ZN => n26017);
   U432 : OAI22_X1 port map( A1 => n27641, A2 => n26238, B1 => n26425, B2 => 
                           n26169, ZN => n26016);
   U433 : AOI211_X1 port map( C1 => n27709, C2 => n26241, A => n26017, B => 
                           n26016, ZN => n1828);
   U434 : INV_X1 port map( A => n1858, ZN => n27564);
   U435 : OAI22_X1 port map( A1 => n27564, A2 => n1847, B1 => n1896, B2 => 
                           n1828, ZN => n26018);
   U436 : INV_X1 port map( A => n26018, ZN => n19005);
   U437 : NAND2_X1 port map( A1 => n24176, A2 => n26719, ZN => n26228);
   U438 : NAND2_X1 port map( A1 => n26019, A2 => n26228, ZN => n26020);
   U439 : NOR4_X1 port map( A1 => n26023, A2 => n26022, A3 => n26021, A4 => 
                           n26020, ZN => n26045);
   U440 : NAND2_X1 port map( A1 => n24177, A2 => n26719, ZN => n26224);
   U441 : NAND2_X1 port map( A1 => n26224, A2 => n26024, ZN => n26025);
   U442 : NOR4_X1 port map( A1 => n26028, A2 => n26027, A3 => n26026, A4 => 
                           n26025, ZN => n26051);
   U443 : INV_X1 port map( A => n26029, ZN => n26032);
   U444 : NAND3_X1 port map( A1 => n26032, A2 => n26031, A3 => n26030, ZN => 
                           n26033);
   U445 : AOI211_X1 port map( C1 => n26704, C2 => n24179, A => n26034, B => 
                           n26033, ZN => n26063);
   U446 : OAI222_X1 port map( A1 => n26769, A2 => n26045, B1 => n26792, B2 => 
                           n26051, C1 => n26446, C2 => n26063, ZN => n22526);
   U447 : INV_X1 port map( A => n26035, ZN => n26037);
   U448 : AOI211_X1 port map( C1 => n26724, C2 => n24176, A => n26037, B => 
                           n26036, ZN => n26038);
   U449 : NAND2_X1 port map( A1 => n24048, A2 => n26704, ZN => n26227);
   U450 : OAI211_X1 port map( C1 => n24165, C2 => n26666, A => n26038, B => 
                           n26227, ZN => n26053);
   U451 : NOR2_X1 port map( A1 => n24165, A2 => n26707, ZN => n26230);
   U452 : AND2_X1 port map( A1 => n24175, A2 => n26848, ZN => n26667);
   U453 : AOI211_X1 port map( C1 => n26847, C2 => n24173, A => n26230, B => 
                           n26667, ZN => n26040);
   U454 : OAI211_X1 port map( C1 => n24054, C2 => n26750, A => n26040, B => 
                           n26039, ZN => n26044);
   U455 : NOR2_X1 port map( A1 => n24056, A2 => n26461, ZN => n26041);
   U456 : AOI211_X1 port map( C1 => n26847, C2 => n24175, A => n26042, B => 
                           n26041, ZN => n26043);
   U457 : NAND2_X1 port map( A1 => n24048, A2 => n26724, ZN => n26223);
   U458 : OAI211_X1 port map( C1 => n24165, C2 => n26415, A => n26043, B => 
                           n26223, ZN => n26054);
   U459 : AOI222_X1 port map( A1 => n26053, A2 => n26209, B1 => n26044, B2 => 
                           n26207, C1 => n26054, C2 => n26205, ZN => n26050);
   U460 : INV_X1 port map( A => n26045, ZN => n26052);
   U461 : NOR2_X1 port map( A1 => n24054, A2 => n26415, ZN => n26226);
   U462 : NOR4_X1 port map( A1 => n26048, A2 => n26226, A3 => n26047, A4 => 
                           n26046, ZN => n26049);
   U463 : OAI21_X1 port map( B1 => n27682, B2 => n26666, A => n26049, ZN => 
                           n26055);
   U464 : AOI222_X1 port map( A1 => n26052, A2 => n26209, B1 => n26053, B2 => 
                           n26207, C1 => n26055, C2 => n26205, ZN => n26854);
   U465 : OAI22_X1 port map( A1 => n27641, A2 => n26050, B1 => n26854, B2 => 
                           n27636, ZN => n26057);
   U466 : INV_X1 port map( A => n26051, ZN => n26083);
   U467 : AOI222_X1 port map( A1 => n26083, A2 => n26209, B1 => n26055, B2 => 
                           n26207, C1 => n26052, C2 => n26205, ZN => n26853);
   U468 : AOI222_X1 port map( A1 => n26055, A2 => n26209, B1 => n26054, B2 => 
                           n26207, C1 => n26053, C2 => n26205, ZN => n26852);
   U469 : OAI22_X1 port map( A1 => n26853, A2 => n27638, B1 => n26852, B2 => 
                           n27607, ZN => n26056);
   U470 : AOI211_X1 port map( C1 => n27645, C2 => n22526, A => n26057, B => 
                           n26056, ZN => n26058);
   U471 : INV_X1 port map( A => n26058, ZN => n18902);
   U472 : INV_X1 port map( A => DATA1(30), ZN => n27205);
   U473 : XOR2_X1 port map( A => DATA2_I_30_port, B => n27205, Z => n26517);
   U474 : INV_X1 port map( A => n26517, ZN => n1814);
   U475 : INV_X1 port map( A => DATA1(0), ZN => n1855);
   U476 : INV_X1 port map( A => DATA1(1), ZN => n1854);
   U477 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(9), A => n26060, B => 
                           n26059, ZN => n26062);
   U478 : OAI211_X1 port map( C1 => n26707, C2 => n27151, A => n26062, B => 
                           n26061, ZN => n26081);
   U479 : INV_X1 port map( A => n26063, ZN => n26082);
   U480 : NOR2_X1 port map( A1 => n24047, A2 => n26666, ZN => n26067);
   U481 : NOR4_X1 port map( A1 => n26067, A2 => n26066, A3 => n26065, A4 => 
                           n26064, ZN => n26068);
   U482 : OAI21_X1 port map( B1 => n24046, B2 => n26415, A => n26068, ZN => 
                           n26084);
   U483 : AOI222_X1 port map( A1 => n26081, A2 => n26209, B1 => n26082, B2 => 
                           n26207, C1 => n26084, C2 => n26205, ZN => n27640);
   U484 : INV_X1 port map( A => n27640, ZN => n26092);
   U485 : INV_X1 port map( A => n26069, ZN => n26072);
   U486 : NOR3_X1 port map( A1 => n26072, A2 => n26071, A3 => n26070, ZN => 
                           n26074);
   U487 : OAI211_X1 port map( C1 => n26415, C2 => n27151, A => n26074, B => 
                           n26073, ZN => n26089);
   U488 : AOI222_X1 port map( A1 => n26089, A2 => n26209, B1 => n26084, B2 => 
                           n26207, C1 => n26081, C2 => n26205, ZN => n27635);
   U489 : NOR2_X1 port map( A1 => n27151, A2 => n26666, ZN => n26078);
   U490 : NOR4_X1 port map( A1 => n26078, A2 => n26077, A3 => n26076, A4 => 
                           n26075, ZN => n26080);
   U491 : NAND2_X1 port map( A1 => n26080, A2 => n26079, ZN => n26105);
   U492 : AOI222_X1 port map( A1 => n26105, A2 => n26209, B1 => n26081, B2 => 
                           n26207, C1 => n26089, C2 => n26205, ZN => n27637);
   U493 : OAI22_X1 port map( A1 => n27636, A2 => n27635, B1 => n27638, B2 => 
                           n27637, ZN => n26091);
   U494 : AOI222_X1 port map( A1 => n26084, A2 => n26209, B1 => n26083, B2 => 
                           n26207, C1 => n26082, C2 => n26205, ZN => n26857);
   U495 : AOI211_X1 port map( C1 => n26719, C2 => DATA1(11), A => n26086, B => 
                           n26085, ZN => n26088);
   U496 : OAI211_X1 port map( C1 => n26415, C2 => n27547, A => n26088, B => 
                           n26087, ZN => n26107);
   U497 : AOI222_X1 port map( A1 => n26107, A2 => n26209, B1 => n26089, B2 => 
                           n26207, C1 => n26105, C2 => n26205, ZN => n27639);
   U498 : OAI22_X1 port map( A1 => n27641, A2 => n26857, B1 => n26425, B2 => 
                           n27639, ZN => n26090);
   U499 : AOI211_X1 port map( C1 => n26092, C2 => n25892, A => n26091, B => 
                           n26090, ZN => n26860);
   U500 : INV_X1 port map( A => n26860, ZN => n1819);
   U501 : NAND2_X1 port map( A1 => DATA1(12), A2 => n26719, ZN => n26094);
   U502 : OAI211_X1 port map( C1 => n26750, C2 => n26930, A => n26094, B => 
                           n26093, ZN => n26095);
   U503 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(13), A => n26096, B => 
                           n26095, ZN => n26097);
   U504 : INV_X1 port map( A => n26097, ZN => n26106);
   U505 : NOR2_X1 port map( A1 => n26977, A2 => n26666, ZN => n26099);
   U506 : AOI211_X1 port map( C1 => DATA1(17), C2 => n26478, A => n26099, B => 
                           n26098, ZN => n26101);
   U507 : OAI211_X1 port map( C1 => n26415, C2 => n26964, A => n26101, B => 
                           n26100, ZN => n26111);
   U508 : NOR2_X1 port map( A1 => n26943, A2 => n26415, ZN => n26102);
   U509 : NOR2_X1 port map( A1 => n26915, A2 => n26722, ZN => n26198);
   U510 : AOI211_X1 port map( C1 => DATA1(18), C2 => n26478, A => n26102, B => 
                           n26198, ZN => n26104);
   U511 : OAI211_X1 port map( C1 => n26666, C2 => n26964, A => n26104, B => 
                           n26103, ZN => n26128);
   U512 : AOI222_X1 port map( A1 => n26207, A2 => n26106, B1 => n26205, B2 => 
                           n26111, C1 => n26209, C2 => n26128, ZN => n26129);
   U513 : INV_X1 port map( A => n26129, ZN => n27625);
   U514 : AOI222_X1 port map( A1 => n26106, A2 => n26209, B1 => n26105, B2 => 
                           n26207, C1 => n26107, C2 => n26205, ZN => n27628);
   U515 : AOI222_X1 port map( A1 => n26111, A2 => n26209, B1 => n26107, B2 => 
                           n26207, C1 => n26106, C2 => n26205, ZN => n26247);
   U516 : OAI22_X1 port map( A1 => n27628, A2 => n27607, B1 => n26247, B2 => 
                           n27636, ZN => n26113);
   U517 : NOR2_X1 port map( A1 => n26930, A2 => n26415, ZN => n26110);
   U518 : NAND2_X1 port map( A1 => DATA1(15), A2 => n26719, ZN => n26108);
   U519 : NAND2_X1 port map( A1 => DATA1(19), A2 => n26478, ZN => n26216);
   U520 : OAI211_X1 port map( C1 => n26722, C2 => n26903, A => n26108, B => 
                           n26216, ZN => n26109);
   U521 : AOI211_X1 port map( C1 => n26724, C2 => DATA1(17), A => n26110, B => 
                           n26109, ZN => n26135);
   U522 : INV_X1 port map( A => n26135, ZN => n26127);
   U523 : AOI222_X1 port map( A1 => n26127, A2 => n26209, B1 => n26111, B2 => 
                           n26207, C1 => n26128, C2 => n26205, ZN => n26251);
   U524 : OAI22_X1 port map( A1 => n27641, A2 => n27639, B1 => n26425, B2 => 
                           n26251, ZN => n26112);
   U525 : AOI211_X1 port map( C1 => n27709, C2 => n27625, A => n26113, B => 
                           n26112, ZN => n1845);
   U526 : AOI22_X1 port map( A1 => n25892, A2 => n26114, B1 => n26795, B2 => 
                           n26241, ZN => n26116);
   U527 : AOI22_X1 port map( A1 => n27709, A2 => n26118, B1 => n27645, B2 => 
                           n26168, ZN => n26115);
   U528 : OAI211_X1 port map( C1 => n26167, C2 => n27636, A => n26116, B => 
                           n26115, ZN => n1821);
   U529 : NOR3_X1 port map( A1 => n1860, A2 => n26117, A3 => n27594, ZN => 
                           n1894);
   U530 : INV_X1 port map( A => n1894, ZN => n1859);
   U531 : OAI22_X1 port map( A1 => n27636, A2 => n26169, B1 => n27641, B2 => 
                           n26236, ZN => n26121);
   U532 : INV_X1 port map( A => n26241, ZN => n26119);
   U533 : INV_X1 port map( A => n26118, ZN => n26487);
   U534 : OAI22_X1 port map( A1 => n27607, A2 => n26119, B1 => n26425, B2 => 
                           n26487, ZN => n26120);
   U535 : AOI211_X1 port map( C1 => n26122, C2 => n27709, A => n26121, B => 
                           n26120, ZN => n26485);
   U536 : OAI22_X1 port map( A1 => n1836, A2 => n26485, B1 => n1859, B2 => 
                           n1823, ZN => n26123);
   U537 : INV_X1 port map( A => n26123, ZN => n19004);
   U538 : INV_X1 port map( A => DATA1(4), ZN => n1853);
   U539 : NOR2_X1 port map( A1 => n26930, A2 => n26666, ZN => n26126);
   U540 : INV_X1 port map( A => DATA1(20), ZN => n26833);
   U541 : NAND2_X1 port map( A1 => DATA1(17), A2 => n26704, ZN => n26124);
   U542 : NAND2_X1 port map( A1 => DATA1(19), A2 => n26753, ZN => n26186);
   U543 : OAI211_X1 port map( C1 => n26750, C2 => n26833, A => n26124, B => 
                           n26186, ZN => n26125);
   U544 : AOI211_X1 port map( C1 => n26724, C2 => DATA1(18), A => n26126, B => 
                           n26125, ZN => n26134);
   U545 : INV_X1 port map( A => n26134, ZN => n26139);
   U546 : AOI222_X1 port map( A1 => n26139, A2 => n26209, B1 => n26128, B2 => 
                           n26207, C1 => n26127, C2 => n26205, ZN => n27603);
   U547 : INV_X1 port map( A => n27603, ZN => n26248);
   U548 : OAI22_X1 port map( A1 => n26251, A2 => n27638, B1 => n26129, B2 => 
                           n27636, ZN => n26131);
   U549 : OAI22_X1 port map( A1 => n27641, A2 => n27628, B1 => n26247, B2 => 
                           n27607, ZN => n26130);
   U550 : AOI211_X1 port map( C1 => n27645, C2 => n26248, A => n26131, B => 
                           n26130, ZN => n1844);
   U551 : INV_X1 port map( A => DATA1(23), ZN => n1840);
   U552 : NOR2_X1 port map( A1 => n26915, A2 => n26666, ZN => n26133);
   U553 : INV_X1 port map( A => DATA1(21), ZN => n27653);
   U554 : NAND2_X1 port map( A1 => DATA1(19), A2 => n26724, ZN => n26189);
   U555 : NAND2_X1 port map( A1 => DATA1(20), A2 => n26753, ZN => n26215);
   U556 : OAI211_X1 port map( C1 => n26750, C2 => n27653, A => n26189, B => 
                           n26215, ZN => n26132);
   U557 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(18), A => n26133, B => 
                           n26132, ZN => n26138);
   U558 : OAI222_X1 port map( A1 => n26794, A2 => n26135, B1 => n26792, B2 => 
                           n26134, C1 => n26446, C2 => n26138, ZN => n27600);
   U559 : AND2_X1 port map( A1 => DATA1(19), A2 => n26848, ZN => n26197);
   U560 : NOR2_X1 port map( A1 => n27653, A2 => n26722, ZN => n26442);
   U561 : AOI211_X1 port map( C1 => DATA1(22), C2 => n26478, A => n26197, B => 
                           n26442, ZN => n26137);
   U562 : NAND2_X1 port map( A1 => DATA1(18), A2 => n26719, ZN => n26136);
   U563 : OAI211_X1 port map( C1 => n26707, C2 => n26833, A => n26137, B => 
                           n26136, ZN => n26208);
   U564 : INV_X1 port map( A => n26138, ZN => n26142);
   U565 : AOI222_X1 port map( A1 => n26208, A2 => n26209, B1 => n26139, B2 => 
                           n26207, C1 => n26142, C2 => n26205, ZN => n27597);
   U566 : OAI22_X1 port map( A1 => n27597, A2 => n27638, B1 => n27603, B2 => 
                           n27607, ZN => n26144);
   U567 : NOR2_X1 port map( A1 => n26833, A2 => n26415, ZN => n26192);
   U568 : NOR2_X1 port map( A1 => n26461, A2 => n1840, ZN => n26471);
   U569 : AOI211_X1 port map( C1 => n26724, C2 => DATA1(21), A => n26192, B => 
                           n26471, ZN => n26141);
   U570 : OAI211_X1 port map( C1 => n26722, C2 => n27177, A => n26141, B => 
                           n26140, ZN => n26206);
   U571 : AOI222_X1 port map( A1 => n26206, A2 => n26209, B1 => n26142, B2 => 
                           n26207, C1 => n26208, C2 => n26205, ZN => n27596);
   U572 : OAI22_X1 port map( A1 => n27641, A2 => n26251, B1 => n26425, B2 => 
                           n27596, ZN => n26143);
   U573 : AOI211_X1 port map( C1 => n1857, C2 => n27600, A => n26144, B => 
                           n26143, ZN => n1842);
   U574 : NOR2_X1 port map( A1 => n1832, A2 => n26145, ZN => n1830);
   U575 : INV_X2 port map( A => data1_mul_0_port, ZN => n1807);
   U576 : INV_X1 port map( A => n9084, ZN => n1805);
   U577 : INV_X1 port map( A => n9081, ZN => n1804);
   U578 : INV_X1 port map( A => n9078, ZN => n1803);
   U579 : INV_X1 port map( A => n9072, ZN => n1800);
   U580 : INV_X1 port map( A => n9069, ZN => n1799);
   U581 : INV_X1 port map( A => n9066, ZN => n1798);
   U582 : INV_X1 port map( A => n9063, ZN => n1797);
   U583 : INV_X1 port map( A => n9057, ZN => n1795);
   U584 : INV_X1 port map( A => n9054, ZN => n1794);
   U585 : INV_X1 port map( A => n9051, ZN => n1793);
   U586 : INV_X1 port map( A => n9048, ZN => n1792);
   U587 : INV_X1 port map( A => DATA1(6), ZN => n1851);
   U588 : INV_X1 port map( A => DATA1(5), ZN => n1852);
   U589 : OR4_X1 port map( A1 => DATA1(5), A2 => DATA1(4), A3 => DATA1(0), A4 
                           => DATA1(3), ZN => n19010);
   U590 : INV_X1 port map( A => DATA1(8), ZN => n1849);
   U591 : INV_X1 port map( A => DATA1(7), ZN => n1850);
   U592 : NAND2_X1 port map( A1 => n24044, A2 => n25872, ZN => n27474);
   U593 : OAI21_X1 port map( B1 => n24044, B2 => n25872, A => n27474, ZN => 
                           n22802);
   U594 : AOI211_X1 port map( C1 => n24107, C2 => n24116, A => n23699, B => 
                           n23735, ZN => n26152);
   U595 : AOI211_X1 port map( C1 => n24117, C2 => n24107, A => n23696, B => 
                           n23733, ZN => n26955);
   U596 : AOI211_X1 port map( C1 => n24116, C2 => n24058, A => n23697, B => 
                           n23734, ZN => n26153);
   U597 : OAI222_X1 port map( A1 => n24168, A2 => n26152, B1 => n24081, B2 => 
                           n26955, C1 => n23979, C2 => n26153, ZN => n26923);
   U598 : OAI211_X1 port map( C1 => n24158, C2 => n23736, A => n23739, B => 
                           n23738, ZN => n26146);
   U599 : INV_X1 port map( A => n26146, ZN => n26159);
   U600 : OAI22_X1 port map( A1 => n23954, A2 => n24136, B1 => n24156, B2 => 
                           n23736, ZN => n26147);
   U601 : AOI211_X1 port map( C1 => n24106, C2 => n24116, A => n23700, B => 
                           n26147, ZN => n26154);
   U602 : OAI222_X1 port map( A1 => n24168, A2 => n26159, B1 => n24081, B2 => 
                           n26152, C1 => n23979, C2 => n26154, ZN => n26611);
   U603 : INV_X1 port map( A => n26611, ZN => n26893);
   U604 : AOI22_X1 port map( A1 => n24058, A2 => n24117, B1 => n24107, B2 => 
                           n23751, ZN => n26148);
   U605 : OAI211_X1 port map( C1 => n23957, C2 => n23743, A => n25863, B => 
                           n26148, ZN => n26971);
   U606 : OAI22_X1 port map( A1 => n24168, A2 => n26153, B1 => n23979, B2 => 
                           n26955, ZN => n26149);
   U607 : AOI21_X1 port map( B1 => n27670, B2 => n26971, A => n26149, ZN => 
                           n26924);
   U608 : OAI22_X1 port map( A1 => n26893, A2 => n27676, B1 => n26924, B2 => 
                           n27664, ZN => n26156);
   U609 : AOI211_X1 port map( C1 => n24154, C2 => n23600, A => n23747, B => 
                           n23746, ZN => n26536);
   U610 : OAI22_X1 port map( A1 => n26536, A2 => n24156, B1 => n24151, B2 => 
                           n24119, ZN => n26151);
   U611 : OAI21_X1 port map( B1 => n23736, B2 => n23953, A => n23737, ZN => 
                           n26150);
   U612 : NOR2_X1 port map( A1 => n26151, A2 => n26150, ZN => n26543);
   U613 : OAI222_X1 port map( A1 => n24168, A2 => n26543, B1 => n24081, B2 => 
                           n26154, C1 => n23979, C2 => n26159, ZN => n26604);
   U614 : INV_X1 port map( A => n26604, ZN => n26616);
   U615 : OAI222_X1 port map( A1 => n24168, A2 => n26154, B1 => n24081, B2 => 
                           n26153, C1 => n23979, C2 => n26152, ZN => n26910);
   U616 : INV_X1 port map( A => n26910, ZN => n26892);
   U617 : OAI22_X1 port map( A1 => n24113, A2 => n26616, B1 => n26892, B2 => 
                           n27672, ZN => n26155);
   U618 : AOI211_X1 port map( C1 => n24104, C2 => n26923, A => n26156, B => 
                           n26155, ZN => n26822);
   U619 : INV_X1 port map( A => n26822, ZN => n26841);
   U620 : OAI22_X1 port map( A1 => n23954, A2 => n24137, B1 => n24151, B2 => 
                           n23736, ZN => n26158);
   U621 : AOI211_X1 port map( C1 => n24155, C2 => n23600, A => n23745, B => 
                           n23744, ZN => n26537);
   U622 : OAI22_X1 port map( A1 => n26536, A2 => n24158, B1 => n26537, B2 => 
                           n24156, ZN => n26157);
   U623 : AOI211_X1 port map( C1 => n24153, C2 => n23760, A => n26158, B => 
                           n26157, ZN => n26542);
   U624 : OAI222_X1 port map( A1 => n24168, A2 => n26542, B1 => n24081, B2 => 
                           n26159, C1 => n23979, C2 => n26543, ZN => n26612);
   U625 : INV_X1 port map( A => n26612, ZN => n26603);
   U626 : AOI22_X1 port map( A1 => n23963, A2 => n26923, B1 => n23630, B2 => 
                           n26611, ZN => n26161);
   U627 : AOI22_X1 port map( A1 => n24061, A2 => n26604, B1 => n27679, B2 => 
                           n26910, ZN => n26160);
   U628 : OAI211_X1 port map( C1 => n26603, C2 => n27661, A => n26161, B => 
                           n26160, ZN => n26813);
   U629 : AOI22_X1 port map( A1 => n24093, A2 => n26841, B1 => n23962, B2 => 
                           n26813, ZN => n26162);
   U630 : OAI22_X1 port map( A1 => n24029, A2 => n26162, B1 => n24030, B2 => 
                           n23636, ZN => n26163);
   U631 : OR4_X1 port map( A1 => n24166, A2 => n23886, A3 => n25880, A4 => 
                           n26163, ZN => OUTALU(21));
   U632 : NAND2_X1 port map( A1 => n14287, A2 => n19292, ZN => n26164);
   U633 : OR2_X1 port map( A1 => n19293, A2 => n26164, ZN => n22800);
   U634 : INV_X1 port map( A => n19293, ZN => n1808);
   U635 : OAI21_X1 port map( B1 => n14287, B2 => n19292, A => n26164, ZN => 
                           n22765);
   U636 : NOR2_X1 port map( A1 => n1808, A2 => n22765, ZN => n22797);
   U637 : INV_X1 port map( A => n27590, ZN => n27581);
   U638 : OAI21_X1 port map( B1 => DATA2(2), B2 => n27593, A => n27581, ZN => 
                           n1869);
   U639 : NAND2_X1 port map( A1 => n1830, A2 => n1869, ZN => n19271);
   U640 : INV_X1 port map( A => DATA2(4), ZN => n27577);
   U641 : NOR2_X1 port map( A1 => n27592, A2 => n27577, ZN => n27574);
   U642 : NOR2_X1 port map( A1 => n1865, A2 => n27574, ZN => n1866);
   U643 : INV_X1 port map( A => n1865, ZN => n26165);
   U644 : AOI21_X1 port map( B1 => n26166, B2 => n26165, A => n1866, ZN => 
                           n1864);
   U645 : INV_X1 port map( A => n1830, ZN => n26811);
   U646 : NOR2_X1 port map( A1 => n1864, A2 => n26811, ZN => n19261);
   U647 : OAI22_X1 port map( A1 => n26167, A2 => n27607, B1 => n26487, B2 => 
                           n27636, ZN => n26171);
   U648 : INV_X1 port map( A => n26168, ZN => n26489);
   U649 : OAI22_X1 port map( A1 => n27641, A2 => n26169, B1 => n26489, B2 => 
                           n27638, ZN => n26170);
   U650 : AOI211_X1 port map( C1 => n27645, C2 => n26493, A => n26171, B => 
                           n26170, ZN => n26975);
   U651 : INV_X1 port map( A => n1821, ZN => n26494);
   U652 : OAI22_X1 port map( A1 => n26975, A2 => n1856, B1 => n26494, B2 => 
                           n27564, ZN => n21296);
   U653 : NOR2_X1 port map( A1 => n1840, A2 => n26415, ZN => n26440);
   U654 : INV_X1 port map( A => DATA1(26), ZN => n27191);
   U655 : NAND2_X1 port map( A1 => DATA1(24), A2 => n26724, ZN => n26460);
   U656 : NAND2_X1 port map( A1 => DATA1(22), A2 => n26719, ZN => n26185);
   U657 : OAI211_X1 port map( C1 => n26750, C2 => n27191, A => n26460, B => 
                           n26185, ZN => n26172);
   U658 : AOI211_X1 port map( C1 => n26753, C2 => DATA1(25), A => n26440, B => 
                           n26172, ZN => n26178);
   U659 : NOR2_X1 port map( A1 => n26773, A2 => n26707, ZN => n26472);
   U660 : NAND2_X1 port map( A1 => DATA1(24), A2 => n26704, ZN => n26452);
   U661 : NAND2_X1 port map( A1 => DATA1(27), A2 => n26478, ZN => n26495);
   U662 : OAI211_X1 port map( C1 => n26666, C2 => n1840, A => n26452, B => 
                           n26495, ZN => n26173);
   U663 : AOI211_X1 port map( C1 => n26753, C2 => DATA1(26), A => n26472, B => 
                           n26173, ZN => n26182);
   U664 : NOR2_X1 port map( A1 => n27191, A2 => n26707, ZN => n26467);
   U665 : NAND2_X1 port map( A1 => DATA1(27), A2 => n26753, ZN => n26497);
   U666 : NAND2_X1 port map( A1 => DATA1(24), A2 => n26847, ZN => n26444);
   U667 : OAI211_X1 port map( C1 => n26750, C2 => n27198, A => n26497, B => 
                           n26444, ZN => n26174);
   U668 : AOI211_X1 port map( C1 => n26704, C2 => DATA1(25), A => n26467, B => 
                           n26174, ZN => n26793);
   U669 : OAI222_X1 port map( A1 => n26794, A2 => n26178, B1 => n26792, B2 => 
                           n26182, C1 => n26446, C2 => n26793, ZN => n27620);
   U670 : NOR2_X1 port map( A1 => n1840, A2 => n26722, ZN => n26463);
   U671 : NOR2_X1 port map( A1 => n27177, A2 => n26707, ZN => n26441);
   U672 : AOI211_X1 port map( C1 => DATA1(24), C2 => n26478, A => n26463, B => 
                           n26441, ZN => n26175);
   U673 : NAND2_X1 port map( A1 => DATA1(20), A2 => n26847, ZN => n26194);
   U674 : OAI211_X1 port map( C1 => n26415, C2 => n27653, A => n26175, B => 
                           n26194, ZN => n26210);
   U675 : INV_X1 port map( A => DATA1(24), ZN => n27185);
   U676 : NOR2_X1 port map( A1 => n1840, A2 => n26707, ZN => n26455);
   U677 : NOR2_X1 port map( A1 => n27653, A2 => n26666, ZN => n26191);
   U678 : AOI211_X1 port map( C1 => DATA1(25), C2 => n26478, A => n26455, B => 
                           n26191, ZN => n26176);
   U679 : NAND2_X1 port map( A1 => DATA1(22), A2 => n26704, ZN => n26214);
   U680 : OAI211_X1 port map( C1 => n26722, C2 => n27185, A => n26176, B => 
                           n26214, ZN => n26180);
   U681 : AOI22_X1 port map( A1 => n26207, A2 => n26210, B1 => n26205, B2 => 
                           n26180, ZN => n26177);
   U682 : OAI21_X1 port map( B1 => n26178, B2 => n26446, A => n26177, ZN => 
                           n27563);
   U683 : INV_X1 port map( A => n27563, ZN => n27623);
   U684 : OAI22_X1 port map( A1 => n26182, A2 => n26446, B1 => n26178, B2 => 
                           n26754, ZN => n26179);
   U685 : AOI21_X1 port map( B1 => n26207, B2 => n26180, A => n26179, ZN => 
                           n27616);
   U686 : OAI22_X1 port map( A1 => n27623, A2 => n27607, B1 => n27616, B2 => 
                           n27636, ZN => n26184);
   U687 : AOI222_X1 port map( A1 => n26180, A2 => n26209, B1 => n26206, B2 => 
                           n26207, C1 => n26210, C2 => n26205, ZN => n27559);
   U688 : INV_X1 port map( A => DATA1(27), ZN => n26737);
   U689 : NOR2_X1 port map( A1 => n26737, A2 => n26707, ZN => n26481);
   U690 : NAND2_X1 port map( A1 => DATA1(26), A2 => n26704, ZN => n26468);
   U691 : NAND2_X1 port map( A1 => DATA1(25), A2 => n26847, ZN => n26453);
   U692 : OAI211_X1 port map( C1 => n26750, C2 => n26703, A => n26468, B => 
                           n26453, ZN => n26181);
   U693 : AOI211_X1 port map( C1 => n26753, C2 => DATA1(28), A => n26481, B => 
                           n26181, ZN => n26791);
   U694 : OAI222_X1 port map( A1 => n26794, A2 => n26182, B1 => n26792, B2 => 
                           n26793, C1 => n26446, C2 => n26791, ZN => n27619);
   U695 : INV_X1 port map( A => n27619, ZN => n26820);
   U696 : OAI22_X1 port map( A1 => n27641, A2 => n27559, B1 => n26820, B2 => 
                           n26425, ZN => n26183);
   U697 : AOI211_X1 port map( C1 => n27709, C2 => n27620, A => n26184, B => 
                           n26183, ZN => n1816);
   U698 : AOI22_X1 port map( A1 => DATA1(21), A2 => n26704, B1 => DATA1(20), B2
                           => n26724, ZN => n26188);
   U699 : NAND2_X1 port map( A1 => DATA1(18), A2 => n26478, ZN => n26187);
   U700 : AND4_X1 port map( A1 => n26188, A2 => n26187, A3 => n26186, A4 => 
                           n26185, ZN => n26447);
   U701 : NOR2_X1 port map( A1 => n26461, A2 => n26915, ZN => n26193);
   U702 : OAI21_X1 port map( B1 => n26722, B2 => n26903, A => n26189, ZN => 
                           n26190);
   U703 : NOR4_X1 port map( A1 => n26193, A2 => n26192, A3 => n26191, A4 => 
                           n26190, ZN => n26218);
   U704 : NOR2_X1 port map( A1 => n26461, A2 => n26930, ZN => n26196);
   U705 : OAI21_X1 port map( B1 => n26707, B2 => n26903, A => n26194, ZN => 
                           n26195);
   U706 : NOR4_X1 port map( A1 => n26198, A2 => n26197, A3 => n26196, A4 => 
                           n26195, ZN => n26204);
   U707 : OAI222_X1 port map( A1 => n26794, A2 => n26447, B1 => n26792, B2 => 
                           n26218, C1 => n26446, C2 => n26204, ZN => n27604);
   U708 : INV_X1 port map( A => n27604, ZN => n26201);
   U709 : AOI22_X1 port map( A1 => n26209, A2 => n26199, B1 => n26205, B2 => 
                           n26202, ZN => n26200);
   U710 : OAI21_X1 port map( B1 => n26204, B2 => n26794, A => n26200, ZN => 
                           n26448);
   U711 : INV_X1 port map( A => n26448, ZN => n26222);
   U712 : OAI22_X1 port map( A1 => n27641, A2 => n26201, B1 => n26222, B2 => 
                           n27636, ZN => n21379);
   U713 : INV_X1 port map( A => n26202, ZN => n26203);
   U714 : OAI222_X1 port map( A1 => n26794, A2 => n26218, B1 => n26792, B2 => 
                           n26204, C1 => n25967, C2 => n26203, ZN => n26457);
   U715 : INV_X1 port map( A => n26457, ZN => n26221);
   U716 : OAI22_X1 port map( A1 => n26425, A2 => n1848, B1 => n26221, B2 => 
                           n25891, ZN => n21378);
   U717 : INV_X1 port map( A => n27559, ZN => n26211);
   U718 : AOI222_X1 port map( A1 => n26210, A2 => n26209, B1 => n26208, B2 => 
                           n26207, C1 => n26206, C2 => n26205, ZN => n27560);
   U719 : INV_X1 port map( A => n27560, ZN => n27599);
   U720 : AOI22_X1 port map( A1 => n25892, A2 => n26211, B1 => n27624, B2 => 
                           n27599, ZN => n26213);
   U721 : AOI22_X1 port map( A1 => n27632, A2 => n27563, B1 => n27645, B2 => 
                           n27620, ZN => n26212);
   U722 : OAI211_X1 port map( C1 => n27616, C2 => n27638, A => n26213, B => 
                           n26212, ZN => n19399);
   U723 : AOI22_X1 port map( A1 => DATA1(21), A2 => n26724, B1 => DATA1(23), B2
                           => n26847, ZN => n26217);
   U724 : AND4_X1 port map( A1 => n26217, A2 => n26216, A3 => n26215, A4 => 
                           n26214, ZN => n26456);
   U725 : OAI222_X1 port map( A1 => n26794, A2 => n26456, B1 => n26792, B2 => 
                           n26447, C1 => n25967, C2 => n26218, ZN => n27611);
   U726 : AOI22_X1 port map( A1 => n27709, A2 => n26448, B1 => n27624, B2 => 
                           n27611, ZN => n26220);
   U727 : AOI22_X1 port map( A1 => n25892, A2 => n27604, B1 => n1857, B2 => 
                           n26457, ZN => n26219);
   U728 : OAI211_X1 port map( C1 => n26425, C2 => n1846, A => n26220, B => 
                           n26219, ZN => n1826);
   U729 : OAI22_X1 port map( A1 => n27641, A2 => n26222, B1 => n1846, B2 => 
                           n27607, ZN => n21485);
   U730 : OAI22_X1 port map( A1 => n26425, A2 => n26237, B1 => n26238, B2 => 
                           n27638, ZN => n21484);
   U731 : OAI22_X1 port map( A1 => n27641, A2 => n26221, B1 => n1846, B2 => 
                           n27636, ZN => n21491);
   U732 : OAI22_X1 port map( A1 => n26425, A2 => n26238, B1 => n26222, B2 => 
                           n27607, ZN => n21490);
   U733 : OAI211_X1 port map( C1 => n26750, C2 => n24052, A => n26224, B => 
                           n26223, ZN => n26225);
   U734 : AOI211_X1 port map( C1 => n26753, C2 => n24049, A => n26226, B => 
                           n26225, ZN => n26352);
   U735 : OAI211_X1 port map( C1 => n24053, C2 => n26461, A => n26228, B => 
                           n26227, ZN => n26229);
   U736 : AOI211_X1 port map( C1 => n26753, C2 => n24175, A => n26230, B => 
                           n26229, ZN => n26392);
   U737 : OAI222_X1 port map( A1 => n26794, A2 => n26231, B1 => n26792, B2 => 
                           n26352, C1 => n26446, C2 => n26392, ZN => n27536);
   U738 : INV_X1 port map( A => n27536, ZN => n26233);
   U739 : OAI222_X1 port map( A1 => n26794, A2 => n26232, B1 => n26792, B2 => 
                           n26231, C1 => n26446, C2 => n26352, ZN => n26332);
   U740 : INV_X1 port map( A => n26332, ZN => n26490);
   U741 : OAI22_X1 port map( A1 => n26233, A2 => n26425, B1 => n26490, B2 => 
                           n27638, ZN => n26235);
   U742 : INV_X1 port map( A => n26309, ZN => n26488);
   U743 : OAI22_X1 port map( A1 => n27641, A2 => n26489, B1 => n26488, B2 => 
                           n27636, ZN => n26234);
   U744 : AOI211_X1 port map( C1 => n25892, C2 => n26493, A => n26235, B => 
                           n26234, ZN => n12526);
   U745 : OAI22_X1 port map( A1 => n27641, A2 => n1848, B1 => n26236, B2 => 
                           n27638, ZN => n26240);
   U746 : OAI22_X1 port map( A1 => n26238, A2 => n27607, B1 => n26237, B2 => 
                           n27636, ZN => n26239);
   U747 : AOI211_X1 port map( C1 => n27645, C2 => n26241, A => n26240, B => 
                           n26239, ZN => n13963);
   U748 : OAI22_X1 port map( A1 => n26975, A2 => n1836, B1 => n1828, B2 => 
                           n27564, ZN => n19001);
   U749 : OAI22_X1 port map( A1 => n26975, A2 => n1859, B1 => n26485, B2 => 
                           n1856, ZN => n19000);
   U750 : OAI22_X1 port map( A1 => n26975, A2 => n1896, B1 => n26485, B2 => 
                           n27564, ZN => n18999);
   U751 : INV_X1 port map( A => n4302, ZN => n27380);
   U752 : INV_X1 port map( A => n1811, ZN => n27588);
   U753 : NOR2_X1 port map( A1 => n27380, A2 => n27588, ZN => n19280);
   U754 : INV_X1 port map( A => n1813, ZN => n27585);
   U755 : NOR2_X1 port map( A1 => n7769, A2 => n27585, ZN => n21556);
   U756 : INV_X1 port map( A => n1812, ZN => n26242);
   U757 : NOR2_X1 port map( A1 => n26242, A2 => n21556, ZN => n19278);
   U758 : NOR2_X1 port map( A1 => n26932, A2 => n26916, ZN => n19277);
   U759 : AOI22_X1 port map( A1 => n1857, A2 => n26248, B1 => n27709, B2 => 
                           n27600, ZN => n26245);
   U760 : INV_X1 port map( A => n27597, ZN => n26243);
   U761 : AOI22_X1 port map( A1 => n26795, A2 => n27625, B1 => n27645, B2 => 
                           n26243, ZN => n26244);
   U762 : OAI211_X1 port map( C1 => n26251, C2 => n27607, A => n26245, B => 
                           n26244, ZN => n26278);
   U763 : INV_X1 port map( A => n1842, ZN => n26262);
   U764 : AOI22_X1 port map( A1 => n1843, A2 => n26278, B1 => n1861, B2 => 
                           n26262, ZN => n18993);
   U765 : INV_X1 port map( A => n1845, ZN => n26246);
   U766 : AOI22_X1 port map( A1 => n1858, A2 => n26246, B1 => n1894, B2 => 
                           n26278, ZN => n18989);
   U767 : INV_X1 port map( A => n26247, ZN => n27630);
   U768 : AOI22_X1 port map( A1 => n26795, A2 => n27630, B1 => n27645, B2 => 
                           n27600, ZN => n26250);
   U769 : AOI22_X1 port map( A1 => n25892, A2 => n27625, B1 => n27709, B2 => 
                           n26248, ZN => n26249);
   U770 : OAI211_X1 port map( C1 => n26251, C2 => n27636, A => n26250, B => 
                           n26249, ZN => n14004);
   U771 : AOI22_X1 port map( A1 => n1860, A2 => n26262, B1 => n1861, B2 => 
                           n14004, ZN => n18988);
   U772 : INV_X1 port map( A => DATA2(22), ZN => n27259);
   U773 : NOR3_X1 port map( A1 => n27549, A2 => n27259, A3 => n27177, ZN => 
                           n19202);
   U774 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n27587, ZN => n2808);
   U775 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n2808, ZN => n19200);
   U776 : NOR3_X1 port map( A1 => n24170, A2 => n23889, A3 => n1807, ZN => 
                           n3026);
   U777 : AOI221_X1 port map( B1 => n23889, B2 => n24170, C1 => n1807, C2 => 
                           n24170, A => n3026, ZN => n18872);
   U778 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, ZN => 
                           n26252);
   U779 : NOR3_X1 port map( A1 => n23969, A2 => n1807, A3 => n26252, ZN => 
                           n3030);
   U780 : AOI221_X1 port map( B1 => n23969, B2 => n26252, C1 => n1807, C2 => 
                           n26252, A => n3030, ZN => n18867);
   U781 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_4_8_port, ZN => 
                           n26253);
   U782 : NOR3_X1 port map( A1 => n23952, A2 => n1807, A3 => n26253, ZN => 
                           n3029);
   U783 : AOI21_X1 port map( B1 => n24102, B2 => data1_mul_0_port, A => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, ZN => n26254
                           );
   U784 : NOR2_X1 port map( A1 => n3029, A2 => n26254, ZN => n19272);
   U785 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_5_10_port, ZN => 
                           n26255);
   U786 : NOR3_X1 port map( A1 => n23968, A2 => n1807, A3 => n26255, ZN => 
                           n3028);
   U787 : AOI221_X1 port map( B1 => n23968, B2 => n26255, C1 => n1807, C2 => 
                           n26255, A => n3028, ZN => n19194);
   U788 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_6_12_port, ZN => 
                           n26256);
   U789 : NOR3_X1 port map( A1 => n23948, A2 => n1807, A3 => n26256, ZN => 
                           n3027);
   U790 : AOI221_X1 port map( B1 => n23948, B2 => n26256, C1 => n1807, C2 => 
                           n26256, A => n3027, ZN => n18861);
   U791 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n27524);
   U792 : INV_X1 port map( A => n27524, ZN => n27528);
   U793 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN 
                           => n27279);
   U794 : NAND2_X1 port map( A1 => n27279, A2 => data2_mul_1_port, ZN => n27522
                           );
   U795 : INV_X1 port map( A => n27522, ZN => n27526);
   U796 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => n27279, ZN => n27511)
                           ;
   U797 : AOI222_X1 port map( A1 => n27528, A2 => n25898, B1 => n27526, B2 => 
                           n25900, C1 => n27511, C2 => n9081, ZN => n26258);
   U798 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n27318);
   U799 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n27318, ZN => n27280);
   U800 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n27280, ZN => n26257
                           );
   U801 : NOR2_X1 port map( A1 => n26258, A2 => n26257, ZN => n3036);
   U802 : AOI21_X1 port map( B1 => n26258, B2 => n26257, A => n3036, ZN => 
                           n19187);
   U803 : OAI22_X1 port map( A1 => n26488, A2 => n27607, B1 => n26490, B2 => 
                           n27636, ZN => n26261);
   U804 : AOI22_X1 port map( A1 => n27536, A2 => n27709, B1 => n26795, B2 => 
                           n26493, ZN => n26259);
   U805 : INV_X1 port map( A => n26259, ZN => n26260);
   U806 : OAI21_X1 port map( B1 => n26261, B2 => n26260, A => n1831, ZN => 
                           n19186);
   U807 : INV_X1 port map( A => n1844, ZN => n26263);
   U808 : AOI22_X1 port map( A1 => n1858, A2 => n26263, B1 => n1894, B2 => 
                           n26262, ZN => n18982);
   U809 : AOI22_X1 port map( A1 => n1843, A2 => n14004, B1 => n1861, B2 => 
                           n26278, ZN => n18981);
   U810 : NOR2_X1 port map( A1 => n26266, A2 => n26265, ZN => n26264);
   U811 : OR2_X1 port map( A1 => n27710, A2 => n26979, ZN => n27550);
   U812 : AOI211_X1 port map( C1 => n26266, C2 => n26265, A => n26264, B => 
                           n27550, ZN => n26273);
   U813 : INV_X1 port map( A => DATA2(9), ZN => n27271);
   U814 : NAND2_X1 port map( A1 => DATA1(9), A2 => n27271, ZN => n27093);
   U815 : INV_X1 port map( A => n27093, ZN => n27146);
   U816 : NOR2_X1 port map( A1 => DATA1(9), A2 => n27271, ZN => n27144);
   U817 : NOR2_X1 port map( A1 => n27146, A2 => n27144, ZN => n27067);
   U818 : AND2_X1 port map( A1 => n24181, A2 => DATA2_I_8_port, ZN => n26268);
   U819 : INV_X1 port map( A => n1789, ZN => n27021);
   U820 : OAI211_X1 port map( C1 => n26269, C2 => n26268, A => n27021, B => 
                           n26267, ZN => n26271);
   U821 : NAND3_X1 port map( A1 => DATA2(9), A2 => DATA1(9), A3 => n26981, ZN 
                           => n26270);
   U822 : OAI211_X1 port map( C1 => n27067, C2 => n27570, A => n26271, B => 
                           n26270, ZN => n26272);
   U823 : AOI211_X1 port map( C1 => n23846, C2 => n27542, A => n26273, B => 
                           n26272, ZN => n19185);
   U824 : OAI22_X1 port map( A1 => n27641, A2 => n27597, B1 => n27559, B2 => 
                           n27638, ZN => n26275);
   U825 : OAI22_X1 port map( A1 => n27596, A2 => n27607, B1 => n27560, B2 => 
                           n27636, ZN => n26274);
   U826 : AOI211_X1 port map( C1 => n27645, C2 => n27563, A => n26275, B => 
                           n26274, ZN => n1837);
   U827 : OAI22_X1 port map( A1 => n26425, A2 => n27559, B1 => n27596, B2 => 
                           n27636, ZN => n26277);
   U828 : OAI22_X1 port map( A1 => n27597, A2 => n27607, B1 => n27560, B2 => 
                           n27638, ZN => n26276);
   U829 : AOI211_X1 port map( C1 => n27624, C2 => n27600, A => n26277, B => 
                           n26276, ZN => n18992);
   U830 : OAI22_X1 port map( A1 => n18992, A2 => n1856, B1 => n1837, B2 => 
                           n1896, ZN => n21603);
   U831 : OAI22_X1 port map( A1 => n18992, A2 => n27564, B1 => n1837, B2 => 
                           n1856, ZN => n21604);
   U832 : INV_X1 port map( A => n26278, ZN => n26311);
   U833 : OAI22_X1 port map( A1 => n26311, A2 => n27564, B1 => n1837, B2 => 
                           n1836, ZN => n21607);
   U834 : OAI211_X1 port map( C1 => n24057, C2 => n23741, A => n23725, B => 
                           n23724, ZN => n26313);
   U835 : AOI22_X1 port map( A1 => n24149, A2 => n23732, B1 => n23955, B2 => 
                           n24148, ZN => n26279);
   U836 : OAI211_X1 port map( C1 => n23957, C2 => n23730, A => n23731, B => 
                           n26279, ZN => n26303);
   U837 : OAI22_X1 port map( A1 => n23954, A2 => n23741, B1 => n24151, B2 => 
                           n23730, ZN => n26280);
   U838 : AOI211_X1 port map( C1 => n24060, C2 => n23759, A => n23720, B => 
                           n26280, ZN => n26292);
   U839 : INV_X1 port map( A => n26292, ZN => n26291);
   U840 : AOI222_X1 port map( A1 => n27673, A2 => n26313, B1 => n26303, B2 => 
                           n27662, C1 => n26291, C2 => n27663, ZN => n26369);
   U841 : OAI22_X1 port map( A1 => n24151, A2 => n24145, B1 => n23957, B2 => 
                           n25877, ZN => n26281);
   U842 : AOI211_X1 port map( C1 => n24101, C2 => n27694, A => n23722, B => 
                           n26281, ZN => n26293);
   U843 : OAI22_X1 port map( A1 => n23953, A2 => n24146, B1 => n25877, B2 => 
                           n27691, ZN => n26282);
   U844 : AOI211_X1 port map( C1 => n25878, C2 => n27687, A => n23721, B => 
                           n26282, ZN => n26300);
   U845 : INV_X1 port map( A => n26300, ZN => n26284);
   U846 : OAI22_X1 port map( A1 => n23954, A2 => n23730, B1 => n24158, B2 => 
                           n23741, ZN => n26283);
   U847 : AOI211_X1 port map( C1 => n24107, C2 => n23629, A => n23628, B => 
                           n26283, ZN => n26294);
   U848 : INV_X1 port map( A => n26294, ZN => n26290);
   U849 : AOI22_X1 port map( A1 => n27663, A2 => n26284, B1 => n27673, B2 => 
                           n26290, ZN => n26285);
   U850 : OAI21_X1 port map( B1 => n23979, B2 => n26293, A => n26285, ZN => 
                           n26990);
   U851 : AOI22_X1 port map( A1 => n27690, A2 => n24058, B1 => n24153, B2 => 
                           n24126, ZN => n26286);
   U852 : INV_X1 port map( A => n26286, ZN => n26289);
   U853 : AOI22_X1 port map( A1 => n27699, A2 => n25878, B1 => n24060, B2 => 
                           n23753, ZN => n26287);
   U854 : INV_X1 port map( A => n26287, ZN => n26288);
   U855 : AOI211_X1 port map( C1 => n24101, C2 => n23629, A => n26289, B => 
                           n26288, ZN => n26935);
   U856 : OAI222_X1 port map( A1 => n24168, A2 => n26293, B1 => n24081, B2 => 
                           n26935, C1 => n23979, C2 => n26300, ZN => n26988);
   U857 : AOI22_X1 port map( A1 => n24104, A2 => n26990, B1 => n27677, B2 => 
                           n26988, ZN => n26296);
   U858 : AOI222_X1 port map( A1 => n27662, A2 => n26291, B1 => n27663, B2 => 
                           n26290, C1 => n27673, C2 => n26303, ZN => n26304);
   U859 : INV_X1 port map( A => n26304, ZN => n26348);
   U860 : OAI222_X1 port map( A1 => n23979, A2 => n26294, B1 => n24080, B2 => 
                           n26293, C1 => n24105, C2 => n26292, ZN => n26998);
   U861 : AOI22_X1 port map( A1 => n27666, A2 => n26348, B1 => n27683, B2 => 
                           n26998, ZN => n26295);
   U862 : OAI211_X1 port map( C1 => n24113, C2 => n26369, A => n26296, B => 
                           n26295, ZN => n27028);
   U863 : INV_X1 port map( A => n26988, ZN => n26999);
   U864 : INV_X1 port map( A => n26990, ZN => n27002);
   U865 : OAI22_X1 port map( A1 => n23891, A2 => n26999, B1 => n27002, B2 => 
                           n27672, ZN => n26302);
   U866 : NOR2_X1 port map( A1 => n24151, A2 => n23638, ZN => n26297);
   U867 : AOI21_X1 port map( B1 => n24149, B2 => n23753, A => n26297, ZN => 
                           n26299);
   U868 : AOI22_X1 port map( A1 => n24150, A2 => n25878, B1 => n24106, B2 => 
                           n23677, ZN => n26298);
   U869 : OAI211_X1 port map( C1 => n25877, C2 => n27689, A => n26299, B => 
                           n26298, ZN => n26927);
   U870 : INV_X1 port map( A => n26927, ZN => n26934);
   U871 : OAI222_X1 port map( A1 => n23979, A2 => n26935, B1 => n26300, B2 => 
                           n24168, C1 => n26934, C2 => n24081, ZN => n26989);
   U872 : INV_X1 port map( A => n26989, ZN => n27001);
   U873 : OAI22_X1 port map( A1 => n26304, A2 => n27661, B1 => n27001, B2 => 
                           n27664, ZN => n26301);
   U874 : AOI211_X1 port map( C1 => n24123, C2 => n26998, A => n26302, B => 
                           n26301, ZN => n26349);
   U875 : INV_X1 port map( A => n26349, ZN => n27029);
   U876 : OAI211_X1 port map( C1 => n24158, C2 => n24124, A => n23728, B => 
                           n23727, ZN => n26344);
   U877 : AOI222_X1 port map( A1 => n26313, A2 => n24097, B1 => n26303, B2 => 
                           n24038, C1 => n26344, C2 => n23967, ZN => n26374);
   U878 : OAI22_X1 port map( A1 => n23633, A2 => n26369, B1 => n24113, B2 => 
                           n26374, ZN => n26306);
   U879 : OAI22_X1 port map( A1 => n24108, A2 => n26304, B1 => n24090, B2 => 
                           n27002, ZN => n26305);
   U880 : AOI211_X1 port map( C1 => n24104, C2 => n26998, A => n26306, B => 
                           n26305, ZN => n26385);
   U881 : INV_X1 port map( A => n26385, ZN => n26307);
   U882 : AOI222_X1 port map( A1 => n27028, A2 => n24093, B1 => n27029, B2 => 
                           n23632, C1 => n26307, C2 => n23962, ZN => n26308);
   U883 : OAI211_X1 port map( C1 => n24036, C2 => n26308, A => n23935, B => 
                           n23723, ZN => OUTALU(9));
   U884 : CLKBUF_X1 port map( A => n22313, Z => n27567);
   U885 : NAND2_X1 port map( A1 => n24181, A2 => n27272, ZN => n27090);
   U886 : OAI21_X1 port map( B1 => n24181, B2 => n27272, A => n27090, ZN => 
                           n27043);
   U887 : AOI22_X1 port map( A1 => n24020, A2 => n27567, B1 => n27557, B2 => 
                           n27043, ZN => n18980);
   U888 : NOR3_X1 port map( A1 => n24046, A2 => n27549, A3 => n27272, ZN => 
                           n21634);
   U889 : AOI222_X1 port map( A1 => n26309, A2 => n27624, B1 => n27536, B2 => 
                           n1857, C1 => n26332, C2 => n25892, ZN => n26310);
   U890 : INV_X1 port map( A => n1831, ZN => n26391);
   U891 : OAI22_X1 port map( A1 => n21635, A2 => n27550, B1 => n26310, B2 => 
                           n26391, ZN => n21633);
   U892 : OAI22_X1 port map( A1 => n26311, A2 => n1836, B1 => n1844, B2 => 
                           n1896, ZN => n18977);
   U893 : AOI22_X1 port map( A1 => n23632, A2 => n27028, B1 => n24095, B2 => 
                           n27029, ZN => n26320);
   U894 : OAI22_X1 port map( A1 => n24156, A2 => n23726, B1 => n24158, B2 => 
                           n24144, ZN => n26312);
   U895 : AOI211_X1 port map( C1 => n23732, C2 => n24107, A => n23717, B => 
                           n26312, ZN => n26368);
   U896 : INV_X1 port map( A => n26368, ZN => n26345);
   U897 : AOI22_X1 port map( A1 => n27662, A2 => n26344, B1 => n27663, B2 => 
                           n26313, ZN => n26314);
   U898 : INV_X1 port map( A => n26314, ZN => n26315);
   U899 : AOI21_X1 port map( B1 => n27673, B2 => n26345, A => n26315, ZN => 
                           n26399);
   U900 : OAI22_X1 port map( A1 => n23633, A2 => n26374, B1 => n24113, B2 => 
                           n26399, ZN => n26316);
   U901 : INV_X1 port map( A => n26316, ZN => n26318);
   U902 : AOI22_X1 port map( A1 => n23963, A2 => n26998, B1 => n27679, B2 => 
                           n26348, ZN => n26317);
   U903 : OAI211_X1 port map( C1 => n24062, C2 => n26369, A => n26318, B => 
                           n26317, ZN => n26408);
   U904 : NAND2_X1 port map( A1 => n23962, A2 => n26408, ZN => n26319);
   U905 : OAI211_X1 port map( C1 => n23635, C2 => n26385, A => n26320, B => 
                           n26319, ZN => n26321);
   U906 : AOI22_X1 port map( A1 => n23960, A2 => n24019, B1 => n27703, B2 => 
                           n26321, ZN => n26323);
   U907 : NOR2_X1 port map( A1 => n23934, A2 => n23718, ZN => n26322);
   U908 : NAND3_X1 port map( A1 => n23719, A2 => n26323, A3 => n26322, ZN => 
                           OUTALU(8));
   U909 : INV_X1 port map( A => n27033, ZN => n27652);
   U910 : INV_X1 port map( A => n27018, ZN => n27651);
   U911 : AOI21_X1 port map( B1 => n27652, B2 => n27704, A => n27651, ZN => 
                           n26324);
   U912 : OAI21_X1 port map( B1 => n24179, B2 => n27570, A => n26324, ZN => 
                           n26331);
   U913 : INV_X1 port map( A => n26424, ZN => n27036);
   U914 : OAI22_X1 port map( A1 => n26326, A2 => n27036, B1 => n1825, B2 => 
                           n26325, ZN => n26327);
   U915 : INV_X1 port map( A => n26327, ZN => n27538);
   U916 : NOR2_X1 port map( A1 => n26424, A2 => n27040, ZN => n26334);
   U917 : INV_X1 port map( A => n26328, ZN => n26337);
   U918 : AOI211_X1 port map( C1 => n27538, C2 => n26329, A => n26334, B => 
                           n26337, ZN => n26330);
   U919 : AOI22_X1 port map( A1 => DATA2(7), A2 => n26331, B1 => n26330, B2 => 
                           n26333, ZN => n18976);
   U920 : AOI22_X1 port map( A1 => n25892, A2 => n27536, B1 => n27624, B2 => 
                           n26332, ZN => n26339);
   U921 : NOR2_X1 port map( A1 => n24047, A2 => DATA2(7), ZN => n27139);
   U922 : OAI22_X1 port map( A1 => n27539, A2 => n26335, B1 => n26334, B2 => 
                           n26333, ZN => n26336);
   U923 : AOI22_X1 port map( A1 => n27139, A2 => n27557, B1 => n26337, B2 => 
                           n26336, ZN => n26338);
   U924 : OAI21_X1 port map( B1 => n26339, B2 => n26391, A => n26338, ZN => 
                           n26340);
   U925 : AOI21_X1 port map( B1 => n22313, B2 => n23854, A => n26340, ZN => 
                           n19184);
   U926 : OAI22_X1 port map( A1 => n23633, A2 => n26399, B1 => n24108, B2 => 
                           n26374, ZN => n26347);
   U927 : AOI22_X1 port map( A1 => n27669, A2 => n27697, B1 => n23732, B2 => 
                           n24153, ZN => n26343);
   U928 : OAI22_X1 port map( A1 => n24151, A2 => n24143, B1 => n24158, B2 => 
                           n23726, ZN => n26341);
   U929 : INV_X1 port map( A => n26341, ZN => n26342);
   U930 : OAI211_X1 port map( C1 => n23954, C2 => n24144, A => n26343, B => 
                           n26342, ZN => n26364);
   U931 : AOI222_X1 port map( A1 => n27662, A2 => n26345, B1 => n27663, B2 => 
                           n26344, C1 => n26364, C2 => n27673, ZN => n26427);
   U932 : OAI22_X1 port map( A1 => n23891, A2 => n26369, B1 => n26427, B2 => 
                           n24072, ZN => n26346);
   U933 : AOI211_X1 port map( C1 => n23964, C2 => n26348, A => n26347, B => 
                           n26346, ZN => n26407);
   U934 : INV_X1 port map( A => n26408, ZN => n26384);
   U935 : OAI22_X1 port map( A1 => n24112, A2 => n26407, B1 => n23635, B2 => 
                           n26384, ZN => n26351);
   U936 : OAI22_X1 port map( A1 => n24122, A2 => n26385, B1 => n26349, B2 => 
                           n27681, ZN => n26350);
   U937 : AOI211_X1 port map( C1 => n27675, C2 => n27028, A => n26351, B => 
                           n26350, ZN => n27544);
   U938 : OAI211_X1 port map( C1 => n27544, C2 => n24035, A => n23933, B => 
                           n23932, ZN => OUTALU(7));
   U939 : OAI21_X1 port map( B1 => n24056, B2 => n27033, A => n27018, ZN => 
                           n26354);
   U940 : OAI22_X1 port map( A1 => n26352, A2 => n26769, B1 => n26392, B2 => 
                           n26754, ZN => n26353);
   U941 : AOI22_X1 port map( A1 => DATA2(5), A2 => n26354, B1 => n1831, B2 => 
                           n26353, ZN => n18974);
   U942 : NOR2_X1 port map( A1 => n24056, A2 => DATA2(5), ZN => n27087);
   U943 : NOR2_X1 port map( A1 => n27276, A2 => n24177, ZN => n27085);
   U944 : NOR2_X1 port map( A1 => n27087, A2 => n27085, ZN => n27046);
   U945 : INV_X1 port map( A => n27046, ZN => n26355);
   U946 : AOI22_X1 port map( A1 => n27567, A2 => n23861, B1 => n27557, B2 => 
                           n26355, ZN => n18973);
   U947 : OAI22_X1 port map( A1 => n26357, A2 => n27036, B1 => n26356, B2 => 
                           n1825, ZN => n26362);
   U948 : INV_X1 port map( A => n26357, ZN => n26359);
   U949 : OAI22_X1 port map( A1 => n26359, A2 => n27036, B1 => n1825, B2 => 
                           n26358, ZN => n26361);
   U950 : AOI22_X1 port map( A1 => n26363, A2 => n26362, B1 => n26361, B2 => 
                           n26360, ZN => n18972);
   U951 : OAI22_X1 port map( A1 => n24122, A2 => n26384, B1 => n26407, B2 => 
                           n27686, ZN => n26373);
   U952 : INV_X1 port map( A => n26364, ZN => n26378);
   U953 : NOR2_X1 port map( A1 => n24151, A2 => n24144, ZN => n26366);
   U954 : OAI22_X1 port map( A1 => n23954, A2 => n23726, B1 => n24158, B2 => 
                           n23749, ZN => n26365);
   U955 : AOI211_X1 port map( C1 => n23755, C2 => n24101, A => n26366, B => 
                           n26365, ZN => n26367);
   U956 : OAI21_X1 port map( B1 => n23957, B2 => n24143, A => n26367, ZN => 
                           n26380);
   U957 : INV_X1 port map( A => n26380, ZN => n26404);
   U958 : OAI222_X1 port map( A1 => n23979, A2 => n26378, B1 => n24080, B2 => 
                           n26368, C1 => n26404, C2 => n24105, ZN => n26688);
   U959 : OAI22_X1 port map( A1 => n24108, A2 => n26399, B1 => n23891, B2 => 
                           n26374, ZN => n26371);
   U960 : OAI22_X1 port map( A1 => n23633, A2 => n26427, B1 => n24090, B2 => 
                           n26369, ZN => n26370);
   U961 : AOI211_X1 port map( C1 => n23887, C2 => n26688, A => n26371, B => 
                           n26370, ZN => n26409);
   U962 : OAI22_X1 port map( A1 => n24112, A2 => n26409, B1 => n23895, B2 => 
                           n26385, ZN => n26372);
   U963 : AOI211_X1 port map( C1 => n27665, C2 => n27028, A => n26373, B => 
                           n26372, ZN => n27543);
   U964 : OAI22_X1 port map( A1 => n26399, A2 => n27678, B1 => n26374, B2 => 
                           n24090, ZN => n26382);
   U965 : AOI22_X1 port map( A1 => n24149, A2 => n24142, B1 => n23955, B2 => 
                           n24131, ZN => n26376);
   U966 : NAND2_X1 port map( A1 => n24150, A2 => n24141, ZN => n26375);
   U967 : OAI211_X1 port map( C1 => n24158, C2 => n24125, A => n26376, B => 
                           n26375, ZN => n26377);
   U968 : AOI21_X1 port map( B1 => n24152, B2 => n23729, A => n26377, ZN => 
                           n26430);
   U969 : OAI22_X1 port map( A1 => n26430, A2 => n24067, B1 => n24080, B2 => 
                           n26378, ZN => n26379);
   U970 : AOI21_X1 port map( B1 => n27662, B2 => n26380, A => n26379, ZN => 
                           n26686);
   U971 : OAI22_X1 port map( A1 => n26686, A2 => n27661, B1 => n26427, B2 => 
                           n27672, ZN => n26381);
   U972 : AOI211_X1 port map( C1 => n24123, C2 => n26688, A => n26382, B => 
                           n26381, ZN => n26383);
   U973 : INV_X1 port map( A => n26383, ZN => n26872);
   U974 : OAI22_X1 port map( A1 => n23895, A2 => n26384, B1 => n24063, B2 => 
                           n26407, ZN => n26387);
   U975 : OAI22_X1 port map( A1 => n24034, A2 => n26385, B1 => n23635, B2 => 
                           n26409, ZN => n26386);
   U976 : AOI211_X1 port map( C1 => n23962, C2 => n26872, A => n26387, B => 
                           n26386, ZN => n26436);
   U977 : OAI22_X1 port map( A1 => n24110, A2 => n27544, B1 => n23966, B2 => 
                           n26436, ZN => n26388);
   U978 : INV_X1 port map( A => n26388, ZN => n26389);
   U979 : OAI21_X1 port map( B1 => n24103, B2 => n27543, A => n26389, ZN => 
                           n26398);
   U980 : NAND3_X1 port map( A1 => n23888, A2 => n24085, A3 => n26398, ZN => 
                           n26390);
   U981 : NAND4_X1 port map( A1 => n23714, A2 => n23716, A3 => n23715, A4 => 
                           n26390, ZN => OUTALU(5));
   U982 : AOI22_X1 port map( A1 => n26397, A2 => n26424, B1 => n27040, B2 => 
                           n26396, ZN => n18969);
   U983 : NOR3_X1 port map( A1 => n26392, A2 => n26391, A3 => n26769, ZN => 
                           n26395);
   U984 : NAND2_X1 port map( A1 => DATA2(4), A2 => n24054, ZN => n27137);
   U985 : NAND2_X1 port map( A1 => n24176, A2 => n27577, ZN => n27131);
   U986 : AND2_X1 port map( A1 => n27137, A2 => n27131, ZN => n27065);
   U987 : AOI21_X1 port map( B1 => n24176, B2 => n27652, A => n27651, ZN => 
                           n26393);
   U988 : OAI22_X1 port map( A1 => n27065, A2 => n27570, B1 => n26393, B2 => 
                           n27577, ZN => n26394);
   U989 : AOI211_X1 port map( C1 => n27542, C2 => n23623, A => n26395, B => 
                           n26394, ZN => n18968);
   U990 : OAI22_X1 port map( A1 => n26397, A2 => n27036, B1 => n26396, B2 => 
                           n1825, ZN => n18967);
   U991 : INV_X1 port map( A => n26398, ZN => n26861);
   U992 : OAI22_X1 port map( A1 => n27664, A2 => n26399, B1 => n27678, B2 => 
                           n26427, ZN => n26400);
   U993 : INV_X1 port map( A => n26400, ZN => n26406);
   U994 : AOI22_X1 port map( A1 => n24149, A2 => n23710, B1 => n23955, B2 => 
                           n24141, ZN => n26402);
   U995 : NAND2_X1 port map( A1 => n24153, A2 => n24131, ZN => n26401);
   U996 : OAI211_X1 port map( C1 => n23954, C2 => n24125, A => n26402, B => 
                           n26401, ZN => n26403);
   U997 : AOI21_X1 port map( B1 => n24142, B2 => n24040, A => n26403, ZN => 
                           n26685);
   U998 : OAI222_X1 port map( A1 => n23979, A2 => n26430, B1 => n24067, B2 => 
                           n26685, C1 => n24080, C2 => n26404, ZN => n27227);
   U999 : AOI22_X1 port map( A1 => n23887, A2 => n27227, B1 => n23630, B2 => 
                           n26688, ZN => n26405);
   U1000 : OAI211_X1 port map( C1 => n23633, C2 => n26686, A => n26406, B => 
                           n26405, ZN => n27215);
   U1001 : INV_X1 port map( A => n27215, ZN => n26435);
   U1002 : INV_X1 port map( A => n26407, ZN => n26426);
   U1003 : AOI22_X1 port map( A1 => n24082, A2 => n26408, B1 => n27675, B2 => 
                           n26426, ZN => n26411);
   U1004 : INV_X1 port map( A => n26409, ZN => n26691);
   U1005 : AOI22_X1 port map( A1 => n23632, A2 => n26691, B1 => n24092, B2 => 
                           n26872, ZN => n26410);
   U1006 : OAI211_X1 port map( C1 => n26435, C2 => n27674, A => n26411, B => 
                           n26410, ZN => n26695);
   U1007 : OAI22_X1 port map( A1 => n24103, A2 => n26436, B1 => n24110, B2 => 
                           n27543, ZN => n26412);
   U1008 : AOI21_X1 port map( B1 => n24065, B2 => n26695, A => n26412, ZN => 
                           n27212);
   U1009 : OAI22_X1 port map( A1 => n24091, A2 => n26861, B1 => n27212, B2 => 
                           n24111, ZN => n26413);
   U1010 : AOI22_X1 port map( A1 => n24085, A2 => n26413, B1 => n23711, B2 => 
                           n23961, ZN => n26414);
   U1011 : OAI211_X1 port map( C1 => n23961, C2 => n23713, A => n23712, B => 
                           n26414, ZN => OUTALU(4));
   U1012 : AOI22_X1 port map( A1 => n24175, A2 => n26724, B1 => n24048, B2 => 
                           n26847, ZN => n26417);
   U1013 : OR2_X1 port map( A1 => n26415, A2 => n24165, ZN => n26416);
   U1014 : OAI211_X1 port map( C1 => n24076, C2 => n26722, A => n26417, B => 
                           n26416, ZN => n26419);
   U1015 : NOR2_X1 port map( A1 => DATA2(3), A2 => n27682, ZN => n27082);
   U1016 : INV_X1 port map( A => n27082, ZN => n27132);
   U1017 : NAND2_X1 port map( A1 => DATA2(3), A2 => n24164, ZN => n27130);
   U1018 : AOI21_X1 port map( B1 => n27132, B2 => n27130, A => n27570, ZN => 
                           n26418);
   U1019 : AOI21_X1 port map( B1 => n1831, B2 => n26419, A => n26418, ZN => 
                           n18965);
   U1020 : OAI21_X1 port map( B1 => n24164, B2 => n27033, A => n27018, ZN => 
                           n26420);
   U1021 : AOI22_X1 port map( A1 => DATA2(3), A2 => n26420, B1 => n27567, B2 =>
                           n23880, ZN => n18964);
   U1022 : AOI21_X1 port map( B1 => n27532, B2 => n26422, A => n26421, ZN => 
                           n26423);
   U1023 : NAND2_X1 port map( A1 => n26424, A2 => n26423, ZN => n19269);
   U1024 : OAI22_X1 port map( A1 => n27641, A2 => n26853, B1 => n26857, B2 => 
                           n27636, ZN => n21746);
   U1025 : OAI22_X1 port map( A1 => n26425, A2 => n27635, B1 => n27640, B2 => 
                           n27638, ZN => n21745);
   U1026 : AOI22_X1 port map( A1 => n26872, A2 => n23631, B1 => n26426, B2 => 
                           n24082, ZN => n26434);
   U1027 : INV_X1 port map( A => n27227, ZN => n26868);
   U1028 : OAI22_X1 port map( A1 => n23633, A2 => n26868, B1 => n26427, B2 => 
                           n27664, ZN => n26432);
   U1029 : OAI22_X1 port map( A1 => n24151, A2 => n24139, B1 => n24158, B2 => 
                           n24140, ZN => n26429);
   U1030 : AOI211_X1 port map( C1 => n23931, C2 => n24171, A => n23707, B => 
                           n23706, ZN => n26862);
   U1031 : OAI22_X1 port map( A1 => n23954, A2 => n23752, B1 => n24156, B2 => 
                           n26862, ZN => n26428);
   U1032 : AOI211_X1 port map( C1 => n24153, C2 => n24115, A => n26429, B => 
                           n26428, ZN => n26864);
   U1033 : OAI222_X1 port map( A1 => n26864, A2 => n24105, B1 => n26430, B2 => 
                           n27696, C1 => n26685, C2 => n27671, ZN => n26687);
   U1034 : INV_X1 port map( A => n26687, ZN => n27231);
   U1035 : OAI22_X1 port map( A1 => n26686, A2 => n27672, B1 => n27231, B2 => 
                           n27661, ZN => n26431);
   U1036 : AOI211_X1 port map( C1 => n24104, C2 => n26688, A => n26432, B => 
                           n26431, ZN => n27236);
   U1037 : INV_X1 port map( A => n27236, ZN => n26873);
   U1038 : AOI22_X1 port map( A1 => n27684, A2 => n26691, B1 => n26873, B2 => 
                           n23962, ZN => n26433);
   U1039 : OAI211_X1 port map( C1 => n27686, C2 => n26435, A => n26434, B => 
                           n26433, ZN => n26876);
   U1040 : INV_X1 port map( A => n26436, ZN => n26437);
   U1041 : AOI222_X1 port map( A1 => n26876, A2 => n24084, B1 => n26695, B2 => 
                           n23975, C1 => n26437, C2 => n23970, ZN => n27213);
   U1042 : OAI222_X1 port map( A1 => n24091, A2 => n27212, B1 => n23977, B2 => 
                           n26861, C1 => n27213, C2 => n24111, ZN => n26438);
   U1043 : AOI22_X1 port map( A1 => n24085, A2 => n26438, B1 => n23980, B2 => 
                           n24032, ZN => n26439);
   U1044 : NAND4_X1 port map( A1 => n24018, A2 => n23709, A3 => n23708, A4 => 
                           n26439, ZN => OUTALU(3));
   U1045 : INV_X1 port map( A => n27611, ZN => n26451);
   U1046 : NOR2_X1 port map( A1 => n26461, A2 => n26833, ZN => n26443);
   U1047 : NOR4_X1 port map( A1 => n26443, A2 => n26442, A3 => n26441, A4 => 
                           n26440, ZN => n26445);
   U1048 : AND2_X1 port map( A1 => n26445, A2 => n26444, ZN => n26464);
   U1049 : OAI222_X1 port map( A1 => n26447, A2 => n26446, B1 => n26464, B2 => 
                           n26769, C1 => n26456, C2 => n26754, ZN => n27612);
   U1050 : AOI22_X1 port map( A1 => n27709, A2 => n26457, B1 => n27624, B2 => 
                           n27612, ZN => n26450);
   U1051 : AOI22_X1 port map( A1 => n27632, A2 => n27604, B1 => n27645, B2 => 
                           n26448, ZN => n26449);
   U1052 : OAI211_X1 port map( C1 => n26451, C2 => n27607, A => n26450, B => 
                           n26449, ZN => n11966);
   U1053 : INV_X1 port map( A => n27612, ZN => n26477);
   U1054 : OAI211_X1 port map( C1 => n26722, C2 => n27177, A => n26453, B => 
                           n26452, ZN => n26454);
   U1055 : AOI211_X1 port map( C1 => DATA1(21), C2 => n26478, A => n26455, B =>
                           n26454, ZN => n26473);
   U1056 : OAI222_X1 port map( A1 => n26794, A2 => n26473, B1 => n26792, B2 => 
                           n26464, C1 => n26446, C2 => n26456, ZN => n27609);
   U1057 : AOI22_X1 port map( A1 => n27632, A2 => n27611, B1 => n27624, B2 => 
                           n27609, ZN => n26459);
   U1058 : AOI22_X1 port map( A1 => n27709, A2 => n27604, B1 => n27645, B2 => 
                           n26457, ZN => n26458);
   U1059 : OAI211_X1 port map( C1 => n26477, C2 => n27607, A => n26459, B => 
                           n26458, ZN => n21841);
   U1060 : NAND2_X1 port map( A1 => DATA1(26), A2 => n26719, ZN => n26748);
   U1061 : OAI211_X1 port map( C1 => n26461, C2 => n27177, A => n26748, B => 
                           n26460, ZN => n26462);
   U1062 : AOI211_X1 port map( C1 => n26848, C2 => DATA1(25), A => n26463, B =>
                           n26462, ZN => n26474);
   U1063 : OAI222_X1 port map( A1 => n26794, A2 => n26474, B1 => n26792, B2 => 
                           n26473, C1 => n26446, C2 => n26464, ZN => n27610);
   U1064 : NAND2_X1 port map( A1 => DATA1(27), A2 => n26704, ZN => n26749);
   U1065 : NAND2_X1 port map( A1 => DATA1(24), A2 => n26478, ZN => n26465);
   U1066 : OAI211_X1 port map( C1 => n26722, C2 => n26773, A => n26749, B => 
                           n26465, ZN => n26466);
   U1067 : AOI211_X1 port map( C1 => n26847, C2 => DATA1(28), A => n26467, B =>
                           n26466, ZN => n26501);
   U1068 : NOR2_X1 port map( A1 => n27185, A2 => n26722, ZN => n26470);
   U1069 : NAND2_X1 port map( A1 => DATA1(27), A2 => n26719, ZN => n26730);
   U1070 : NAND2_X1 port map( A1 => n26730, A2 => n26468, ZN => n26469);
   U1071 : NOR4_X1 port map( A1 => n26472, A2 => n26471, A3 => n26470, A4 => 
                           n26469, ZN => n26482);
   U1072 : OAI222_X1 port map( A1 => n26769, A2 => n26501, B1 => n26792, B2 => 
                           n26482, C1 => n26446, C2 => n26474, ZN => n26509);
   U1073 : AOI22_X1 port map( A1 => n1857, A2 => n27610, B1 => n26795, B2 => 
                           n26509, ZN => n26476);
   U1074 : OAI222_X1 port map( A1 => n26769, A2 => n26482, B1 => n26754, B2 => 
                           n26474, C1 => n26446, C2 => n26473, ZN => n26507);
   U1075 : AOI22_X1 port map( A1 => n25892, A2 => n26507, B1 => n27709, B2 => 
                           n27609, ZN => n26475);
   U1076 : OAI211_X1 port map( C1 => n26425, C2 => n26477, A => n26476, B => 
                           n26475, ZN => n21843);
   U1077 : INV_X1 port map( A => n27609, ZN => n27608);
   U1078 : NAND2_X1 port map( A1 => DATA1(28), A2 => n26704, ZN => n26731);
   U1079 : NAND2_X1 port map( A1 => DATA1(25), A2 => n26478, ZN => n26479);
   U1080 : OAI211_X1 port map( C1 => n26722, C2 => n27191, A => n26731, B => 
                           n26479, ZN => n26480);
   U1081 : AOI211_X1 port map( C1 => n26847, C2 => DATA1(29), A => n26481, B =>
                           n26480, ZN => n26502);
   U1082 : OAI222_X1 port map( A1 => n26769, A2 => n26502, B1 => n26792, B2 => 
                           n26501, C1 => n26446, C2 => n26482, ZN => n26510);
   U1083 : AOI22_X1 port map( A1 => n1857, A2 => n26507, B1 => n26795, B2 => 
                           n26510, ZN => n26484);
   U1084 : AOI22_X1 port map( A1 => n25892, A2 => n26509, B1 => n27709, B2 => 
                           n27610, ZN => n26483);
   U1085 : OAI211_X1 port map( C1 => n26425, C2 => n27608, A => n26484, B => 
                           n26483, ZN => n26526);
   U1086 : AOI22_X1 port map( A1 => n1843, A2 => n21843, B1 => n1858, B2 => 
                           n26526, ZN => n18954);
   U1087 : OAI22_X1 port map( A1 => n1828, A2 => n1856, B1 => n26485, B2 => 
                           n1859, ZN => n18952);
   U1088 : OAI22_X1 port map( A1 => n1823, A2 => n1856, B1 => n26485, B2 => 
                           n1896, ZN => n18950);
   U1089 : INV_X1 port map( A => n1822, ZN => n26486);
   U1090 : OAI22_X1 port map( A1 => n1823, A2 => n27564, B1 => n26486, B2 => 
                           n1836, ZN => n18949);
   U1091 : OAI22_X1 port map( A1 => n26488, A2 => n27638, B1 => n27641, B2 => 
                           n26487, ZN => n26492);
   U1092 : OAI22_X1 port map( A1 => n26490, A2 => n26425, B1 => n26489, B2 => 
                           n27607, ZN => n26491);
   U1093 : AOI211_X1 port map( C1 => n1857, C2 => n26493, A => n26492, B => 
                           n26491, ZN => n1820);
   U1094 : OAI22_X1 port map( A1 => n26494, A2 => n1856, B1 => n1820, B2 => 
                           n1836, ZN => n18948);
   U1095 : NOR2_X1 port map( A1 => n26703, A2 => n26707, ZN => n26734);
   U1096 : NAND2_X1 port map( A1 => DATA1(31), A2 => n26719, ZN => n26518);
   U1097 : OAI211_X1 port map( C1 => n27198, C2 => n26722, A => n26518, B => 
                           n26495, ZN => n26496);
   U1098 : AOI211_X1 port map( C1 => DATA1(30), C2 => n26704, A => n26734, B =>
                           n26496, ZN => n26499);
   U1099 : NOR2_X1 port map( A1 => n27198, A2 => n26707, ZN => n26752);
   U1100 : NAND2_X1 port map( A1 => DATA1(29), A2 => n26704, ZN => n26720);
   U1101 : OAI211_X1 port map( C1 => n26750, C2 => n27191, A => n26497, B => 
                           n26720, ZN => n26498);
   U1102 : AOI211_X1 port map( C1 => n26847, C2 => DATA1(30), A => n26752, B =>
                           n26498, ZN => n26503);
   U1103 : OAI222_X1 port map( A1 => n26794, A2 => n26499, B1 => n26792, B2 => 
                           n26503, C1 => n25967, C2 => n26502, ZN => n26500);
   U1104 : AOI22_X1 port map( A1 => n27709, A2 => n26509, B1 => n27624, B2 => 
                           n26500, ZN => n26505);
   U1105 : OAI222_X1 port map( A1 => n26769, A2 => n26503, B1 => n26754, B2 => 
                           n26502, C1 => n25967, C2 => n26501, ZN => n26508);
   U1106 : AOI22_X1 port map( A1 => n25892, A2 => n26508, B1 => n27645, B2 => 
                           n26507, ZN => n26504);
   U1107 : NAND2_X1 port map( A1 => n26505, A2 => n26504, ZN => n26506);
   U1108 : AOI21_X1 port map( B1 => n27632, B2 => n26510, A => n26506, ZN => 
                           n19183);
   U1109 : INV_X1 port map( A => n26507, ZN => n27615);
   U1110 : AOI22_X1 port map( A1 => n27624, A2 => n26508, B1 => n27645, B2 => 
                           n27610, ZN => n26512);
   U1111 : AOI22_X1 port map( A1 => n25892, A2 => n26510, B1 => n1857, B2 => 
                           n26509, ZN => n26511);
   U1112 : OAI211_X1 port map( C1 => n27615, C2 => n27638, A => n26512, B => 
                           n26511, ZN => n21842);
   U1113 : AOI22_X1 port map( A1 => n1843, A2 => n21842, B1 => n1861, B2 => 
                           n26526, ZN => n18946);
   U1114 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n26712);
   U1115 : AOI21_X1 port map( B1 => n26712, B2 => n27659, A => n26713, ZN => 
                           n26515);
   U1116 : AOI21_X1 port map( B1 => n26712, B2 => n27657, A => n26713, ZN => 
                           n26514);
   U1117 : AOI22_X1 port map( A1 => n26786, A2 => n26515, B1 => n26788, B2 => 
                           n26514, ZN => n1787);
   U1118 : NAND2_X1 port map( A1 => DATA1(29), A2 => n4395, ZN => n26661);
   U1119 : INV_X1 port map( A => n26661, ZN => n26513);
   U1120 : AOI22_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, B1 => 
                           n26513, B2 => n1814, ZN => n26516);
   U1121 : OAI22_X1 port map( A1 => n26516, A2 => n27710, B1 => n1787, B2 => 
                           n26517, ZN => n26525);
   U1122 : XNOR2_X1 port map( A => DATA1(31), B => n4293, ZN => n26524);
   U1123 : INV_X1 port map( A => n26786, ZN => n27660);
   U1124 : OAI22_X1 port map( A1 => n26515, A2 => n27660, B1 => n26514, B2 => 
                           n27658, ZN => n26710);
   U1125 : OAI211_X1 port map( C1 => n26517, C2 => n26710, A => n27249, B => 
                           n26516, ZN => n26522);
   U1126 : INV_X1 port map( A => DATA2(31), ZN => n27250);
   U1127 : INV_X1 port map( A => DATA1(31), ZN => n26732);
   U1128 : AOI211_X1 port map( C1 => n27018, C2 => n27033, A => n27250, B => 
                           n26732, ZN => n26520);
   U1129 : NAND2_X1 port map( A1 => DATA1(31), A2 => n27250, ZN => n27210);
   U1130 : INV_X1 port map( A => n27210, ZN => n27204);
   U1131 : NAND2_X1 port map( A1 => DATA2(31), A2 => n26732, ZN => n27122);
   U1132 : INV_X1 port map( A => n27122, ZN => n27207);
   U1133 : NOR2_X1 port map( A1 => n27204, A2 => n27207, ZN => n27056);
   U1134 : OAI22_X1 port map( A1 => n27056, A2 => n27570, B1 => n26811, B2 => 
                           n26518, ZN => n26519);
   U1135 : AOI211_X1 port map( C1 => n23763, C2 => n27542, A => n26520, B => 
                           n26519, ZN => n26521);
   U1136 : OAI21_X1 port map( B1 => n26522, B2 => n26524, A => n26521, ZN => 
                           n26523);
   U1137 : AOI21_X1 port map( B1 => n26525, B2 => n26524, A => n26523, ZN => 
                           n18945);
   U1138 : AOI22_X1 port map( A1 => n1843, A2 => n26526, B1 => n1861, B2 => 
                           n21843, ZN => n21845);
   U1139 : NOR2_X1 port map( A1 => n23958, A2 => n24137, ZN => n26528);
   U1140 : AOI211_X1 port map( C1 => n23601, C2 => n24155, A => n23757, B => 
                           n23756, ZN => n26538);
   U1141 : OAI22_X1 port map( A1 => n26538, A2 => n24158, B1 => n26537, B2 => 
                           n23953, ZN => n26527);
   U1142 : AOI211_X1 port map( C1 => n24101, C2 => n23750, A => n26528, B => 
                           n26527, ZN => n26529);
   U1143 : OAI21_X1 port map( B1 => n26536, B2 => n24151, A => n26529, ZN => 
                           n26535);
   U1144 : AOI22_X1 port map( A1 => n23705, A2 => n24060, B1 => n27669, B2 => 
                           n27685, ZN => n26531);
   U1145 : INV_X1 port map( A => n26538, ZN => n26551);
   U1146 : AOI22_X1 port map( A1 => n23750, A2 => n27693, B1 => n26551, B2 => 
                           n27668, ZN => n26530);
   U1147 : OAI211_X1 port map( C1 => n23958, C2 => n26537, A => n26531, B => 
                           n26530, ZN => n26558);
   U1148 : AOI22_X1 port map( A1 => n24149, A2 => n23705, B1 => n23750, B2 => 
                           n24041, ZN => n26534);
   U1149 : OAI22_X1 port map( A1 => n23954, A2 => n26538, B1 => n24151, B2 => 
                           n26537, ZN => n26532);
   U1150 : INV_X1 port map( A => n26532, ZN => n26533);
   U1151 : OAI211_X1 port map( C1 => n26536, C2 => n23958, A => n26534, B => 
                           n26533, ZN => n26559);
   U1152 : AOI222_X1 port map( A1 => n27670, A2 => n26535, B1 => n26558, B2 => 
                           n27680, C1 => n27662, C2 => n26559, ZN => n26570);
   U1153 : INV_X1 port map( A => n26535, ZN => n26544);
   U1154 : INV_X1 port map( A => n26536, ZN => n26541);
   U1155 : OAI22_X1 port map( A1 => n24151, A2 => n24137, B1 => n23957, B2 => 
                           n23736, ZN => n26540);
   U1156 : OAI22_X1 port map( A1 => n26538, A2 => n24156, B1 => n26537, B2 => 
                           n24158, ZN => n26539);
   U1157 : AOI211_X1 port map( C1 => n24058, C2 => n26541, A => n26540, B => 
                           n26539, ZN => n26545);
   U1158 : OAI222_X1 port map( A1 => n24168, A2 => n26544, B1 => n24081, B2 => 
                           n26542, C1 => n26545, C2 => n23979, ZN => n26605);
   U1159 : AOI22_X1 port map( A1 => n23630, A2 => n26605, B1 => n27677, B2 => 
                           n26612, ZN => n26548);
   U1160 : OAI222_X1 port map( A1 => n24168, A2 => n26545, B1 => n24081, B2 => 
                           n26543, C1 => n23979, C2 => n26542, ZN => n26613);
   U1161 : INV_X1 port map( A => n26559, ZN => n26546);
   U1162 : OAI222_X1 port map( A1 => n24168, A2 => n26546, B1 => n24081, B2 => 
                           n26545, C1 => n23979, C2 => n26544, ZN => n26567);
   U1163 : AOI22_X1 port map( A1 => n24104, A2 => n26613, B1 => n24123, B2 => 
                           n26567, ZN => n26547);
   U1164 : OAI211_X1 port map( C1 => n26570, C2 => n27661, A => n26548, B => 
                           n26547, ZN => n26628);
   U1165 : INV_X1 port map( A => n26570, ZN => n26563);
   U1166 : AOI22_X1 port map( A1 => n23750, A2 => n24153, B1 => n27667, B2 => 
                           n27695, ZN => n26550);
   U1167 : AOI22_X1 port map( A1 => n24149, A2 => n24134, B1 => n23705, B2 => 
                           n23955, ZN => n26549);
   U1168 : OAI211_X1 port map( C1 => n25861, C2 => n27692, A => n26550, B => 
                           n26549, ZN => n26557);
   U1169 : AOI22_X1 port map( A1 => n23750, A2 => n23956, B1 => n24041, B2 => 
                           n27685, ZN => n26553);
   U1170 : AOI22_X1 port map( A1 => n24150, A2 => n23705, B1 => n24153, B2 => 
                           n26551, ZN => n26552);
   U1171 : OAI211_X1 port map( C1 => n24156, C2 => n23748, A => n26553, B => 
                           n26552, ZN => n26560);
   U1172 : AOI222_X1 port map( A1 => n26557, A2 => n24051, B1 => n26560, B2 => 
                           n24097, C1 => n26558, C2 => n24039, ZN => n26575);
   U1173 : AOI22_X1 port map( A1 => n24138, A2 => n24150, B1 => n27667, B2 => 
                           n27698, ZN => n26555);
   U1174 : AOI22_X1 port map( A1 => n24149, A2 => n23702, B1 => n23705, B2 => 
                           n24152, ZN => n26554);
   U1175 : OAI211_X1 port map( C1 => n25861, C2 => n27688, A => n26555, B => 
                           n26554, ZN => n26577);
   U1176 : AOI22_X1 port map( A1 => n24153, A2 => n23703, B1 => n23955, B2 => 
                           n24138, ZN => n26556);
   U1177 : OAI211_X1 port map( C1 => n23954, C2 => n23740, A => n23701, B => 
                           n26556, ZN => n26584);
   U1178 : AOI222_X1 port map( A1 => n26577, A2 => n24097, B1 => n26584, B2 => 
                           n24051, C1 => n26557, C2 => n24039, ZN => n26590);
   U1179 : OAI22_X1 port map( A1 => n26575, A2 => n27672, B1 => n24113, B2 => 
                           n26590, ZN => n26562);
   U1180 : AOI222_X1 port map( A1 => n26557, A2 => n24097, B1 => n26577, B2 => 
                           n24051, C1 => n26560, C2 => n24039, ZN => n26589);
   U1181 : AOI222_X1 port map( A1 => n26560, A2 => n24051, B1 => n26559, B2 => 
                           n24039, C1 => n26558, C2 => n24097, ZN => n26578);
   U1182 : OAI22_X1 port map( A1 => n23633, A2 => n26589, B1 => n26578, B2 => 
                           n23891, ZN => n26561);
   U1183 : AOI211_X1 port map( C1 => n26563, C2 => n27677, A => n26562, B => 
                           n26561, ZN => n26596);
   U1184 : OAI22_X1 port map( A1 => n23633, A2 => n26575, B1 => n24113, B2 => 
                           n26589, ZN => n26565);
   U1185 : OAI22_X1 port map( A1 => n26570, A2 => n23891, B1 => n26578, B2 => 
                           n24108, ZN => n26564);
   U1186 : AOI211_X1 port map( C1 => n23963, C2 => n26567, A => n26565, B => 
                           n26564, ZN => n26625);
   U1187 : OAI22_X1 port map( A1 => n24112, A2 => n26596, B1 => n26625, B2 => 
                           n23635, ZN => n26574);
   U1188 : INV_X1 port map( A => n26613, ZN => n26566);
   U1189 : OAI22_X1 port map( A1 => n24089, A2 => n26566, B1 => n24113, B2 => 
                           n26578, ZN => n26569);
   U1190 : INV_X1 port map( A => n26567, ZN => n26608);
   U1191 : OAI22_X1 port map( A1 => n24062, A2 => n26608, B1 => n23633, B2 => 
                           n26570, ZN => n26568);
   U1192 : AOI211_X1 port map( C1 => n24069, C2 => n26605, A => n26569, B => 
                           n26568, ZN => n26619);
   U1193 : OAI22_X1 port map( A1 => n23633, A2 => n26578, B1 => n24113, B2 => 
                           n26575, ZN => n26572);
   U1194 : OAI22_X1 port map( A1 => n26608, A2 => n23891, B1 => n26570, B2 => 
                           n24108, ZN => n26571);
   U1195 : AOI211_X1 port map( C1 => n23963, C2 => n26605, A => n26572, B => 
                           n26571, ZN => n26631);
   U1196 : OAI22_X1 port map( A1 => n26619, A2 => n23894, B1 => n26631, B2 => 
                           n24121, ZN => n26573);
   U1197 : AOI211_X1 port map( C1 => n24082, C2 => n26628, A => n26574, B => 
                           n26573, ZN => n26623);
   U1198 : INV_X1 port map( A => n26619, ZN => n26627);
   U1199 : INV_X1 port map( A => n26575, ZN => n26593);
   U1200 : AOI22_X1 port map( A1 => n24149, A2 => n23695, B1 => n23955, B2 => 
                           n24134, ZN => n26576);
   U1201 : OAI211_X1 port map( C1 => n23957, C2 => n23748, A => n23692, B => 
                           n26576, ZN => n26586);
   U1202 : AOI222_X1 port map( A1 => n26584, A2 => n24097, B1 => n26586, B2 => 
                           n24051, C1 => n26577, C2 => n24039, ZN => n26588);
   U1203 : OAI22_X1 port map( A1 => n23633, A2 => n26590, B1 => n24113, B2 => 
                           n26588, ZN => n26580);
   U1204 : OAI22_X1 port map( A1 => n24089, A2 => n26578, B1 => n24108, B2 => 
                           n26589, ZN => n26579);
   U1205 : AOI211_X1 port map( C1 => n24104, C2 => n26593, A => n26580, B => 
                           n26579, ZN => n26594);
   U1206 : OAI22_X1 port map( A1 => n24112, A2 => n26594, B1 => n24122, B2 => 
                           n26625, ZN => n26582);
   U1207 : OAI22_X1 port map( A1 => n26631, A2 => n23895, B1 => n23634, B2 => 
                           n26596, ZN => n26581);
   U1208 : AOI211_X1 port map( C1 => n24082, C2 => n26627, A => n26582, B => 
                           n26581, ZN => n26632);
   U1209 : INV_X1 port map( A => n26631, ZN => n26599);
   U1210 : AOI22_X1 port map( A1 => n24153, A2 => n24134, B1 => n23955, B2 => 
                           n23702, ZN => n26583);
   U1211 : OAI211_X1 port map( C1 => n24156, C2 => n23930, A => n23694, B => 
                           n26583, ZN => n26585);
   U1212 : AOI222_X1 port map( A1 => n26586, A2 => n24097, B1 => n26585, B2 => 
                           n23967, C1 => n26584, C2 => n24038, ZN => n26587);
   U1213 : OAI22_X1 port map( A1 => n23633, A2 => n26588, B1 => n24113, B2 => 
                           n26587, ZN => n26592);
   U1214 : OAI22_X1 port map( A1 => n24108, A2 => n26590, B1 => n23891, B2 => 
                           n26589, ZN => n26591);
   U1215 : AOI211_X1 port map( C1 => n23963, C2 => n26593, A => n26592, B => 
                           n26591, ZN => n26595);
   U1216 : OAI22_X1 port map( A1 => n24112, A2 => n26595, B1 => n23635, B2 => 
                           n26594, ZN => n26598);
   U1217 : OAI22_X1 port map( A1 => n23895, A2 => n26625, B1 => n24121, B2 => 
                           n26596, ZN => n26597);
   U1218 : AOI211_X1 port map( C1 => n24082, C2 => n26599, A => n26598, B => 
                           n26597, ZN => n26600);
   U1219 : OAI222_X1 port map( A1 => n26623, A2 => n24071, B1 => n26632, B2 => 
                           n24103, C1 => n23965, C2 => n26600, ZN => n26642);
   U1220 : AOI22_X1 port map( A1 => n23963, A2 => n26611, B1 => n24104, B2 => 
                           n26604, ZN => n26602);
   U1221 : AOI22_X1 port map( A1 => n24123, A2 => n26613, B1 => n23887, B2 => 
                           n26605, ZN => n26601);
   U1222 : OAI211_X1 port map( C1 => n24108, C2 => n26603, A => n26602, B => 
                           n26601, ZN => n26646);
   U1223 : AOI22_X1 port map( A1 => n24069, A2 => n26612, B1 => n27677, B2 => 
                           n26604, ZN => n26607);
   U1224 : AOI22_X1 port map( A1 => n23630, A2 => n26613, B1 => n24061, B2 => 
                           n26605, ZN => n26606);
   U1225 : OAI211_X1 port map( C1 => n26608, C2 => n27661, A => n26607, B => 
                           n26606, ZN => n26624);
   U1226 : AOI22_X1 port map( A1 => n24082, A2 => n26646, B1 => n24094, B2 => 
                           n26624, ZN => n26610);
   U1227 : AOI22_X1 port map( A1 => n24093, A2 => n26627, B1 => n23632, B2 => 
                           n26628, ZN => n26609);
   U1228 : OAI211_X1 port map( C1 => n24112, C2 => n26631, A => n26610, B => 
                           n26609, ZN => n26639);
   U1229 : AOI22_X1 port map( A1 => n23963, A2 => n26910, B1 => n24104, B2 => 
                           n26611, ZN => n26615);
   U1230 : AOI22_X1 port map( A1 => n23887, A2 => n26613, B1 => n27666, B2 => 
                           n26612, ZN => n26614);
   U1231 : OAI211_X1 port map( C1 => n24108, C2 => n26616, A => n26615, B => 
                           n26614, ZN => n26645);
   U1232 : AOI22_X1 port map( A1 => n26624, A2 => n27708, B1 => n27665, B2 => 
                           n26645, ZN => n26618);
   U1233 : AOI22_X1 port map( A1 => n24092, A2 => n26628, B1 => n26646, B2 => 
                           n27675, ZN => n26617);
   U1234 : OAI211_X1 port map( C1 => n26619, C2 => n24064, A => n26618, B => 
                           n26617, ZN => n26635);
   U1235 : INV_X1 port map( A => n26628, ZN => n26622);
   U1236 : AOI22_X1 port map( A1 => n24094, A2 => n26645, B1 => n27665, B2 => 
                           n26813, ZN => n26621);
   U1237 : AOI22_X1 port map( A1 => n23632, A2 => n26646, B1 => n24066, B2 => 
                           n26624, ZN => n26620);
   U1238 : OAI211_X1 port map( C1 => n26622, C2 => n27674, A => n26621, B => 
                           n26620, ZN => n26781);
   U1239 : AOI222_X1 port map( A1 => n26639, A2 => n24084, B1 => n26635, B2 => 
                           n23975, C1 => n26781, C2 => n23970, ZN => n26652);
   U1240 : INV_X1 port map( A => n26623, ZN => n26633);
   U1241 : INV_X1 port map( A => n26624, ZN => n26647);
   U1242 : OAI22_X1 port map( A1 => n24112, A2 => n26625, B1 => n26647, B2 => 
                           n24034, ZN => n26626);
   U1243 : INV_X1 port map( A => n26626, ZN => n26630);
   U1244 : AOI22_X1 port map( A1 => n24095, A2 => n26628, B1 => n26627, B2 => 
                           n27706, ZN => n26629);
   U1245 : OAI211_X1 port map( C1 => n26631, C2 => n23634, A => n26630, B => 
                           n26629, ZN => n26636);
   U1246 : AOI222_X1 port map( A1 => n26633, A2 => n24084, B1 => n26639, B2 => 
                           n23970, C1 => n26636, C2 => n23975, ZN => n26644);
   U1247 : OAI22_X1 port map( A1 => n26652, A2 => n24098, B1 => n26644, B2 => 
                           n23977, ZN => n26641);
   U1248 : INV_X1 port map( A => n26632, ZN => n26634);
   U1249 : AOI222_X1 port map( A1 => n26634, A2 => n24084, B1 => n26633, B2 => 
                           n23975, C1 => n26636, C2 => n23970, ZN => n26655);
   U1250 : INV_X1 port map( A => n26635, ZN => n26651);
   U1251 : INV_X1 port map( A => n26636, ZN => n26637);
   U1252 : OAI22_X1 port map( A1 => n26651, A2 => n24070, B1 => n26637, B2 => 
                           n23966, ZN => n26638);
   U1253 : AOI21_X1 port map( B1 => n23975, B2 => n26639, A => n26638, ZN => 
                           n26643);
   U1254 : OAI22_X1 port map( A1 => n26655, A2 => n24091, B1 => n26643, B2 => 
                           n23893, ZN => n26640);
   U1255 : AOI211_X1 port map( C1 => n23888, C2 => n26642, A => n26641, B => 
                           n26640, ZN => n26657);
   U1256 : INV_X1 port map( A => n26643, ZN => n26728);
   U1257 : INV_X1 port map( A => n26644, ZN => n26714);
   U1258 : AOI22_X1 port map( A1 => n24096, A2 => n26728, B1 => n27702, B2 => 
                           n26714, ZN => n26654);
   U1259 : INV_X1 port map( A => n26781, ZN => n26650);
   U1260 : INV_X1 port map( A => n26645, ZN => n26824);
   U1261 : OAI22_X1 port map( A1 => n26824, A2 => n24122, B1 => n26822, B2 => 
                           n27681, ZN => n26649);
   U1262 : INV_X1 port map( A => n26646, ZN => n26814);
   U1263 : OAI22_X1 port map( A1 => n24112, A2 => n26647, B1 => n26814, B2 => 
                           n23635, ZN => n26648);
   U1264 : AOI211_X1 port map( C1 => n27675, C2 => n26813, A => n26649, B => 
                           n26648, ZN => n26799);
   U1265 : OAI222_X1 port map( A1 => n26651, A2 => n23966, B1 => n26650, B2 => 
                           n24103, C1 => n24110, C2 => n26799, ZN => n26766);
   U1266 : INV_X1 port map( A => n26652, ZN => n26746);
   U1267 : AOI22_X1 port map( A1 => n23976, A2 => n26766, B1 => n24099, B2 => 
                           n26746, ZN => n26653);
   U1268 : OAI211_X1 port map( C1 => n26655, C2 => n27705, A => n26654, B => 
                           n26653, ZN => n26662);
   U1269 : NAND3_X1 port map( A1 => n24012, A2 => n24167, A3 => n26662, ZN => 
                           n26656);
   U1270 : OAI211_X1 port map( C1 => n24029, C2 => n26657, A => n23693, B => 
                           n26656, ZN => OUTALU(31));
   U1271 : AOI22_X1 port map( A1 => DATA2(30), A2 => n26981, B1 => n26847, B2 
                           => n1830, ZN => n26660);
   U1272 : INV_X1 port map( A => DATA2(30), ZN => n27251);
   U1273 : AOI22_X1 port map( A1 => DATA1(30), A2 => n27251, B1 => DATA2(30), 
                           B2 => n27205, ZN => n27120);
   U1274 : INV_X1 port map( A => n27120, ZN => n27199);
   U1275 : AOI22_X1 port map( A1 => n23766, A2 => n27567, B1 => n27557, B2 => 
                           n27199, ZN => n26659);
   U1276 : NAND3_X1 port map( A1 => DATA1(31), A2 => n1830, A3 => n26848, ZN =>
                           n26658);
   U1277 : OAI211_X1 port map( C1 => n26660, C2 => n27205, A => n26659, B => 
                           n26658, ZN => n18935);
   U1278 : NOR3_X1 port map( A1 => n1814, A2 => n26661, A3 => n27710, ZN => 
                           n19182);
   U1279 : NAND3_X1 port map( A1 => n1814, A2 => n26661, A3 => n26710, ZN => 
                           n19268);
   U1280 : AOI21_X1 port map( B1 => n26662, B2 => n24086, A => n23929, ZN => 
                           n26663);
   U1281 : NAND2_X1 port map( A1 => n23928, A2 => n26663, ZN => n26664);
   U1282 : NOR2_X1 port map( A1 => n26664, A2 => n23691, ZN => n26665);
   U1283 : OAI21_X1 port map( B1 => n24159, B2 => n24114, A => n26665, ZN => 
                           OUTALU(30));
   U1284 : NOR2_X1 port map( A1 => n24165, A2 => n26666, ZN => n26668);
   U1285 : AOI211_X1 port map( C1 => n26724, C2 => n24173, A => n26668, B => 
                           n26667, ZN => n18934);
   U1286 : AOI211_X1 port map( C1 => n26671, C2 => n26670, A => n26669, B => 
                           n27036, ZN => n26679);
   U1287 : NAND2_X1 port map( A1 => DATA2(2), A2 => n24049, ZN => n26677);
   U1288 : OAI211_X1 port map( C1 => n26674, C2 => n26673, A => n27040, B => 
                           n26672, ZN => n26676);
   U1289 : AOI22_X1 port map( A1 => DATA2(2), A2 => n24049, B1 => n24165, B2 =>
                           n27592, ZN => n27127);
   U1290 : NAND2_X1 port map( A1 => n27127, A2 => n27557, ZN => n26675);
   U1291 : OAI211_X1 port map( C1 => n27549, C2 => n26677, A => n26676, B => 
                           n26675, ZN => n26678);
   U1292 : AOI211_X1 port map( C1 => n23936, C2 => n27567, A => n26679, B => 
                           n26678, ZN => n18933);
   U1293 : OAI22_X1 port map( A1 => n26857, A2 => n27638, B1 => n26853, B2 => 
                           n25891, ZN => n26681);
   U1294 : OAI22_X1 port map( A1 => n27641, A2 => n26854, B1 => n26425, B2 => 
                           n27640, ZN => n26680);
   U1295 : AOI211_X1 port map( C1 => n27632, C2 => n22526, A => n26681, B => 
                           n26680, ZN => n1806);
   U1296 : OAI22_X1 port map( A1 => n23893, A2 => n26861, B1 => n23977, B2 => 
                           n27212, ZN => n26699);
   U1297 : INV_X1 port map( A => n26862, ZN => n27223);
   U1298 : NAND2_X1 port map( A1 => n24118, A2 => n24107, ZN => n26682);
   U1299 : OAI21_X1 port map( B1 => n23954, B2 => n24140, A => n26682, ZN => 
                           n26684);
   U1300 : OAI22_X1 port map( A1 => n24156, A2 => n23687, B1 => n23957, B2 => 
                           n24139, ZN => n26683);
   U1301 : AOI211_X1 port map( C1 => n27667, C2 => n27223, A => n26684, B => 
                           n26683, ZN => n27225);
   U1302 : OAI222_X1 port map( A1 => n23979, A2 => n26864, B1 => n26685, B2 => 
                           n24080, C1 => n24105, C2 => n27225, ZN => n27218);
   U1303 : INV_X1 port map( A => n27218, ZN => n26867);
   U1304 : INV_X1 port map( A => n26686, ZN => n26871);
   U1305 : AOI22_X1 port map( A1 => n27666, A2 => n26687, B1 => n26871, B2 => 
                           n24069, ZN => n26690);
   U1306 : AOI22_X1 port map( A1 => n27227, A2 => n23630, B1 => n26688, B2 => 
                           n23963, ZN => n26689);
   U1307 : OAI211_X1 port map( C1 => n27661, C2 => n26867, A => n26690, B => 
                           n26689, ZN => n27214);
   U1308 : INV_X1 port map( A => n27214, ZN => n26694);
   U1309 : AOI22_X1 port map( A1 => n24094, A2 => n26872, B1 => n27665, B2 => 
                           n26691, ZN => n26693);
   U1310 : AOI22_X1 port map( A1 => n24092, A2 => n26873, B1 => n23631, B2 => 
                           n27215, ZN => n26692);
   U1311 : OAI211_X1 port map( C1 => n26694, C2 => n27674, A => n26693, B => 
                           n26692, ZN => n27238);
   U1312 : AOI22_X1 port map( A1 => n24084, A2 => n27238, B1 => n23970, B2 => 
                           n26695, ZN => n26696);
   U1313 : INV_X1 port map( A => n26696, ZN => n26697);
   U1314 : AOI21_X1 port map( B1 => n26876, B2 => n23975, A => n26697, ZN => 
                           n27241);
   U1315 : OAI22_X1 port map( A1 => n24091, A2 => n27213, B1 => n27241, B2 => 
                           n24111, ZN => n26698);
   U1316 : OAI21_X1 port map( B1 => n26699, B2 => n26698, A => n24085, ZN => 
                           n26700);
   U1317 : OAI211_X1 port map( C1 => n24029, C2 => n23690, A => n23689, B => 
                           n26700, ZN => OUTALU(2));
   U1318 : NOR2_X1 port map( A1 => DATA2(29), A2 => n26703, ZN => n27200);
   U1319 : NAND2_X1 port map( A1 => DATA2(29), A2 => n26703, ZN => n27201);
   U1320 : INV_X1 port map( A => n27201, ZN => n26701);
   U1321 : NOR2_X1 port map( A1 => n27200, A2 => n26701, ZN => n27044);
   U1322 : INV_X1 port map( A => n27044, ZN => n26702);
   U1323 : AOI22_X1 port map( A1 => n27567, A2 => n23769, B1 => n27557, B2 => 
                           n26702, ZN => n18930);
   U1324 : OAI21_X1 port map( B1 => n26703, B2 => n27033, A => n27018, ZN => 
                           n26709);
   U1325 : NAND2_X1 port map( A1 => DATA1(29), A2 => n26719, ZN => n26706);
   U1326 : NAND2_X1 port map( A1 => DATA1(30), A2 => n26704, ZN => n26705);
   U1327 : OAI211_X1 port map( C1 => n26707, C2 => n26732, A => n26706, B => 
                           n26705, ZN => n26708);
   U1328 : AOI22_X1 port map( A1 => DATA2(29), A2 => n26709, B1 => n1830, B2 =>
                           n26708, ZN => n18929);
   U1329 : INV_X1 port map( A => n26710, ZN => n26711);
   U1330 : AOI21_X1 port map( B1 => n26713, B2 => n26712, A => n26711, ZN => 
                           n19181);
   U1331 : AOI22_X1 port map( A1 => n23892, A2 => n26728, B1 => n24096, B2 => 
                           n26746, ZN => n26716);
   U1332 : AOI22_X1 port map( A1 => n24099, A2 => n26766, B1 => n23888, B2 => 
                           n26714, ZN => n26715);
   U1333 : AOI21_X1 port map( B1 => n26716, B2 => n26715, A => n24029, ZN => 
                           n26717);
   U1334 : AOI211_X1 port map( C1 => n24162, C2 => n23959, A => n23927, B => 
                           n26717, ZN => n26718);
   U1335 : NAND3_X1 port map( A1 => n23686, A2 => n23685, A3 => n26718, ZN => 
                           OUTALU(29));
   U1336 : INV_X1 port map( A => DATA2(28), ZN => n27253);
   U1337 : NOR3_X1 port map( A1 => n27549, A2 => n27253, A3 => n27198, ZN => 
                           n26727);
   U1338 : AOI22_X1 port map( A1 => DATA1(28), A2 => n27253, B1 => DATA2(28), 
                           B2 => n27198, ZN => n27192);
   U1339 : NAND2_X1 port map( A1 => DATA1(28), A2 => n26719, ZN => n26721);
   U1340 : OAI211_X1 port map( C1 => n26722, C2 => n26732, A => n26721, B => 
                           n26720, ZN => n26723);
   U1341 : AOI21_X1 port map( B1 => DATA1(30), B2 => n26724, A => n26723, ZN =>
                           n26725);
   U1342 : OAI22_X1 port map( A1 => n27192, A2 => n27570, B1 => n26725, B2 => 
                           n26811, ZN => n26726);
   U1343 : AOI211_X1 port map( C1 => n27542, C2 => n23772, A => n26727, B => 
                           n26726, ZN => n18927);
   U1344 : AOI222_X1 port map( A1 => n26766, A2 => n24096, B1 => n26728, B2 => 
                           n23888, C1 => n26746, C2 => n23892, ZN => n26729);
   U1345 : OAI211_X1 port map( C1 => n24029, C2 => n26729, A => n23684, B => 
                           n24028, ZN => OUTALU(28));
   U1346 : OAI22_X1 port map( A1 => n26736, A2 => n27660, B1 => n26735, B2 => 
                           n27658, ZN => n26744);
   U1347 : OAI211_X1 port map( C1 => n26750, C2 => n26732, A => n26731, B => 
                           n26730, ZN => n26733);
   U1348 : AOI211_X1 port map( C1 => n26753, C2 => DATA1(30), A => n26734, B =>
                           n26733, ZN => n26768);
   U1349 : NOR3_X1 port map( A1 => n26768, A2 => n26769, A3 => n26811, ZN => 
                           n26743);
   U1350 : AOI22_X1 port map( A1 => n26786, A2 => n26736, B1 => n26788, B2 => 
                           n26735, ZN => n26741);
   U1351 : NOR2_X1 port map( A1 => DATA2(27), A2 => n26737, ZN => n27194);
   U1352 : INV_X1 port map( A => n27194, ZN => n26738);
   U1353 : NAND2_X1 port map( A1 => DATA2(27), A2 => n26737, ZN => n27195);
   U1354 : NAND2_X1 port map( A1 => n26738, A2 => n27195, ZN => n27058);
   U1355 : AOI22_X1 port map( A1 => n27567, A2 => n23777, B1 => n27557, B2 => 
                           n27058, ZN => n26740);
   U1356 : NAND3_X1 port map( A1 => DATA2(27), A2 => DATA1(27), A3 => n26981, 
                           ZN => n26739);
   U1357 : OAI211_X1 port map( C1 => n26741, C2 => n26745, A => n26740, B => 
                           n26739, ZN => n26742);
   U1358 : AOI211_X1 port map( C1 => n26745, C2 => n26744, A => n26743, B => 
                           n26742, ZN => n18926);
   U1359 : AOI22_X1 port map( A1 => n23892, A2 => n26766, B1 => n23888, B2 => 
                           n26746, ZN => n26747);
   U1360 : OAI21_X1 port map( B1 => n24029, B2 => n26747, A => n23683, ZN => 
                           OUTALU(27));
   U1361 : OAI211_X1 port map( C1 => n26750, C2 => n27205, A => n26749, B => 
                           n26748, ZN => n26751);
   U1362 : AOI211_X1 port map( C1 => n26753, C2 => DATA1(29), A => n26752, B =>
                           n26751, ZN => n26790);
   U1363 : OAI22_X1 port map( A1 => n26768, A2 => n26754, B1 => n26790, B2 => 
                           n26769, ZN => n26755);
   U1364 : NAND2_X1 port map( A1 => n1830, A2 => n26755, ZN => n19267);
   U1365 : AND2_X1 port map( A1 => n26757, A2 => n26756, ZN => n26760);
   U1366 : AOI211_X1 port map( C1 => n26760, C2 => n26770, A => n26758, B => 
                           n27660, ZN => n26765);
   U1367 : INV_X1 port map( A => DATA2(26), ZN => n27255);
   U1368 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2(26), B1 => n27255, 
                           B2 => n27191, ZN => n27186);
   U1369 : INV_X1 port map( A => n27186, ZN => n27074);
   U1370 : NAND3_X1 port map( A1 => DATA2(26), A2 => DATA1(26), A3 => n26981, 
                           ZN => n26763);
   U1371 : AOI211_X1 port map( C1 => n26775, C2 => n26760, A => n27658, B => 
                           n26759, ZN => n26761);
   U1372 : INV_X1 port map( A => n26761, ZN => n26762);
   U1373 : OAI211_X1 port map( C1 => n27074, C2 => n27570, A => n26763, B => 
                           n26762, ZN => n26764);
   U1374 : AOI211_X1 port map( C1 => n27542, C2 => n23781, A => n26765, B => 
                           n26764, ZN => n18925);
   U1375 : NAND3_X1 port map( A1 => n23888, A2 => n24086, A3 => n26766, ZN => 
                           n26767);
   U1376 : NAND3_X1 port map( A1 => n24017, A2 => n23682, A3 => n26767, ZN => 
                           OUTALU(26));
   U1377 : OAI222_X1 port map( A1 => n26769, A2 => n26791, B1 => n26792, B2 => 
                           n26790, C1 => n26446, C2 => n26768, ZN => n26827);
   U1378 : NAND3_X1 port map( A1 => n1830, A2 => n27624, A3 => n26827, ZN => 
                           n19180);
   U1379 : INV_X1 port map( A => n26776, ZN => n26772);
   U1380 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n26785);
   U1381 : INV_X1 port map( A => n26770, ZN => n26771);
   U1382 : AOI211_X1 port map( C1 => n26772, C2 => n26785, A => n26771, B => 
                           n27660, ZN => n26780);
   U1383 : NOR2_X1 port map( A1 => DATA2(25), A2 => n26773, ZN => n27187);
   U1384 : NAND2_X1 port map( A1 => DATA2(25), A2 => n26773, ZN => n27188);
   U1385 : INV_X1 port map( A => n27188, ZN => n26774);
   U1386 : NOR2_X1 port map( A1 => n27187, A2 => n26774, ZN => n27062);
   U1387 : OAI211_X1 port map( C1 => n26776, C2 => n26784, A => n26788, B => 
                           n26775, ZN => n26778);
   U1388 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n26981, 
                           ZN => n26777);
   U1389 : OAI211_X1 port map( C1 => n27062, C2 => n27570, A => n26778, B => 
                           n26777, ZN => n26779);
   U1390 : AOI211_X1 port map( C1 => n27542, C2 => n23785, A => n26780, B => 
                           n26779, ZN => n19179);
   U1391 : INV_X1 port map( A => n26799, ZN => n26782);
   U1392 : AOI22_X1 port map( A1 => n23975, A2 => n26782, B1 => n24065, B2 => 
                           n26781, ZN => n26783);
   U1393 : OAI211_X1 port map( C1 => n24029, C2 => n26783, A => n23926, B => 
                           n23681, ZN => OUTALU(25));
   U1394 : NAND3_X1 port map( A1 => n26786, A2 => n26785, A3 => n26784, ZN => 
                           n19178);
   U1395 : NAND2_X1 port map( A1 => n26788, A2 => n26787, ZN => n19266);
   U1396 : AOI22_X1 port map( A1 => DATA2(24), A2 => n27652, B1 => 
                           DATA2_I_24_port, B2 => n26788, ZN => n26789);
   U1397 : AOI21_X1 port map( B1 => n26789, B2 => n27018, A => n27185, ZN => 
                           n26798);
   U1398 : INV_X1 port map( A => DATA2(24), ZN => n27257);
   U1399 : AOI22_X1 port map( A1 => DATA1(24), A2 => DATA2(24), B1 => n27257, 
                           B2 => n27185, ZN => n27180);
   U1400 : INV_X1 port map( A => n27180, ZN => n27057);
   U1401 : OAI222_X1 port map( A1 => n26794, A2 => n26793, B1 => n26792, B2 => 
                           n26791, C1 => n26446, C2 => n26790, ZN => n27617);
   U1402 : AOI22_X1 port map( A1 => n25892, A2 => n26827, B1 => n26795, B2 => 
                           n27617, ZN => n26796);
   U1403 : OAI22_X1 port map( A1 => n27057, A2 => n27570, B1 => n26796, B2 => 
                           n26811, ZN => n26797);
   U1404 : AOI211_X1 port map( C1 => n23789, C2 => n27542, A => n26798, B => 
                           n26797, ZN => n22091);
   U1405 : OR3_X1 port map( A1 => n26799, A2 => n23966, A3 => n24029, ZN => 
                           n26800);
   U1406 : NAND4_X1 port map( A1 => n23680, A2 => n23925, A3 => n24016, A4 => 
                           n26800, ZN => OUTALU(24));
   U1407 : AOI21_X1 port map( B1 => DATA2(23), B2 => n27652, A => n27651, ZN =>
                           n19176);
   U1408 : NAND2_X1 port map( A1 => n22313, A2 => n23793, ZN => n19265);
   U1409 : AOI222_X1 port map( A1 => n27619, A2 => n27624, B1 => n27617, B2 => 
                           n25892, C1 => n26827, C2 => n1857, ZN => n26812);
   U1410 : NOR2_X1 port map( A1 => DATA2(23), A2 => n1840, ZN => n27181);
   U1411 : INV_X1 port map( A => n27181, ZN => n26801);
   U1412 : NAND2_X1 port map( A1 => DATA2(23), A2 => n1840, ZN => n27182);
   U1413 : NAND2_X1 port map( A1 => n26801, A2 => n27182, ZN => n27059);
   U1414 : AOI21_X1 port map( B1 => n26802, B2 => n26804, A => n26807, ZN => 
                           n26803);
   U1415 : AOI211_X1 port map( C1 => n26807, C2 => n26804, A => n27710, B => 
                           n26803, ZN => n26805);
   U1416 : AOI21_X1 port map( B1 => n27557, B2 => n27059, A => n26805, ZN => 
                           n26810);
   U1417 : NAND3_X1 port map( A1 => n26808, A2 => n26807, A3 => n26806, ZN => 
                           n26809);
   U1418 : OAI211_X1 port map( C1 => n26812, C2 => n26811, A => n26810, B => 
                           n26809, ZN => n18923);
   U1419 : INV_X1 port map( A => n26813, ZN => n26823);
   U1420 : OAI22_X1 port map( A1 => n23895, A2 => n26822, B1 => n26823, B2 => 
                           n24122, ZN => n26816);
   U1421 : OAI22_X1 port map( A1 => n24112, A2 => n26814, B1 => n26824, B2 => 
                           n23635, ZN => n26815);
   U1422 : AOI221_X1 port map( B1 => n26816, B2 => n24086, C1 => n26815, C2 => 
                           n24086, A => n23679, ZN => n26817);
   U1423 : OAI211_X1 port map( C1 => n23924, C2 => n24163, A => n24015, B => 
                           n26817, ZN => OUTALU(23));
   U1424 : AOI22_X1 port map( A1 => DATA1(22), A2 => n27259, B1 => DATA2(22), 
                           B2 => n27177, ZN => n27179);
   U1425 : INV_X1 port map( A => n27179, ZN => n26818);
   U1426 : AOI22_X1 port map( A1 => n23797, A2 => n27567, B1 => n27557, B2 => 
                           n26818, ZN => n18922);
   U1427 : AOI22_X1 port map( A1 => n27632, A2 => n27617, B1 => n27624, B2 => 
                           n27620, ZN => n26819);
   U1428 : OAI21_X1 port map( B1 => n26820, B2 => n27607, A => n26819, ZN => 
                           n26821);
   U1429 : AOI21_X1 port map( B1 => n27709, B2 => n26827, A => n26821, ZN => 
                           n19174);
   U1430 : OAI222_X1 port map( A1 => n24112, A2 => n26824, B1 => n26823, B2 => 
                           n23635, C1 => n24122, C2 => n26822, ZN => n26825);
   U1431 : AOI211_X1 port map( C1 => n24086, C2 => n26825, A => n23923, B => 
                           n23951, ZN => n26826);
   U1432 : OAI211_X1 port map( C1 => n24036, C2 => n23922, A => n23678, B => 
                           n26826, ZN => OUTALU(22));
   U1433 : AOI22_X1 port map( A1 => n25892, A2 => n27620, B1 => n27709, B2 => 
                           n27617, ZN => n26829);
   U1434 : AOI22_X1 port map( A1 => n27632, A2 => n27619, B1 => n26827, B2 => 
                           n27645, ZN => n26828);
   U1435 : OAI211_X1 port map( C1 => n27641, C2 => n27616, A => n26829, B => 
                           n26828, ZN => n18921);
   U1436 : NAND3_X1 port map( A1 => n1858, A2 => n1830, A3 => n18921, ZN => 
                           n12313);
   U1437 : AOI211_X1 port map( C1 => n26832, C2 => n26831, A => n26830, B => 
                           n26919, ZN => n26840);
   U1438 : INV_X1 port map( A => DATA2(20), ZN => n27261);
   U1439 : NAND2_X1 port map( A1 => DATA1(20), A2 => n27261, ZN => n27173);
   U1440 : NAND2_X1 port map( A1 => DATA2(20), A2 => n26833, ZN => n27176);
   U1441 : AND2_X1 port map( A1 => n27173, A2 => n27176, ZN => n27055);
   U1442 : OAI211_X1 port map( C1 => n26836, C2 => n26835, A => n27648, B => 
                           n26834, ZN => n26838);
   U1443 : NAND3_X1 port map( A1 => DATA2(20), A2 => DATA1(20), A3 => n26981, 
                           ZN => n26837);
   U1444 : OAI211_X1 port map( C1 => n27055, C2 => n27570, A => n26838, B => 
                           n26837, ZN => n26839);
   U1445 : AOI211_X1 port map( C1 => n27542, C2 => n23805, A => n26840, B => 
                           n26839, ZN => n19172);
   U1446 : AOI22_X1 port map( A1 => n24101, A2 => n24126, B1 => n24060, B2 => 
                           n23677, ZN => n26843);
   U1447 : NAND3_X1 port map( A1 => n23962, A2 => n24086, A3 => n26841, ZN => 
                           n26842);
   U1448 : OAI211_X1 port map( C1 => n24036, C2 => n26843, A => n23676, B => 
                           n26842, ZN => OUTALU(20));
   U1449 : AOI211_X1 port map( C1 => n27034, C2 => n26849, A => n26844, B => 
                           n27036, ZN => n26846);
   U1450 : NOR2_X1 port map( A1 => n24175, A2 => n27571, ZN => n27125);
   U1451 : NAND2_X1 port map( A1 => n24175, A2 => n27571, ZN => n27080);
   U1452 : INV_X1 port map( A => n27080, ZN => n27126);
   U1453 : NOR2_X1 port map( A1 => n27125, A2 => n27126, ZN => n27045);
   U1454 : NOR2_X1 port map( A1 => n27045, A2 => n27570, ZN => n26845);
   U1455 : AOI211_X1 port map( C1 => n23591, C2 => n27542, A => n26846, B => 
                           n26845, ZN => n18920);
   U1456 : AOI21_X1 port map( B1 => n26847, B2 => n1831, A => n27651, ZN => 
                           n27032);
   U1457 : OAI21_X1 port map( B1 => n27571, B2 => n27033, A => n27032, ZN => 
                           n19171);
   U1458 : NAND3_X1 port map( A1 => n24173, A2 => n26848, A3 => n1831, ZN => 
                           n19170);
   U1459 : INV_X1 port map( A => n26849, ZN => n26851);
   U1460 : OAI221_X1 port map( B1 => n27035, B2 => n26851, C1 => n26850, C2 => 
                           n26849, A => n27040, ZN => n18860);
   U1461 : OAI22_X1 port map( A1 => n27641, A2 => n26852, B1 => n26425, B2 => 
                           n26857, ZN => n26856);
   U1462 : OAI22_X1 port map( A1 => n26854, A2 => n27607, B1 => n26853, B2 => 
                           n27636, ZN => n26855);
   U1463 : AOI211_X1 port map( C1 => n27709, C2 => n22526, A => n26856, B => 
                           n26855, ZN => n22532);
   U1464 : OAI22_X1 port map( A1 => n26425, A2 => n27637, B1 => n27635, B2 => 
                           n27638, ZN => n26859);
   U1465 : OAI22_X1 port map( A1 => n26857, A2 => n27607, B1 => n27640, B2 => 
                           n27636, ZN => n26858);
   U1466 : AOI211_X1 port map( C1 => n27624, C2 => n22526, A => n26859, B => 
                           n26858, ZN => n1817);
   U1467 : OAI22_X1 port map( A1 => n1817, A2 => n1859, B1 => n26860, B2 => 
                           n1836, ZN => n18918);
   U1468 : INV_X1 port map( A => n27241, ZN => n26879);
   U1469 : OAI22_X1 port map( A1 => n23893, A2 => n27212, B1 => n26861, B2 => 
                           n27707, ZN => n26878);
   U1470 : INV_X1 port map( A => n27225, ZN => n26866);
   U1471 : OAI22_X1 port map( A1 => n23954, A2 => n26862, B1 => n24156, B2 => 
                           n23674, ZN => n26863);
   U1472 : AOI211_X1 port map( C1 => n25864, C2 => n24060, A => n23673, B => 
                           n26863, ZN => n27226);
   U1473 : OAI22_X1 port map( A1 => n24080, A2 => n26864, B1 => n24105, B2 => 
                           n27226, ZN => n26865);
   U1474 : AOI21_X1 port map( B1 => n27662, B2 => n26866, A => n26865, ZN => 
                           n27217);
   U1475 : OAI22_X1 port map( A1 => n26867, A2 => n27676, B1 => n27217, B2 => 
                           n27661, ZN => n26870);
   U1476 : OAI22_X1 port map( A1 => n23891, A2 => n26868, B1 => n27231, B2 => 
                           n27672, ZN => n26869);
   U1477 : AOI211_X1 port map( C1 => n23964, C2 => n26871, A => n26870, B => 
                           n26869, ZN => n27216);
   U1478 : AOI22_X1 port map( A1 => n24075, A2 => n26872, B1 => n27684, B2 => 
                           n27215, ZN => n26875);
   U1479 : AOI22_X1 port map( A1 => n24093, A2 => n27214, B1 => n23631, B2 => 
                           n26873, ZN => n26874);
   U1480 : OAI211_X1 port map( C1 => n27216, C2 => n27674, A => n26875, B => 
                           n26874, ZN => n27239);
   U1481 : AOI222_X1 port map( A1 => n27238, A2 => n23975, B1 => n26876, B2 => 
                           n23971, C1 => n27239, C2 => n24073, ZN => n27211);
   U1482 : OAI22_X1 port map( A1 => n23977, A2 => n27213, B1 => n24074, B2 => 
                           n27211, ZN => n26877);
   U1483 : AOI211_X1 port map( C1 => n27702, C2 => n26879, A => n26878, B => 
                           n26877, ZN => n27248);
   U1484 : INV_X1 port map( A => n27248, ZN => n26880);
   U1485 : AOI22_X1 port map( A1 => n24174, A2 => n23920, B1 => n24085, B2 => 
                           n26880, ZN => n26881);
   U1486 : NAND4_X1 port map( A1 => n23612, A2 => n23675, A3 => n23919, A4 => 
                           n26881, ZN => OUTALU(1));
   U1487 : INV_X1 port map( A => n26884, ZN => n26883);
   U1488 : INV_X1 port map( A => n26919, ZN => n27649);
   U1489 : AOI22_X1 port map( A1 => n26883, A2 => n27649, B1 => n27648, B2 => 
                           n26882, ZN => n26888);
   U1490 : AOI22_X1 port map( A1 => n27648, A2 => n26885, B1 => n27649, B2 => 
                           n26884, ZN => n26887);
   U1491 : INV_X1 port map( A => n26889, ZN => n26886);
   U1492 : AOI22_X1 port map( A1 => n26889, A2 => n26888, B1 => n26887, B2 => 
                           n26886, ZN => n18917);
   U1493 : INV_X1 port map( A => DATA2(19), ZN => n27262);
   U1494 : NAND2_X1 port map( A1 => DATA1(19), A2 => n27262, ZN => n27172);
   U1495 : NOR2_X1 port map( A1 => n27262, A2 => DATA1(19), ZN => n27166);
   U1496 : INV_X1 port map( A => n27166, ZN => n27109);
   U1497 : AND2_X1 port map( A1 => n27172, A2 => n27109, ZN => n27064);
   U1498 : OAI21_X1 port map( B1 => n27262, B2 => n27033, A => n27018, ZN => 
                           n26890);
   U1499 : AOI22_X1 port map( A1 => DATA1(19), A2 => n26890, B1 => n27542, B2 
                           => n23809, ZN => n26891);
   U1500 : OAI21_X1 port map( B1 => n27064, B2 => n27570, A => n26891, ZN => 
                           n19264);
   U1501 : AOI222_X1 port map( A1 => n24058, A2 => n23677, B1 => n24101, B2 => 
                           n25878, C1 => n24060, C2 => n24126, ZN => n26898);
   U1502 : OAI22_X1 port map( A1 => n26893, A2 => n27661, B1 => n26892, B2 => 
                           n27676, ZN => n26894);
   U1503 : AOI21_X1 port map( B1 => n23630, B2 => n26923, A => n26894, ZN => 
                           n26895);
   U1504 : OAI21_X1 port map( B1 => n26924, B2 => n27678, A => n26895, ZN => 
                           n26896);
   U1505 : AOI211_X1 port map( C1 => n27701, C2 => n26896, A => n23918, B => 
                           n23917, ZN => n26897);
   U1506 : OAI21_X1 port map( B1 => n24036, B2 => n26898, A => n26897, ZN => 
                           OUTALU(19));
   U1507 : OR2_X1 port map( A1 => n26900, A2 => n26899, ZN => n26905);
   U1508 : OAI211_X1 port map( C1 => n26905, C2 => n26920, A => n26901, B => 
                           n27649, ZN => n26902);
   U1509 : INV_X1 port map( A => n26902, ZN => n26909);
   U1510 : INV_X1 port map( A => DATA2(18), ZN => n27263);
   U1511 : NOR2_X1 port map( A1 => DATA1(18), A2 => n27263, ZN => n27167);
   U1512 : NOR2_X1 port map( A1 => DATA2(18), A2 => n26903, ZN => n27163);
   U1513 : NOR2_X1 port map( A1 => n27167, A2 => n27163, ZN => n27060);
   U1514 : OAI211_X1 port map( C1 => n26917, C2 => n26905, A => n27648, B => 
                           n26904, ZN => n26907);
   U1515 : NAND3_X1 port map( A1 => DATA2(18), A2 => DATA1(18), A3 => n26981, 
                           ZN => n26906);
   U1516 : OAI211_X1 port map( C1 => n27060, C2 => n27570, A => n26907, B => 
                           n26906, ZN => n26908);
   U1517 : AOI211_X1 port map( C1 => n27542, C2 => n23813, A => n26909, B => 
                           n26908, ZN => n18916);
   U1518 : INV_X1 port map( A => n26924, ZN => n26937);
   U1519 : AOI222_X1 port map( A1 => n26923, A2 => n24123, B1 => n26910, B2 => 
                           n23887, C1 => n26937, C2 => n23630, ZN => n26914);
   U1520 : AOI22_X1 port map( A1 => n24060, A2 => n25878, B1 => n23956, B2 => 
                           n23677, ZN => n26911);
   U1521 : OAI21_X1 port map( B1 => n24156, B2 => n25877, A => n26911, ZN => 
                           n26912);
   U1522 : OAI221_X1 port map( B1 => n26912, B2 => n24126, C1 => n26912, C2 => 
                           n24058, A => n24085, ZN => n26913);
   U1523 : OAI211_X1 port map( C1 => n24029, C2 => n26914, A => n23672, B => 
                           n26913, ZN => OUTALU(18));
   U1524 : NOR2_X1 port map( A1 => DATA2(17), A2 => n26915, ZN => n27105);
   U1525 : INV_X1 port map( A => n27105, ZN => n27169);
   U1526 : NAND2_X1 port map( A1 => DATA2(17), A2 => n26915, ZN => n27165);
   U1527 : NAND2_X1 port map( A1 => n27169, A2 => n27165, ZN => n27049);
   U1528 : AOI22_X1 port map( A1 => n27567, A2 => n23817, B1 => n27557, B2 => 
                           n27049, ZN => n18915);
   U1529 : AOI211_X1 port map( C1 => n26918, C2 => n26922, A => n26917, B => 
                           n26916, ZN => n18914);
   U1530 : AOI211_X1 port map( C1 => n26922, C2 => n26921, A => n26920, B => 
                           n26919, ZN => n18913);
   U1531 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n26981, 
                           ZN => n19169);
   U1532 : INV_X1 port map( A => n26923, ZN => n26925);
   U1533 : OAI22_X1 port map( A1 => n26925, A2 => n27661, B1 => n26924, B2 => 
                           n27676, ZN => n26926);
   U1534 : AOI211_X1 port map( C1 => n24086, C2 => n26926, A => n23670, B => 
                           n23669, ZN => n26929);
   U1535 : NAND3_X1 port map( A1 => n24051, A2 => n24085, A3 => n26927, ZN => 
                           n26928);
   U1536 : NAND4_X1 port map( A1 => n23671, A2 => n23916, A3 => n26929, A4 => 
                           n26928, ZN => OUTALU(17));
   U1537 : INV_X1 port map( A => DATA2(16), ZN => n27265);
   U1538 : NAND2_X1 port map( A1 => n27265, A2 => DATA1(16), ZN => n27159);
   U1539 : INV_X1 port map( A => n27159, ZN => n27107);
   U1540 : AOI21_X1 port map( B1 => DATA2(16), B2 => n26930, A => n27107, ZN =>
                           n27053);
   U1541 : INV_X1 port map( A => n27053, ZN => n26931);
   U1542 : AOI22_X1 port map( A1 => n27567, A2 => n23821, B1 => n27557, B2 => 
                           n26931, ZN => n18912);
   U1543 : OAI21_X1 port map( B1 => n27265, B2 => n27033, A => n27018, ZN => 
                           n26933);
   U1544 : AOI22_X1 port map( A1 => DATA1(16), A2 => n26933, B1 => n26932, B2 
                           => n27649, ZN => n18911);
   U1545 : OAI22_X1 port map( A1 => n24168, A2 => n26935, B1 => n23979, B2 => 
                           n26934, ZN => n26936);
   U1546 : AOI21_X1 port map( B1 => n24085, B2 => n26936, A => n24025, ZN => 
                           n26939);
   U1547 : NAND3_X1 port map( A1 => n23887, A2 => n24086, A3 => n26937, ZN => 
                           n26938);
   U1548 : NAND4_X1 port map( A1 => n23667, A2 => n23668, A3 => n26939, A4 => 
                           n26938, ZN => OUTALU(16));
   U1549 : INV_X1 port map( A => n26940, ZN => n26942);
   U1550 : INV_X1 port map( A => n26950, ZN => n26941);
   U1551 : AOI221_X1 port map( B1 => n26942, B2 => n26941, C1 => n26940, C2 => 
                           n26950, A => n1789, ZN => n26954);
   U1552 : AOI22_X1 port map( A1 => DATA1(15), A2 => n27266, B1 => DATA2(15), 
                           B2 => n26943, ZN => n27066);
   U1553 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n26944);
   U1554 : AND2_X1 port map( A1 => n26944, A2 => n17503, ZN => n27553);
   U1555 : OAI21_X1 port map( B1 => n27553, B2 => n26946, A => n26945, ZN => 
                           n26959);
   U1556 : NOR2_X1 port map( A1 => n26962, A2 => n26959, ZN => n26965);
   U1557 : OAI21_X1 port map( B1 => n26965, B2 => n26968, A => n26947, ZN => 
                           n26949);
   U1558 : AOI21_X1 port map( B1 => n26950, B2 => n26949, A => n27550, ZN => 
                           n26948);
   U1559 : OAI21_X1 port map( B1 => n26950, B2 => n26949, A => n26948, ZN => 
                           n26952);
   U1560 : NAND3_X1 port map( A1 => DATA2(15), A2 => DATA1(15), A3 => n26981, 
                           ZN => n26951);
   U1561 : OAI211_X1 port map( C1 => n27066, C2 => n27570, A => n26952, B => 
                           n26951, ZN => n26953);
   U1562 : AOI211_X1 port map( C1 => n27542, C2 => n23825, A => n26954, B => 
                           n26953, ZN => n18910);
   U1563 : INV_X1 port map( A => n26955, ZN => n26956);
   U1564 : AOI22_X1 port map( A1 => n24097, A2 => n26971, B1 => n24051, B2 => 
                           n26956, ZN => n26958);
   U1565 : NAND3_X1 port map( A1 => n23887, A2 => n24085, A3 => n26989, ZN => 
                           n26957);
   U1566 : OAI211_X1 port map( C1 => n24029, C2 => n26958, A => n23666, B => 
                           n26957, ZN => OUTALU(15));
   U1567 : OAI22_X1 port map( A1 => n26960, A2 => n1789, B1 => n27550, B2 => 
                           n26959, ZN => n26986);
   U1568 : INV_X1 port map( A => n26986, ZN => n26961);
   U1569 : NOR3_X1 port map( A1 => n26968, A2 => n26962, A3 => n26961, ZN => 
                           n19168);
   U1570 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_7_14_port, ZN =>
                           n26963);
   U1571 : NOR3_X1 port map( A1 => n24161, A2 => n23914, A3 => n26963, ZN => 
                           n3020);
   U1572 : AOI221_X1 port map( B1 => n24161, B2 => n26963, C1 => n23914, C2 => 
                           n26963, A => n3020, ZN => n18856);
   U1573 : AOI22_X1 port map( A1 => DATA1(14), A2 => n27267, B1 => DATA2(14), 
                           B2 => n26964, ZN => n27102);
   U1574 : OAI22_X1 port map( A1 => n26966, A2 => n1789, B1 => n26965, B2 => 
                           n27550, ZN => n26967);
   U1575 : AOI22_X1 port map( A1 => n23608, A2 => n27567, B1 => n26968, B2 => 
                           n26967, ZN => n26970);
   U1576 : NAND3_X1 port map( A1 => DATA2(14), A2 => DATA1(14), A3 => n26981, 
                           ZN => n26969);
   U1577 : OAI211_X1 port map( C1 => n27102, C2 => n27570, A => n26970, B => 
                           n26969, ZN => n18909);
   U1578 : NAND2_X1 port map( A1 => n1831, A2 => n1841, ZN => n19262);
   U1579 : INV_X1 port map( A => n26971, ZN => n26974);
   U1580 : OAI22_X1 port map( A1 => n23633, A2 => n27001, B1 => n24113, B2 => 
                           n26999, ZN => n26972);
   U1581 : AOI211_X1 port map( C1 => n24085, C2 => n26972, A => n23915, B => 
                           n23665, ZN => n26973);
   U1582 : OAI21_X1 port map( B1 => n26974, B2 => n24013, A => n26973, ZN => 
                           OUTALU(14));
   U1583 : OAI22_X1 port map( A1 => n26975, A2 => n27564, B1 => n1820, B2 => 
                           n1896, ZN => n22276);
   U1584 : INV_X1 port map( A => n26976, ZN => n26985);
   U1585 : NOR2_X1 port map( A1 => DATA2(13), A2 => n26977, ZN => n27158);
   U1586 : NAND2_X1 port map( A1 => DATA2(13), A2 => n26977, ZN => n27152);
   U1587 : INV_X1 port map( A => n27152, ZN => n26978);
   U1588 : NOR2_X1 port map( A1 => n27158, A2 => n26978, ZN => n27047);
   U1589 : NOR2_X1 port map( A1 => n27553, A2 => n27552, ZN => n27551);
   U1590 : AOI211_X1 port map( C1 => n26979, C2 => n26994, A => n26987, B => 
                           n27710, ZN => n26980);
   U1591 : AOI22_X1 port map( A1 => n27567, A2 => n23830, B1 => n27551, B2 => 
                           n26980, ZN => n26983);
   U1592 : NAND3_X1 port map( A1 => DATA2(13), A2 => DATA1(13), A3 => n26981, 
                           ZN => n26982);
   U1593 : OAI211_X1 port map( C1 => n27047, C2 => n27570, A => n26983, B => 
                           n26982, ZN => n26984);
   U1594 : AOI221_X1 port map( B1 => n26987, B2 => n26986, C1 => n26985, C2 => 
                           n26986, A => n26984, ZN => n22281);
   U1595 : AOI222_X1 port map( A1 => n26990, A2 => n23887, B1 => n26989, B2 => 
                           n23630, C1 => n26988, C2 => n24061, ZN => n26993);
   U1596 : OAI22_X1 port map( A1 => n24151, A2 => n23743, B1 => n24158, B2 => 
                           n23698, ZN => n26991);
   U1597 : OAI21_X1 port map( B1 => n23664, B2 => n26991, A => n24147, ZN => 
                           n26992);
   U1598 : OAI211_X1 port map( C1 => n24036, C2 => n26993, A => n23913, B => 
                           n26992, ZN => OUTALU(13));
   U1599 : INV_X1 port map( A => n26994, ZN => n26995);
   U1600 : OAI221_X1 port map( B1 => n26996, B2 => n26995, C1 => n27552, C2 => 
                           n26994, A => n27021, ZN => n18855);
   U1601 : OAI222_X1 port map( A1 => n23954, A2 => n23743, B1 => n24156, B2 => 
                           n23698, C1 => n24158, C2 => n24135, ZN => n26997);
   U1602 : AOI22_X1 port map( A1 => n24086, A2 => n26997, B1 => n24160, B2 => 
                           n23942, ZN => n27006);
   U1603 : INV_X1 port map( A => n26998, ZN => n27000);
   U1604 : OAI22_X1 port map( A1 => n24113, A2 => n27000, B1 => n24108, B2 => 
                           n26999, ZN => n27004);
   U1605 : OAI22_X1 port map( A1 => n23633, A2 => n27002, B1 => n23891, B2 => 
                           n27001, ZN => n27003);
   U1606 : OAI21_X1 port map( B1 => n27004, B2 => n27003, A => n24085, ZN => 
                           n27005);
   U1607 : NAND4_X1 port map( A1 => n23607, A2 => n23637, A3 => n27006, A4 => 
                           n27005, ZN => OUTALU(12));
   U1608 : INV_X1 port map( A => n27008, ZN => n27007);
   U1609 : AOI221_X1 port map( B1 => n27009, B2 => n27008, C1 => n27011, C2 => 
                           n27007, A => n1789, ZN => n18854);
   U1610 : INV_X1 port map( A => n27010, ZN => n27012);
   U1611 : AOI21_X1 port map( B1 => n27012, B2 => n27011, A => n27550, ZN => 
                           n19165);
   U1612 : OAI22_X1 port map( A1 => n24156, A2 => n24135, B1 => n23742, B2 => 
                           n24157, ZN => n27013);
   U1613 : AOI211_X1 port map( C1 => n24086, C2 => n27013, A => n23606, B => 
                           n24120, ZN => n27015);
   U1614 : AOI22_X1 port map( A1 => n23912, A2 => n24014, B1 => n24033, B2 => 
                           n27029, ZN => n27014);
   U1615 : NAND2_X1 port map( A1 => n27015, A2 => n27014, ZN => OUTALU(11));
   U1616 : OAI21_X1 port map( B1 => n27023, B2 => n27017, A => n27016, ZN => 
                           n27026);
   U1617 : OAI21_X1 port map( B1 => n27270, B2 => n27033, A => n27018, ZN => 
                           n27019);
   U1618 : AOI22_X1 port map( A1 => DATA1(10), A2 => n27270, B1 => DATA2(10), 
                           B2 => n27151, ZN => n27098);
   U1619 : INV_X1 port map( A => n27098, ZN => n27145);
   U1620 : AOI22_X1 port map( A1 => DATA1(10), A2 => n27019, B1 => n27557, B2 
                           => n27145, ZN => n27025);
   U1621 : OAI211_X1 port map( C1 => n27023, C2 => n27022, A => n27021, B => 
                           n27020, ZN => n27024);
   U1622 : OAI211_X1 port map( C1 => n27550, C2 => n27026, A => n27025, B => 
                           n27024, ZN => n27027);
   U1623 : AOI21_X1 port map( B1 => n22313, B2 => n23613, A => n27027, ZN => 
                           n19164);
   U1624 : AOI22_X1 port map( A1 => n24092, A2 => n27029, B1 => n23962, B2 => 
                           n27028, ZN => n27031);
   U1625 : OR3_X1 port map( A1 => n24156, A2 => n23743, A3 => n24029, ZN => 
                           n27030);
   U1626 : OAI211_X1 port map( C1 => n24036, C2 => n27031, A => n23663, B => 
                           n27030, ZN => OUTALU(10));
   U1627 : OAI21_X1 port map( B1 => n27573, B2 => n27033, A => n27032, ZN => 
                           n27038);
   U1628 : NAND2_X1 port map( A1 => n24173, A2 => n27573, ZN => n27079);
   U1629 : NAND2_X1 port map( A1 => DATA2(0), A2 => n24053, ZN => n27128);
   U1630 : AND2_X1 port map( A1 => n27079, A2 => n27128, ZN => n27054);
   U1631 : NOR2_X1 port map( A1 => n27035, A2 => n27034, ZN => n27039);
   U1632 : OAI22_X1 port map( A1 => n27054, A2 => n27570, B1 => n27039, B2 => 
                           n27036, ZN => n27037);
   U1633 : AOI21_X1 port map( B1 => n24173, B2 => n27038, A => n27037, ZN => 
                           n18848);
   U1634 : AOI22_X1 port map( A1 => n27567, A2 => n24005, B1 => n27040, B2 => 
                           n27039, ZN => n18904);
   U1635 : NOR2_X1 port map( A1 => n27042, A2 => n27041, ZN => n8626);
   U1636 : NAND2_X1 port map( A1 => FUNC(3), A2 => n8626, ZN => n19259);
   U1637 : AOI21_X1 port map( B1 => n24047, B2 => DATA2(7), A => n27043, ZN => 
                           n27092);
   U1638 : NAND4_X1 port map( A1 => n27047, A2 => n27046, A3 => n27045, A4 => 
                           n27044, ZN => n27048);
   U1639 : NOR4_X1 port map( A1 => n27150, A2 => n27082, A3 => n27049, A4 => 
                           n27048, ZN => n27050);
   U1640 : INV_X1 port map( A => n27139, ZN => n27089);
   U1641 : NAND4_X1 port map( A1 => n27092, A2 => n27050, A3 => n27130, A4 => 
                           n27089, ZN => n27076);
   U1642 : INV_X1 port map( A => DATA2(12), ZN => n27548);
   U1643 : NOR2_X1 port map( A1 => DATA1(12), A2 => n27548, ZN => n27099);
   U1644 : INV_X1 port map( A => n27099, ZN => n27153);
   U1645 : OAI21_X1 port map( B1 => n27547, B2 => DATA2(12), A => n27153, ZN =>
                           n27556);
   U1646 : OR2_X1 port map( A1 => n27556, A2 => n27096, ZN => n27154);
   U1647 : INV_X1 port map( A => DATA2(21), ZN => n27260);
   U1648 : NAND2_X1 port map( A1 => DATA1(21), A2 => n27260, ZN => n27124);
   U1649 : NOR2_X1 port map( A1 => DATA1(21), A2 => n27260, ZN => n27565);
   U1650 : INV_X1 port map( A => n27565, ZN => n27174);
   U1651 : INV_X1 port map( A => DATA2(6), ZN => n27534);
   U1652 : OAI22_X1 port map( A1 => n27534, A2 => n24178, B1 => n24077, B2 => 
                           DATA2(6), ZN => n27051);
   U1653 : INV_X1 port map( A => n27051, ZN => n27533);
   U1654 : NAND3_X1 port map( A1 => n27124, A2 => n27174, A3 => n27533, ZN => 
                           n27052);
   U1655 : NOR4_X1 port map( A1 => n27127, A2 => n27145, A3 => n27154, A4 => 
                           n27052, ZN => n27073);
   U1656 : NAND4_X1 port map( A1 => n27056, A2 => n27055, A3 => n27054, A4 => 
                           n27053, ZN => n27071);
   U1657 : NAND4_X1 port map( A1 => n27102, A2 => n27057, A3 => n27192, A4 => 
                           n27120, ZN => n27070);
   U1658 : INV_X1 port map( A => n27058, ZN => n27063);
   U1659 : INV_X1 port map( A => n27059, ZN => n27061);
   U1660 : NAND4_X1 port map( A1 => n27063, A2 => n27062, A3 => n27061, A4 => 
                           n27060, ZN => n27069);
   U1661 : NAND4_X1 port map( A1 => n27067, A2 => n27066, A3 => n27065, A4 => 
                           n27064, ZN => n27068);
   U1662 : NOR4_X1 port map( A1 => n27071, A2 => n27070, A3 => n27069, A4 => 
                           n27068, ZN => n27072);
   U1663 : NAND4_X1 port map( A1 => n27074, A2 => n27179, A3 => n27073, A4 => 
                           n27072, ZN => n27075);
   U1664 : OAI21_X1 port map( B1 => n27076, B2 => n27075, A => n1832, ZN => 
                           n27078);
   U1665 : AOI211_X1 port map( C1 => FUNC(2), C2 => n27078, A => FUNC(1), B => 
                           n27077, ZN => n18903);
   U1666 : NOR2_X1 port map( A1 => DATA2(24), A2 => n27185, ZN => n27116);
   U1667 : AOI22_X1 port map( A1 => DATA1(15), A2 => n27266, B1 => DATA1(14), 
                           B2 => n27267, ZN => n27160);
   U1668 : NAND2_X1 port map( A1 => DATA1(12), A2 => n27548, ZN => n27101);
   U1669 : NAND2_X1 port map( A1 => n27137, A2 => n27130, ZN => n27084);
   U1670 : AOI211_X1 port map( C1 => n27080, C2 => n27079, A => n27127, B => 
                           n27125, ZN => n27081);
   U1671 : AOI211_X1 port map( C1 => n24049, C2 => n27592, A => n27082, B => 
                           n27081, ZN => n27083);
   U1672 : OAI21_X1 port map( B1 => n27084, B2 => n27083, A => n27131, ZN => 
                           n27086);
   U1673 : INV_X1 port map( A => n27085, ZN => n27136);
   U1674 : OAI211_X1 port map( C1 => n27087, C2 => n27086, A => n27533, B => 
                           n27136, ZN => n27088);
   U1675 : OAI211_X1 port map( C1 => DATA2(6), C2 => n24055, A => n27089, B => 
                           n27088, ZN => n27091);
   U1676 : INV_X1 port map( A => n27090, ZN => n27140);
   U1677 : AOI21_X1 port map( B1 => n27092, B2 => n27091, A => n27140, ZN => 
                           n27094);
   U1678 : OAI21_X1 port map( B1 => n27144, B2 => n27094, A => n27093, ZN => 
                           n27097);
   U1679 : NOR2_X1 port map( A1 => DATA2(10), A2 => n27151, ZN => n27095);
   U1680 : AOI211_X1 port map( C1 => n27098, C2 => n27097, A => n27096, B => 
                           n27095, ZN => n27100);
   U1681 : AOI221_X1 port map( B1 => n27150, B2 => n27101, C1 => n27100, C2 => 
                           n27101, A => n27099, ZN => n27103);
   U1682 : OAI211_X1 port map( C1 => n27158, C2 => n27103, A => n27102, B => 
                           n27152, ZN => n27104);
   U1683 : OAI22_X1 port map( A1 => DATA1(15), A2 => n27266, B1 => DATA1(16), 
                           B2 => n27265, ZN => n27161);
   U1684 : AOI21_X1 port map( B1 => n27160, B2 => n27104, A => n27161, ZN => 
                           n27106);
   U1685 : AOI221_X1 port map( B1 => n27107, B2 => n27165, C1 => n27106, C2 => 
                           n27165, A => n27105, ZN => n27108);
   U1686 : OAI21_X1 port map( B1 => n27167, B2 => n27108, A => n27172, ZN => 
                           n27110);
   U1687 : OAI211_X1 port map( C1 => n27163, C2 => n27110, A => n27109, B => 
                           n27176, ZN => n27111);
   U1688 : OAI221_X1 port map( B1 => n27565, B2 => n27173, C1 => n27565, C2 => 
                           n27111, A => n27124, ZN => n27113);
   U1689 : NOR2_X1 port map( A1 => DATA2(22), A2 => n27177, ZN => n27112);
   U1690 : AOI211_X1 port map( C1 => n27179, C2 => n27113, A => n27112, B => 
                           n27181, ZN => n27114);
   U1691 : AOI211_X1 port map( C1 => DATA2(23), C2 => n1840, A => n27114, B => 
                           n27180, ZN => n27115);
   U1692 : AOI221_X1 port map( B1 => n27116, B2 => n27188, C1 => n27115, C2 => 
                           n27188, A => n27187, ZN => n27117);
   U1693 : OAI22_X1 port map( A1 => DATA2(26), A2 => n27191, B1 => n27117, B2 
                           => n27186, ZN => n27118);
   U1694 : OAI211_X1 port map( C1 => n27194, C2 => n27118, A => n27192, B => 
                           n27195, ZN => n27119);
   U1695 : OAI21_X1 port map( B1 => DATA2(28), B2 => n27198, A => n27119, ZN =>
                           n27121);
   U1696 : OAI211_X1 port map( C1 => n27200, C2 => n27121, A => n27120, B => 
                           n27201, ZN => n27123);
   U1697 : OAI211_X1 port map( C1 => DATA2(30), C2 => n27205, A => n27123, B =>
                           n27122, ZN => n27209);
   U1698 : INV_X1 port map( A => n27124, ZN => n27566);
   U1699 : AOI22_X1 port map( A1 => DATA2(6), A2 => n24055, B1 => n24047, B2 =>
                           DATA2(7), ZN => n27142);
   U1700 : INV_X1 port map( A => n27125, ZN => n27129);
   U1701 : AOI211_X1 port map( C1 => n27129, C2 => n27128, A => n27127, B => 
                           n27126, ZN => n27134);
   U1702 : OAI21_X1 port map( B1 => n24049, B2 => n27592, A => n27130, ZN => 
                           n27133);
   U1703 : OAI211_X1 port map( C1 => n27134, C2 => n27133, A => n27132, B => 
                           n27131, ZN => n27135);
   U1704 : NAND3_X1 port map( A1 => n27137, A2 => n27136, A3 => n27135, ZN => 
                           n27138);
   U1705 : OAI211_X1 port map( C1 => n24056, C2 => DATA2(5), A => n27533, B => 
                           n27138, ZN => n27141);
   U1706 : AOI211_X1 port map( C1 => n27142, C2 => n27141, A => n27140, B => 
                           n27139, ZN => n27143);
   U1707 : AOI21_X1 port map( B1 => DATA2(8), B2 => n24046, A => n27143, ZN => 
                           n27148);
   U1708 : INV_X1 port map( A => n27144, ZN => n27147);
   U1709 : AOI211_X1 port map( C1 => n27148, C2 => n27147, A => n27146, B => 
                           n27145, ZN => n27149);
   U1710 : AOI211_X1 port map( C1 => DATA2(10), C2 => n27151, A => n27150, B =>
                           n27149, ZN => n27155);
   U1711 : OAI211_X1 port map( C1 => n27155, C2 => n27154, A => n27153, B => 
                           n27152, ZN => n27156);
   U1712 : INV_X1 port map( A => n27156, ZN => n27157);
   U1713 : OAI22_X1 port map( A1 => n27267, A2 => DATA1(14), B1 => n27158, B2 
                           => n27157, ZN => n27162);
   U1714 : OAI221_X1 port map( B1 => n27162, B2 => n27161, C1 => n27160, C2 => 
                           n27161, A => n27159, ZN => n27164);
   U1715 : AOI21_X1 port map( B1 => n27165, B2 => n27164, A => n27163, ZN => 
                           n27168);
   U1716 : AOI211_X1 port map( C1 => n27169, C2 => n27168, A => n27167, B => 
                           n27166, ZN => n27170);
   U1717 : INV_X1 port map( A => n27170, ZN => n27171);
   U1718 : NAND3_X1 port map( A1 => n27173, A2 => n27172, A3 => n27171, ZN => 
                           n27175);
   U1719 : OAI221_X1 port map( B1 => n27566, B2 => n27176, C1 => n27566, C2 => 
                           n27175, A => n27174, ZN => n27178);
   U1720 : AOI22_X1 port map( A1 => n27179, A2 => n27178, B1 => DATA2(22), B2 
                           => n27177, ZN => n27183);
   U1721 : AOI211_X1 port map( C1 => n27183, C2 => n27182, A => n27181, B => 
                           n27180, ZN => n27184);
   U1722 : AOI21_X1 port map( B1 => DATA2(24), B2 => n27185, A => n27184, ZN =>
                           n27189);
   U1723 : AOI211_X1 port map( C1 => n27189, C2 => n27188, A => n27187, B => 
                           n27186, ZN => n27190);
   U1724 : AOI21_X1 port map( B1 => DATA2(26), B2 => n27191, A => n27190, ZN =>
                           n27196);
   U1725 : INV_X1 port map( A => n27192, ZN => n27193);
   U1726 : AOI211_X1 port map( C1 => n27196, C2 => n27195, A => n27194, B => 
                           n27193, ZN => n27197);
   U1727 : AOI21_X1 port map( B1 => DATA2(28), B2 => n27198, A => n27197, ZN =>
                           n27202);
   U1728 : AOI211_X1 port map( C1 => n27202, C2 => n27201, A => n27200, B => 
                           n27199, ZN => n27203);
   U1729 : AOI211_X1 port map( C1 => DATA2(30), C2 => n27205, A => n27204, B =>
                           n27203, ZN => n27206);
   U1730 : AOI221_X1 port map( B1 => n27207, B2 => n1832, C1 => n27206, C2 => 
                           n1832, A => FUNC(2), ZN => n27208);
   U1731 : OAI221_X1 port map( B1 => n1832, B2 => n27210, C1 => n1832, C2 => 
                           n27209, A => n27208, ZN => n18853);
   U1732 : INV_X1 port map( A => n27211, ZN => n27244);
   U1733 : OAI22_X1 port map( A1 => n23893, A2 => n27213, B1 => n27212, B2 => 
                           n24068, ZN => n27243);
   U1734 : AOI22_X1 port map( A1 => n24082, A2 => n27215, B1 => n23631, B2 => 
                           n27214, ZN => n27235);
   U1735 : INV_X1 port map( A => n27216, ZN => n27233);
   U1736 : INV_X1 port map( A => n27217, ZN => n27219);
   U1737 : AOI22_X1 port map( A1 => n24123, A2 => n27219, B1 => n23630, B2 => 
                           n27218, ZN => n27230);
   U1738 : NAND2_X1 port map( A1 => n23660, A2 => n24101, ZN => n27220);
   U1739 : OAI21_X1 port map( B1 => n24158, B2 => n23674, A => n27220, ZN => 
                           n27222);
   U1740 : OAI22_X1 port map( A1 => n23954, A2 => n23687, B1 => n23957, B2 => 
                           n24140, ZN => n27221);
   U1741 : AOI211_X1 port map( C1 => n27668, C2 => n27223, A => n27222, B => 
                           n27221, ZN => n27224);
   U1742 : OAI222_X1 port map( A1 => n23979, A2 => n27226, B1 => n24080, B2 => 
                           n27225, C1 => n24105, C2 => n27224, ZN => n27228);
   U1743 : AOI22_X1 port map( A1 => n23887, A2 => n27228, B1 => n23964, B2 => 
                           n27227, ZN => n27229);
   U1744 : OAI211_X1 port map( C1 => n23891, C2 => n27231, A => n27230, B => 
                           n27229, ZN => n27232);
   U1745 : AOI22_X1 port map( A1 => n24093, A2 => n27233, B1 => n23962, B2 => 
                           n27232, ZN => n27234);
   U1746 : OAI211_X1 port map( C1 => n23894, C2 => n27236, A => n27235, B => 
                           n27234, ZN => n27237);
   U1747 : AOI222_X1 port map( A1 => n27239, A2 => n23975, B1 => n27238, B2 => 
                           n23971, C1 => n27237, C2 => n24083, ZN => n27240);
   U1748 : OAI22_X1 port map( A1 => n23977, A2 => n27241, B1 => n24111, B2 => 
                           n27240, ZN => n27242);
   U1749 : AOI211_X1 port map( C1 => n23892, C2 => n27244, A => n27243, B => 
                           n27242, ZN => n27245);
   U1750 : OAI211_X1 port map( C1 => n24036, C2 => n27245, A => n23599, B => 
                           n23662, ZN => n27246);
   U1751 : AOI21_X1 port map( B1 => n23605, B2 => n23661, A => n27246, ZN => 
                           n27247);
   U1752 : OAI21_X1 port map( B1 => n24011, B2 => n27248, A => n27247, ZN => 
                           OUTALU(0));
   U1753 : NAND2_X1 port map( A1 => n27249, A2 => n1832, ZN => n27278);
   U1754 : CLKBUF_X1 port map( A => n27278, Z => n27274);
   U1755 : NAND2_X1 port map( A1 => FUNC(3), A2 => n27249, ZN => n27277);
   U1756 : CLKBUF_X1 port map( A => n27277, Z => n27273);
   U1757 : AOI22_X1 port map( A1 => DATA2(31), A2 => n27274, B1 => n27273, B2 
                           => n27250, ZN => N2548);
   U1758 : AOI22_X1 port map( A1 => DATA2(30), A2 => n27278, B1 => n27277, B2 
                           => n27251, ZN => N2547);
   U1759 : INV_X1 port map( A => DATA2(29), ZN => n27252);
   U1760 : AOI22_X1 port map( A1 => DATA2(29), A2 => n27274, B1 => n27273, B2 
                           => n27252, ZN => N2546);
   U1761 : AOI22_X1 port map( A1 => DATA2(28), A2 => n27278, B1 => n27277, B2 
                           => n27253, ZN => N2545);
   U1762 : INV_X1 port map( A => DATA2(27), ZN => n27254);
   U1763 : AOI22_X1 port map( A1 => DATA2(27), A2 => n27274, B1 => n27273, B2 
                           => n27254, ZN => N2544);
   U1764 : AOI22_X1 port map( A1 => DATA2(26), A2 => n27278, B1 => n27277, B2 
                           => n27255, ZN => N2543);
   U1765 : INV_X1 port map( A => DATA2(25), ZN => n27256);
   U1766 : AOI22_X1 port map( A1 => DATA2(25), A2 => n27274, B1 => n27273, B2 
                           => n27256, ZN => N2542);
   U1767 : AOI22_X1 port map( A1 => DATA2(24), A2 => n27278, B1 => n27277, B2 
                           => n27257, ZN => N2541);
   U1768 : INV_X1 port map( A => DATA2(23), ZN => n27258);
   U1769 : AOI22_X1 port map( A1 => DATA2(23), A2 => n27274, B1 => n27273, B2 
                           => n27258, ZN => N2540);
   U1770 : AOI22_X1 port map( A1 => DATA2(22), A2 => n27278, B1 => n27277, B2 
                           => n27259, ZN => N2539);
   U1771 : AOI22_X1 port map( A1 => DATA2(21), A2 => n27278, B1 => n27277, B2 
                           => n27260, ZN => N2538);
   U1772 : AOI22_X1 port map( A1 => DATA2(20), A2 => n27278, B1 => n27277, B2 
                           => n27261, ZN => N2537);
   U1773 : AOI22_X1 port map( A1 => DATA2(19), A2 => n27274, B1 => n27273, B2 
                           => n27262, ZN => N2536);
   U1774 : AOI22_X1 port map( A1 => DATA2(18), A2 => n27274, B1 => n27273, B2 
                           => n27263, ZN => N2535);
   U1775 : INV_X1 port map( A => DATA2(17), ZN => n27264);
   U1776 : AOI22_X1 port map( A1 => DATA2(17), A2 => n27274, B1 => n27273, B2 
                           => n27264, ZN => N2534);
   U1777 : AOI22_X1 port map( A1 => DATA2(16), A2 => n27274, B1 => n27273, B2 
                           => n27265, ZN => N2533);
   U1778 : AOI22_X1 port map( A1 => DATA2(15), A2 => n27274, B1 => n27273, B2 
                           => n27266, ZN => N2532);
   U1779 : AOI22_X1 port map( A1 => DATA2(14), A2 => n27274, B1 => n27273, B2 
                           => n27267, ZN => N2531);
   U1780 : INV_X1 port map( A => DATA2(13), ZN => n27268);
   U1781 : AOI22_X1 port map( A1 => DATA2(13), A2 => n27274, B1 => n27273, B2 
                           => n27268, ZN => N2530);
   U1782 : AOI22_X1 port map( A1 => DATA2(12), A2 => n27274, B1 => n27273, B2 
                           => n27548, ZN => N2529);
   U1783 : AOI22_X1 port map( A1 => DATA2(11), A2 => n27274, B1 => n27273, B2 
                           => n27269, ZN => N2528);
   U1784 : AOI22_X1 port map( A1 => DATA2(10), A2 => n27274, B1 => n27273, B2 
                           => n27270, ZN => N2527);
   U1785 : AOI22_X1 port map( A1 => DATA2(9), A2 => n27274, B1 => n27273, B2 =>
                           n27271, ZN => N2526);
   U1786 : AOI22_X1 port map( A1 => DATA2(8), A2 => n27274, B1 => n27273, B2 =>
                           n27272, ZN => N2525);
   U1787 : INV_X1 port map( A => DATA2(7), ZN => n27275);
   U1788 : AOI22_X1 port map( A1 => DATA2(7), A2 => n27278, B1 => n27277, B2 =>
                           n27275, ZN => N2524);
   U1789 : AOI22_X1 port map( A1 => DATA2(6), A2 => n27278, B1 => n27277, B2 =>
                           n27534, ZN => N2523);
   U1790 : AOI22_X1 port map( A1 => DATA2(5), A2 => n27278, B1 => n27277, B2 =>
                           n27276, ZN => N2522);
   U1791 : AOI22_X1 port map( A1 => DATA2(4), A2 => n27278, B1 => n27277, B2 =>
                           n27577, ZN => N2521);
   U1792 : AOI22_X1 port map( A1 => DATA2(3), A2 => n27278, B1 => n27277, B2 =>
                           n27594, ZN => N2520);
   U1793 : AOI22_X1 port map( A1 => DATA2(2), A2 => n27278, B1 => n27277, B2 =>
                           n27592, ZN => N2519);
   U1794 : AOI22_X1 port map( A1 => DATA2(1), A2 => n27278, B1 => n27277, B2 =>
                           n27571, ZN => N2518);
   U1795 : AOI22_X1 port map( A1 => DATA2(0), A2 => n27278, B1 => n27277, B2 =>
                           n27573, ZN => N2517);
   U1796 : NOR2_X1 port map( A1 => n27279, A2 => n1807, ZN => n19253);
   U1797 : NAND2_X1 port map( A1 => n27318, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n27283);
   U1798 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , ZN => n27314);
   U1799 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n27314, ZN => n27313);
   U1800 : INV_X1 port map( A => n27280, ZN => n27281);
   U1801 : AOI22_X1 port map( A1 => n25900, A2 => n27316, B1 => n9084, B2 => 
                           n27310, ZN => n27282);
   U1802 : OAI221_X1 port map( B1 => n1807, B2 => n27283, C1 => n1807, C2 => 
                           n27313, A => n27282, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1803 : INV_X1 port map( A => n27283, ZN => n27315);
   U1804 : AOI22_X1 port map( A1 => n25898, A2 => n27316, B1 => n25900, B2 => 
                           n27315, ZN => n27285);
   U1805 : NAND2_X1 port map( A1 => n9081, A2 => n27310, ZN => n27284);
   U1806 : OAI211_X1 port map( C1 => n1805, C2 => n27313, A => n27285, B => 
                           n27284, ZN => boothmul_pipelined_i_mux_out_1_4_port)
                           ;
   U1807 : AOI22_X1 port map( A1 => n25898, A2 => n27315, B1 => n27316, B2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n27287);
   U1808 : NAND2_X1 port map( A1 => n27310, A2 => n9078, ZN => n27286);
   U1809 : OAI211_X1 port map( C1 => n27313, C2 => n1804, A => n27287, B => 
                           n27286, ZN => boothmul_pipelined_i_mux_out_1_5_port)
                           ;
   U1810 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n27289);
   U1811 : NAND2_X1 port map( A1 => n27310, A2 => n9075, ZN => n27288);
   U1812 : OAI211_X1 port map( C1 => n1803, C2 => n27313, A => n27289, B => 
                           n27288, ZN => boothmul_pipelined_i_mux_out_1_6_port)
                           ;
   U1813 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n27291);
   U1814 : NAND2_X1 port map( A1 => n27310, A2 => n9072, ZN => n27290);
   U1815 : OAI211_X1 port map( C1 => n1802, C2 => n27313, A => n27291, B => 
                           n27290, ZN => boothmul_pipelined_i_mux_out_1_7_port)
                           ;
   U1816 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n27293);
   U1817 : NAND2_X1 port map( A1 => n27310, A2 => n9069, ZN => n27292);
   U1818 : OAI211_X1 port map( C1 => n1800, C2 => n27313, A => n27293, B => 
                           n27292, ZN => boothmul_pipelined_i_mux_out_1_8_port)
                           ;
   U1819 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n27295);
   U1820 : NAND2_X1 port map( A1 => n27310, A2 => n9066, ZN => n27294);
   U1821 : OAI211_X1 port map( C1 => n1799, C2 => n27313, A => n27295, B => 
                           n27294, ZN => boothmul_pipelined_i_mux_out_1_9_port)
                           ;
   U1822 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n27297);
   U1823 : NAND2_X1 port map( A1 => n27310, A2 => n9063, ZN => n27296);
   U1824 : OAI211_X1 port map( C1 => n1798, C2 => n27313, A => n27297, B => 
                           n27296, ZN => boothmul_pipelined_i_mux_out_1_10_port
                           );
   U1825 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n27299);
   U1826 : NAND2_X1 port map( A1 => n27310, A2 => n9060, ZN => n27298);
   U1827 : OAI211_X1 port map( C1 => n1797, C2 => n27313, A => n27299, B => 
                           n27298, ZN => boothmul_pipelined_i_mux_out_1_11_port
                           );
   U1828 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n27301);
   U1829 : NAND2_X1 port map( A1 => n27310, A2 => n9057, ZN => n27300);
   U1830 : OAI211_X1 port map( C1 => n1796, C2 => n27313, A => n27301, B => 
                           n27300, ZN => boothmul_pipelined_i_mux_out_1_12_port
                           );
   U1831 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n27303);
   U1832 : NAND2_X1 port map( A1 => n27310, A2 => n9054, ZN => n27302);
   U1833 : OAI211_X1 port map( C1 => n1795, C2 => n27313, A => n27303, B => 
                           n27302, ZN => boothmul_pipelined_i_mux_out_1_13_port
                           );
   U1834 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n27305);
   U1835 : NAND2_X1 port map( A1 => n27310, A2 => n9051, ZN => n27304);
   U1836 : OAI211_X1 port map( C1 => n1794, C2 => n27313, A => n27305, B => 
                           n27304, ZN => boothmul_pipelined_i_mux_out_1_14_port
                           );
   U1837 : AOI22_X1 port map( A1 => n27316, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n27307);
   U1838 : NAND2_X1 port map( A1 => n27310, A2 => n9048, ZN => n27306);
   U1839 : OAI211_X1 port map( C1 => n1793, C2 => n27313, A => n27307, B => 
                           n27306, ZN => boothmul_pipelined_i_mux_out_1_15_port
                           );
   U1840 : AOI22_X1 port map( A1 => n27316, A2 => n25894, B1 => n27315, B2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n27309);
   U1841 : NAND2_X1 port map( A1 => n27310, A2 => n9045, ZN => n27308);
   U1842 : OAI211_X1 port map( C1 => n1792, C2 => n27313, A => n27309, B => 
                           n27308, ZN => boothmul_pipelined_i_mux_out_1_16_port
                           );
   U1843 : AOI22_X1 port map( A1 => n27316, A2 => n25896, B1 => n27315, B2 => 
                           n25894, ZN => n27312);
   U1844 : NAND2_X1 port map( A1 => n27310, A2 => data1_mul_15_port, ZN => 
                           n27311);
   U1845 : OAI211_X1 port map( C1 => n1791, C2 => n27313, A => n27312, B => 
                           n27311, ZN => boothmul_pipelined_i_mux_out_1_17_port
                           );
   U1846 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n27314, ZN => 
                           n27319);
   U1847 : XOR2_X1 port map( A => data1_mul_15_port, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => n27443);
   U1848 : INV_X1 port map( A => n27443, ZN => n27527);
   U1849 : AOI22_X1 port map( A1 => n27316, A2 => n27527, B1 => n27315, B2 => 
                           n25896, ZN => n27317);
   U1850 : OAI21_X1 port map( B1 => n27319, B2 => n27318, A => n27317, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1851 : OR2_X1 port map( A1 => n27320, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n19252);
   U1852 : AOI22_X1 port map( A1 => n25900, A2 => n23972, B1 => n9084, B2 => 
                           n23949, ZN => n27321);
   U1853 : OAI221_X1 port map( B1 => n1807, B2 => n23974, C1 => n1807, C2 => 
                           n24004, A => n27321, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1854 : AOI22_X1 port map( A1 => n25900, A2 => n24109, B1 => n9081, B2 => 
                           n23949, ZN => n27323);
   U1855 : NAND2_X1 port map( A1 => n25898, A2 => n23972, ZN => n27322);
   U1856 : OAI211_X1 port map( C1 => n24004, C2 => n1805, A => n27323, B => 
                           n27322, ZN => boothmul_pipelined_i_mux_out_2_6_port)
                           ;
   U1857 : AOI22_X1 port map( A1 => n9078, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n23972, ZN => n27325);
   U1858 : NAND2_X1 port map( A1 => n25898, A2 => n24109, ZN => n27324);
   U1859 : OAI211_X1 port map( C1 => n24004, C2 => n1804, A => n27325, B => 
                           n27324, ZN => boothmul_pipelined_i_mux_out_2_7_port)
                           ;
   U1860 : AOI22_X1 port map( A1 => n9075, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n23972, ZN => n27327);
   U1861 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n24109, ZN => n27326);
   U1862 : OAI211_X1 port map( C1 => n24004, C2 => n1803, A => n27327, B => 
                           n27326, ZN => boothmul_pipelined_i_mux_out_2_8_port)
                           ;
   U1863 : AOI22_X1 port map( A1 => n9072, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n23972, ZN => n27329);
   U1864 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n24109, ZN => n27328);
   U1865 : OAI211_X1 port map( C1 => n24004, C2 => n1802, A => n27329, B => 
                           n27328, ZN => boothmul_pipelined_i_mux_out_2_9_port)
                           ;
   U1866 : AOI22_X1 port map( A1 => n9069, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n23972, ZN => n27331);
   U1867 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n24109, ZN => n27330);
   U1868 : OAI211_X1 port map( C1 => n24004, C2 => n1800, A => n27331, B => 
                           n27330, ZN => boothmul_pipelined_i_mux_out_2_10_port
                           );
   U1869 : AOI22_X1 port map( A1 => n9066, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n23972, ZN => n27333);
   U1870 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n24109, ZN => n27332);
   U1871 : OAI211_X1 port map( C1 => n24004, C2 => n1799, A => n27333, B => 
                           n27332, ZN => boothmul_pipelined_i_mux_out_2_11_port
                           );
   U1872 : AOI22_X1 port map( A1 => n9063, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n23972, ZN => n27335);
   U1873 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n24109, ZN => n27334);
   U1874 : OAI211_X1 port map( C1 => n24004, C2 => n1798, A => n27335, B => 
                           n27334, ZN => boothmul_pipelined_i_mux_out_2_12_port
                           );
   U1875 : AOI22_X1 port map( A1 => n9060, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n23972, ZN => n27337);
   U1876 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n24109, ZN => n27336);
   U1877 : OAI211_X1 port map( C1 => n24004, C2 => n1797, A => n27337, B => 
                           n27336, ZN => boothmul_pipelined_i_mux_out_2_13_port
                           );
   U1878 : AOI22_X1 port map( A1 => n9057, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n23972, ZN => n27339);
   U1879 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n24109, ZN => n27338);
   U1880 : OAI211_X1 port map( C1 => n24004, C2 => n1796, A => n27339, B => 
                           n27338, ZN => boothmul_pipelined_i_mux_out_2_14_port
                           );
   U1881 : AOI22_X1 port map( A1 => n9054, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n23972, ZN => n27341);
   U1882 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n24109, ZN => n27340);
   U1883 : OAI211_X1 port map( C1 => n24004, C2 => n1795, A => n27341, B => 
                           n27340, ZN => boothmul_pipelined_i_mux_out_2_15_port
                           );
   U1884 : AOI22_X1 port map( A1 => n9051, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n23972, ZN => n27343);
   U1885 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n24109, ZN => n27342);
   U1886 : OAI211_X1 port map( C1 => n24004, C2 => n1794, A => n27343, B => 
                           n27342, ZN => boothmul_pipelined_i_mux_out_2_16_port
                           );
   U1887 : AOI22_X1 port map( A1 => n9048, A2 => n23949, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n23972, ZN => n27345);
   U1888 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n24109, ZN => n27344);
   U1889 : OAI211_X1 port map( C1 => n24004, C2 => n1793, A => n27345, B => 
                           n27344, ZN => boothmul_pipelined_i_mux_out_2_17_port
                           );
   U1890 : AOI22_X1 port map( A1 => n9045, A2 => n23949, B1 => n25894, B2 => 
                           n23972, ZN => n27347);
   U1891 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n24109, ZN => n27346);
   U1892 : OAI211_X1 port map( C1 => n24004, C2 => n1792, A => n27347, B => 
                           n27346, ZN => boothmul_pipelined_i_mux_out_2_18_port
                           );
   U1893 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n23949, B1 => 
                           n25896, B2 => n23972, ZN => n27349);
   U1894 : NAND2_X1 port map( A1 => n25894, A2 => n24109, ZN => n27348);
   U1895 : OAI211_X1 port map( C1 => n24004, C2 => n1791, A => n27349, B => 
                           n27348, ZN => boothmul_pipelined_i_mux_out_2_19_port
                           );
   U1896 : OAI222_X1 port map( A1 => n25895, A2 => n23974, B1 => n1790, B2 => 
                           n23950, C1 => n24079, C2 => n27443, ZN => n18847);
   U1897 : NAND2_X1 port map( A1 => n7769, A2 => n27350, ZN => n19251);
   U1898 : AOI22_X1 port map( A1 => n25900, A2 => n24130, B1 => n9084, B2 => 
                           n24087, ZN => n27351);
   U1899 : OAI221_X1 port map( B1 => n1807, B2 => n24003, C1 => n1807, C2 => 
                           n24129, A => n27351, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1900 : OAI22_X1 port map( A1 => n24003, A2 => n25899, B1 => n24129, B2 => 
                           n1805, ZN => n27352);
   U1901 : AOI21_X1 port map( B1 => n25898, B2 => n24130, A => n27352, ZN => 
                           n27353);
   U1902 : OAI21_X1 port map( B1 => n24169, B2 => n1804, A => n27353, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1903 : OAI22_X1 port map( A1 => n24129, A2 => n1804, B1 => n24169, B2 => 
                           n1803, ZN => n27354);
   U1904 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           B2 => n24130, A => n27354, ZN => n27355);
   U1905 : OAI21_X1 port map( B1 => n24003, B2 => n25897, A => n27355, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1906 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN 
                           => n27512);
   U1907 : OAI22_X1 port map( A1 => n24003, A2 => n27512, B1 => n24169, B2 => 
                           n1802, ZN => n27356);
   U1908 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           B2 => n24130, A => n27356, ZN => n27357);
   U1909 : OAI21_X1 port map( B1 => n24129, B2 => n1803, A => n27357, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1910 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN 
                           => n27513);
   U1911 : OAI22_X1 port map( A1 => n24003, A2 => n27513, B1 => n24169, B2 => 
                           n1800, ZN => n27358);
   U1912 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           B2 => n24130, A => n27358, ZN => n27359);
   U1913 : OAI21_X1 port map( B1 => n24129, B2 => n1802, A => n27359, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1914 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN 
                           => n27514);
   U1915 : OAI22_X1 port map( A1 => n24003, A2 => n27514, B1 => n24169, B2 => 
                           n1799, ZN => n27360);
   U1916 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           B2 => n24130, A => n27360, ZN => n27361);
   U1917 : OAI21_X1 port map( B1 => n24129, B2 => n1800, A => n27361, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1918 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN 
                           => n27515);
   U1919 : OAI22_X1 port map( A1 => n24003, A2 => n27515, B1 => n24169, B2 => 
                           n1798, ZN => n27362);
   U1920 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           B2 => n24130, A => n27362, ZN => n27363);
   U1921 : OAI21_X1 port map( B1 => n24129, B2 => n1799, A => n27363, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1922 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN 
                           => n27516);
   U1923 : OAI22_X1 port map( A1 => n24003, A2 => n27516, B1 => n24169, B2 => 
                           n1797, ZN => n27364);
   U1924 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           B2 => n24130, A => n27364, ZN => n27365);
   U1925 : OAI21_X1 port map( B1 => n24129, B2 => n1798, A => n27365, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U1926 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN 
                           => n27517);
   U1927 : OAI22_X1 port map( A1 => n24003, A2 => n27517, B1 => n24169, B2 => 
                           n1796, ZN => n27366);
   U1928 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           B2 => n24130, A => n27366, ZN => n27367);
   U1929 : OAI21_X1 port map( B1 => n24129, B2 => n1797, A => n27367, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U1930 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN 
                           => n27518);
   U1931 : OAI22_X1 port map( A1 => n24003, A2 => n27518, B1 => n24169, B2 => 
                           n1795, ZN => n27368);
   U1932 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           B2 => n24130, A => n27368, ZN => n27369);
   U1933 : OAI21_X1 port map( B1 => n24129, B2 => n1796, A => n27369, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U1934 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN 
                           => n27519);
   U1935 : OAI22_X1 port map( A1 => n24003, A2 => n27519, B1 => n24169, B2 => 
                           n1794, ZN => n27370);
   U1936 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           B2 => n24130, A => n27370, ZN => n27371);
   U1937 : OAI21_X1 port map( B1 => n24129, B2 => n1795, A => n27371, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U1938 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN 
                           => n27520);
   U1939 : OAI22_X1 port map( A1 => n24003, A2 => n27520, B1 => n24169, B2 => 
                           n1793, ZN => n27372);
   U1940 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           B2 => n24130, A => n27372, ZN => n27373);
   U1941 : OAI21_X1 port map( B1 => n24129, B2 => n1794, A => n27373, ZN => 
                           n14145);
   U1942 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN 
                           => n27521);
   U1943 : OAI22_X1 port map( A1 => n24003, A2 => n27521, B1 => n24169, B2 => 
                           n1792, ZN => n27374);
   U1944 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           B2 => n24130, A => n27374, ZN => n27375);
   U1945 : OAI21_X1 port map( B1 => n24129, B2 => n1793, A => n27375, ZN => 
                           n19163);
   U1946 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN 
                           => n27523);
   U1947 : OAI22_X1 port map( A1 => n24003, A2 => n27523, B1 => n24169, B2 => 
                           n1791, ZN => n27376);
   U1948 : AOI21_X1 port map( B1 => n25894, B2 => n24130, A => n27376, ZN => 
                           n27377);
   U1949 : OAI21_X1 port map( B1 => n24129, B2 => n1792, A => n27377, ZN => 
                           n19162);
   U1950 : OAI22_X1 port map( A1 => n24003, A2 => n25893, B1 => n24169, B2 => 
                           n1790, ZN => n27378);
   U1951 : AOI21_X1 port map( B1 => n25896, B2 => n24130, A => n27378, ZN => 
                           n27379);
   U1952 : OAI21_X1 port map( B1 => n24129, B2 => n1791, A => n27379, ZN => 
                           n19161);
   U1953 : OAI222_X1 port map( A1 => n25895, A2 => n24003, B1 => n1790, B2 => 
                           n24026, C1 => n23973, C2 => n27443, ZN => n18846);
   U1954 : NAND3_X1 port map( A1 => n7769, A2 => n8978, A3 => n27380, ZN => 
                           n19160);
   U1955 : AOI22_X1 port map( A1 => n25900, A2 => n24027, B1 => n9084, B2 => 
                           n24128, ZN => n27381);
   U1956 : OAI221_X1 port map( B1 => n1807, B2 => n24002, C1 => n1807, C2 => 
                           n24100, A => n27381, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U1957 : AOI22_X1 port map( A1 => n25900, A2 => n23890, B1 => n9081, B2 => 
                           n24128, ZN => n27383);
   U1958 : NAND2_X1 port map( A1 => n25898, A2 => n24027, ZN => n27382);
   U1959 : OAI211_X1 port map( C1 => n24002, C2 => n1805, A => n27383, B => 
                           n27382, ZN => boothmul_pipelined_i_mux_out_4_10_port
                           );
   U1960 : AOI22_X1 port map( A1 => n9078, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n24027, ZN => n27385);
   U1961 : NAND2_X1 port map( A1 => n25898, A2 => n23890, ZN => n27384);
   U1962 : OAI211_X1 port map( C1 => n24002, C2 => n1804, A => n27385, B => 
                           n27384, ZN => boothmul_pipelined_i_mux_out_4_11_port
                           );
   U1963 : AOI22_X1 port map( A1 => n9075, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n24027, ZN => n27387);
   U1964 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n23890, ZN => n27386);
   U1965 : OAI211_X1 port map( C1 => n24002, C2 => n1803, A => n27387, B => 
                           n27386, ZN => boothmul_pipelined_i_mux_out_4_12_port
                           );
   U1966 : AOI22_X1 port map( A1 => n9072, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n24027, ZN => n27389);
   U1967 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n23890, ZN => n27388);
   U1968 : OAI211_X1 port map( C1 => n24002, C2 => n1802, A => n27389, B => 
                           n27388, ZN => boothmul_pipelined_i_mux_out_4_13_port
                           );
   U1969 : AOI22_X1 port map( A1 => n9069, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n24027, ZN => n27391);
   U1970 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n23890, ZN => n27390);
   U1971 : OAI211_X1 port map( C1 => n24002, C2 => n1800, A => n27391, B => 
                           n27390, ZN => boothmul_pipelined_i_mux_out_4_14_port
                           );
   U1972 : AOI22_X1 port map( A1 => n9066, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n24027, ZN => n27393);
   U1973 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n23890, ZN => n27392);
   U1974 : OAI211_X1 port map( C1 => n24002, C2 => n1799, A => n27393, B => 
                           n27392, ZN => boothmul_pipelined_i_mux_out_4_15_port
                           );
   U1975 : AOI22_X1 port map( A1 => n9063, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n24027, ZN => n27395);
   U1976 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n23890, ZN => n27394);
   U1977 : OAI211_X1 port map( C1 => n24002, C2 => n1798, A => n27395, B => 
                           n27394, ZN => n8928);
   U1978 : AOI22_X1 port map( A1 => n9060, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n24027, ZN => n27397);
   U1979 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n23890, ZN => n27396);
   U1980 : OAI211_X1 port map( C1 => n24002, C2 => n1797, A => n27397, B => 
                           n27396, ZN => n18899);
   U1981 : AOI22_X1 port map( A1 => n9057, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n24027, ZN => n27399);
   U1982 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n23890, ZN => n27398);
   U1983 : OAI211_X1 port map( C1 => n24002, C2 => n1796, A => n27399, B => 
                           n27398, ZN => n18898);
   U1984 : AOI22_X1 port map( A1 => n9054, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n24027, ZN => n27401);
   U1985 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n23890, ZN => n27400);
   U1986 : OAI211_X1 port map( C1 => n24002, C2 => n1795, A => n27401, B => 
                           n27400, ZN => n18897);
   U1987 : AOI22_X1 port map( A1 => n9051, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n24027, ZN => n27403);
   U1988 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n23890, ZN => n27402);
   U1989 : OAI211_X1 port map( C1 => n24002, C2 => n1794, A => n27403, B => 
                           n27402, ZN => n18896);
   U1990 : AOI22_X1 port map( A1 => n9048, A2 => n24128, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n24027, ZN => n27405);
   U1991 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n23890, ZN => n27404);
   U1992 : OAI211_X1 port map( C1 => n24002, C2 => n1793, A => n27405, B => 
                           n27404, ZN => n18895);
   U1993 : AOI22_X1 port map( A1 => n9045, A2 => n24128, B1 => n25894, B2 => 
                           n24027, ZN => n27407);
   U1994 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n23890, ZN => n27406);
   U1995 : OAI211_X1 port map( C1 => n24002, C2 => n1792, A => n27407, B => 
                           n27406, ZN => n18894);
   U1996 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n24128, B1 => 
                           n25896, B2 => n24027, ZN => n27409);
   U1997 : NAND2_X1 port map( A1 => n25894, A2 => n23890, ZN => n27408);
   U1998 : OAI211_X1 port map( C1 => n24002, C2 => n1791, A => n27409, B => 
                           n27408, ZN => n18893);
   U1999 : AOI22_X1 port map( A1 => n25896, A2 => n23890, B1 => n24027, B2 => 
                           n27527, ZN => n27410);
   U2000 : OAI221_X1 port map( B1 => n1790, B2 => n24002, C1 => n1790, C2 => 
                           n23978, A => n27410, ZN => n18852);
   U2001 : NOR2_X1 port map( A1 => n4302, A2 => n14286, ZN => n27411);
   U2002 : NAND2_X1 port map( A1 => n14287, A2 => n27411, ZN => n19250);
   U2003 : AOI22_X1 port map( A1 => n25900, A2 => n24088, B1 => n9084, B2 => 
                           n24000, ZN => n27412);
   U2004 : OAI221_X1 port map( B1 => n1807, B2 => n24001, C1 => n1807, C2 => 
                           n24127, A => n27412, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2005 : OAI22_X1 port map( A1 => n24001, A2 => n25899, B1 => n24127, B2 => 
                           n1805, ZN => n27413);
   U2006 : AOI21_X1 port map( B1 => n9081, B2 => n24000, A => n27413, ZN => 
                           n27414);
   U2007 : OAI21_X1 port map( B1 => n24037, B2 => n25897, A => n27414, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2008 : OAI22_X1 port map( A1 => n24037, A2 => n27512, B1 => n24127, B2 => 
                           n1804, ZN => n27415);
   U2009 : AOI21_X1 port map( B1 => n9078, B2 => n24000, A => n27415, ZN => 
                           n27416);
   U2010 : OAI21_X1 port map( B1 => n24001, B2 => n25897, A => n27416, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2011 : OAI22_X1 port map( A1 => n24037, A2 => n27513, B1 => n24001, B2 => 
                           n27512, ZN => n27417);
   U2012 : AOI21_X1 port map( B1 => n9075, B2 => n24000, A => n27417, ZN => 
                           n27418);
   U2013 : OAI21_X1 port map( B1 => n24127, B2 => n1803, A => n27418, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2014 : OAI22_X1 port map( A1 => n24037, A2 => n27514, B1 => n24001, B2 => 
                           n27513, ZN => n27419);
   U2015 : AOI21_X1 port map( B1 => n9072, B2 => n24000, A => n27419, ZN => 
                           n27420);
   U2016 : OAI21_X1 port map( B1 => n24127, B2 => n1802, A => n27420, ZN => 
                           n19158);
   U2017 : OAI22_X1 port map( A1 => n24037, A2 => n27515, B1 => n24001, B2 => 
                           n27514, ZN => n27421);
   U2018 : AOI21_X1 port map( B1 => n9069, B2 => n24000, A => n27421, ZN => 
                           n27422);
   U2019 : OAI21_X1 port map( B1 => n24127, B2 => n1800, A => n27422, ZN => 
                           n19157);
   U2020 : OAI22_X1 port map( A1 => n24037, A2 => n27516, B1 => n24001, B2 => 
                           n27515, ZN => n27423);
   U2021 : AOI21_X1 port map( B1 => n9066, B2 => n24000, A => n27423, ZN => 
                           n27424);
   U2022 : OAI21_X1 port map( B1 => n24127, B2 => n1799, A => n27424, ZN => 
                           n19156);
   U2023 : OAI22_X1 port map( A1 => n24037, A2 => n27517, B1 => n24001, B2 => 
                           n27516, ZN => n27425);
   U2024 : AOI21_X1 port map( B1 => n9063, B2 => n24000, A => n27425, ZN => 
                           n27426);
   U2025 : OAI21_X1 port map( B1 => n24127, B2 => n1798, A => n27426, ZN => 
                           n19155);
   U2026 : OAI22_X1 port map( A1 => n24037, A2 => n27518, B1 => n24001, B2 => 
                           n27517, ZN => n27427);
   U2027 : AOI21_X1 port map( B1 => n9060, B2 => n24000, A => n27427, ZN => 
                           n27428);
   U2028 : OAI21_X1 port map( B1 => n24127, B2 => n1797, A => n27428, ZN => 
                           n19154);
   U2029 : OAI22_X1 port map( A1 => n24037, A2 => n27519, B1 => n24001, B2 => 
                           n27518, ZN => n27429);
   U2030 : AOI21_X1 port map( B1 => n9057, B2 => n24000, A => n27429, ZN => 
                           n27430);
   U2031 : OAI21_X1 port map( B1 => n24127, B2 => n1796, A => n27430, ZN => 
                           n19153);
   U2032 : OAI22_X1 port map( A1 => n24037, A2 => n27520, B1 => n24001, B2 => 
                           n27519, ZN => n27431);
   U2033 : AOI21_X1 port map( B1 => n9054, B2 => n24000, A => n27431, ZN => 
                           n27432);
   U2034 : OAI21_X1 port map( B1 => n24127, B2 => n1795, A => n27432, ZN => 
                           n19152);
   U2035 : OAI22_X1 port map( A1 => n24037, A2 => n27521, B1 => n24001, B2 => 
                           n27520, ZN => n27433);
   U2036 : AOI21_X1 port map( B1 => n9051, B2 => n24000, A => n27433, ZN => 
                           n27434);
   U2037 : OAI21_X1 port map( B1 => n24127, B2 => n1794, A => n27434, ZN => 
                           n19151);
   U2038 : OAI22_X1 port map( A1 => n24037, A2 => n27523, B1 => n24001, B2 => 
                           n27521, ZN => n27435);
   U2039 : AOI21_X1 port map( B1 => n9048, B2 => n24000, A => n27435, ZN => 
                           n27436);
   U2040 : OAI21_X1 port map( B1 => n24127, B2 => n1793, A => n27436, ZN => 
                           n19150);
   U2041 : OAI22_X1 port map( A1 => n24037, A2 => n25893, B1 => n24001, B2 => 
                           n27523, ZN => n27437);
   U2042 : AOI21_X1 port map( B1 => n9045, B2 => n24000, A => n27437, ZN => 
                           n27438);
   U2043 : OAI21_X1 port map( B1 => n24127, B2 => n1792, A => n27438, ZN => 
                           n19149);
   U2044 : OAI22_X1 port map( A1 => n24037, A2 => n25895, B1 => n24001, B2 => 
                           n25893, ZN => n27439);
   U2045 : AOI21_X1 port map( B1 => data1_mul_15_port, B2 => n24000, A => 
                           n27439, ZN => n27440);
   U2046 : OAI21_X1 port map( B1 => n24127, B2 => n1791, A => n27440, ZN => 
                           n19148);
   U2047 : NAND2_X1 port map( A1 => n4302, A2 => n14286, ZN => n27441);
   U2048 : OAI21_X1 port map( B1 => n4302, B2 => n14286, A => n27441, ZN => 
                           n17932);
   U2049 : NOR2_X1 port map( A1 => n14287, A2 => n17932, ZN => n19291);
   U2050 : INV_X1 port map( A => n1810, ZN => n27442);
   U2051 : NOR2_X1 port map( A1 => n27442, A2 => n19291, ZN => n19248);
   U2052 : OAI222_X1 port map( A1 => n25895, A2 => n24001, B1 => n1790, B2 => 
                           n23999, C1 => n24037, C2 => n27443, ZN => n18845);
   U2053 : AOI22_X1 port map( A1 => n25900, A2 => n24043, B1 => n9084, B2 => 
                           n24042, ZN => n27444);
   U2054 : OAI221_X1 port map( B1 => n1807, B2 => n23897, C1 => n1807, C2 => 
                           n23998, A => n27444, ZN => n18851);
   U2055 : AOI22_X1 port map( A1 => n25900, A2 => n24133, B1 => n9081, B2 => 
                           n24042, ZN => n27446);
   U2056 : NAND2_X1 port map( A1 => n25898, A2 => n24043, ZN => n27445);
   U2057 : OAI211_X1 port map( C1 => n23897, C2 => n1805, A => n27446, B => 
                           n27445, ZN => n19247);
   U2058 : AOI22_X1 port map( A1 => n9078, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n24043, ZN => n27448);
   U2059 : NAND2_X1 port map( A1 => n25898, A2 => n24133, ZN => n27447);
   U2060 : OAI211_X1 port map( C1 => n23897, C2 => n1804, A => n27448, B => 
                           n27447, ZN => n19246);
   U2061 : AOI22_X1 port map( A1 => n9075, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n24043, ZN => n27450);
   U2062 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n24133, ZN => n27449);
   U2063 : OAI211_X1 port map( C1 => n23897, C2 => n1803, A => n27450, B => 
                           n27449, ZN => n19245);
   U2064 : AOI22_X1 port map( A1 => n9072, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n24043, ZN => n27452);
   U2065 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n24133, ZN => n27451);
   U2066 : OAI211_X1 port map( C1 => n23897, C2 => n1802, A => n27452, B => 
                           n27451, ZN => n19244);
   U2067 : AOI22_X1 port map( A1 => n9069, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n24043, ZN => n27454);
   U2068 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n24133, ZN => n27453);
   U2069 : OAI211_X1 port map( C1 => n23897, C2 => n1800, A => n27454, B => 
                           n27453, ZN => n19243);
   U2070 : AOI22_X1 port map( A1 => n9066, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n24043, ZN => n27456);
   U2071 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n24133, ZN => n27455);
   U2072 : OAI211_X1 port map( C1 => n23897, C2 => n1799, A => n27456, B => 
                           n27455, ZN => n19242);
   U2073 : AOI22_X1 port map( A1 => n9063, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n24043, ZN => n27458);
   U2074 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n24133, ZN => n27457);
   U2075 : OAI211_X1 port map( C1 => n23897, C2 => n1798, A => n27458, B => 
                           n27457, ZN => n19241);
   U2076 : AOI22_X1 port map( A1 => n9060, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n24043, ZN => n27460);
   U2077 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n24133, ZN => n27459);
   U2078 : OAI211_X1 port map( C1 => n23897, C2 => n1797, A => n27460, B => 
                           n27459, ZN => n19240);
   U2079 : AOI22_X1 port map( A1 => n9057, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n24043, ZN => n27462);
   U2080 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n24133, ZN => n27461);
   U2081 : OAI211_X1 port map( C1 => n23897, C2 => n1796, A => n27462, B => 
                           n27461, ZN => n19239);
   U2082 : AOI22_X1 port map( A1 => n9054, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n24043, ZN => n27464);
   U2083 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n24133, ZN => n27463);
   U2084 : OAI211_X1 port map( C1 => n23897, C2 => n1795, A => n27464, B => 
                           n27463, ZN => n19238);
   U2085 : AOI22_X1 port map( A1 => n9051, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n24043, ZN => n27466);
   U2086 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n24133, ZN => n27465);
   U2087 : OAI211_X1 port map( C1 => n23897, C2 => n1794, A => n27466, B => 
                           n27465, ZN => n19237);
   U2088 : AOI22_X1 port map( A1 => n9048, A2 => n24042, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n24043, ZN => n27468);
   U2089 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n24133, ZN => n27467);
   U2090 : OAI211_X1 port map( C1 => n23897, C2 => n1793, A => n27468, B => 
                           n27467, ZN => n19236);
   U2091 : AOI22_X1 port map( A1 => n9045, A2 => n24042, B1 => n25894, B2 => 
                           n24043, ZN => n27470);
   U2092 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n24133, ZN => n27469);
   U2093 : OAI211_X1 port map( C1 => n23897, C2 => n1792, A => n27470, B => 
                           n27469, ZN => n19235);
   U2094 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n24042, B1 => 
                           n25896, B2 => n24043, ZN => n27472);
   U2095 : NAND2_X1 port map( A1 => n25894, A2 => n24133, ZN => n27471);
   U2096 : OAI211_X1 port map( C1 => n23897, C2 => n1791, A => n27472, B => 
                           n27471, ZN => n18892);
   U2097 : AOI22_X1 port map( A1 => n25896, A2 => n24133, B1 => n24043, B2 => 
                           n27527, ZN => n27473);
   U2098 : OAI221_X1 port map( B1 => n1790, B2 => n23897, C1 => n1790, C2 => 
                           n24132, A => n27473, ZN => n18850);
   U2099 : OR2_X1 port map( A1 => n27474, A2 => n27700, ZN => n27509);
   U2100 : INV_X1 port map( A => n27507, ZN => n27476);
   U2101 : AOI22_X1 port map( A1 => n25900, A2 => n27506, B1 => n9084, B2 => 
                           n27505, ZN => n27475);
   U2102 : OAI221_X1 port map( B1 => n1807, B2 => n27509, C1 => n1807, C2 => 
                           n27476, A => n27475, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2103 : AOI22_X1 port map( A1 => n25898, A2 => n27506, B1 => n25900, B2 => 
                           n27507, ZN => n27478);
   U2104 : NAND2_X1 port map( A1 => n9081, A2 => n27505, ZN => n27477);
   U2105 : OAI211_X1 port map( C1 => n27509, C2 => n1805, A => n27478, B => 
                           n27477, ZN => boothmul_pipelined_i_mux_out_7_16_port
                           );
   U2106 : AOI22_X1 port map( A1 => n25898, A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n27506, ZN => n27480);
   U2107 : NAND2_X1 port map( A1 => n9078, A2 => n27505, ZN => n27479);
   U2108 : OAI211_X1 port map( C1 => n27509, C2 => n1804, A => n27480, B => 
                           n27479, ZN => boothmul_pipelined_i_mux_out_7_17_port
                           );
   U2109 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n27506, ZN => n27482);
   U2110 : NAND2_X1 port map( A1 => n9075, A2 => n27505, ZN => n27481);
   U2111 : OAI211_X1 port map( C1 => n27509, C2 => n1803, A => n27482, B => 
                           n27481, ZN => boothmul_pipelined_i_mux_out_7_18_port
                           );
   U2112 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n27506, ZN => n27484);
   U2113 : NAND2_X1 port map( A1 => n9072, A2 => n27505, ZN => n27483);
   U2114 : OAI211_X1 port map( C1 => n27509, C2 => n1802, A => n27484, B => 
                           n27483, ZN => boothmul_pipelined_i_mux_out_7_19_port
                           );
   U2115 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n27506, ZN => n27486);
   U2116 : NAND2_X1 port map( A1 => n9069, A2 => n27505, ZN => n27485);
   U2117 : OAI211_X1 port map( C1 => n27509, C2 => n1800, A => n27486, B => 
                           n27485, ZN => boothmul_pipelined_i_mux_out_7_20_port
                           );
   U2118 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n27506, ZN => n27488);
   U2119 : NAND2_X1 port map( A1 => n9066, A2 => n27505, ZN => n27487);
   U2120 : OAI211_X1 port map( C1 => n27509, C2 => n1799, A => n27488, B => 
                           n27487, ZN => boothmul_pipelined_i_mux_out_7_21_port
                           );
   U2121 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n27506, ZN => n27490);
   U2122 : NAND2_X1 port map( A1 => n9063, A2 => n27505, ZN => n27489);
   U2123 : OAI211_X1 port map( C1 => n27509, C2 => n1798, A => n27490, B => 
                           n27489, ZN => boothmul_pipelined_i_mux_out_7_22_port
                           );
   U2124 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n27506, ZN => n27492);
   U2125 : NAND2_X1 port map( A1 => n9060, A2 => n27505, ZN => n27491);
   U2126 : OAI211_X1 port map( C1 => n27509, C2 => n1797, A => n27492, B => 
                           n27491, ZN => boothmul_pipelined_i_mux_out_7_23_port
                           );
   U2127 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n27506, ZN => n27494);
   U2128 : NAND2_X1 port map( A1 => n9057, A2 => n27505, ZN => n27493);
   U2129 : OAI211_X1 port map( C1 => n27509, C2 => n1796, A => n27494, B => 
                           n27493, ZN => boothmul_pipelined_i_mux_out_7_24_port
                           );
   U2130 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n27506, ZN => n27496);
   U2131 : NAND2_X1 port map( A1 => n9054, A2 => n27505, ZN => n27495);
   U2132 : OAI211_X1 port map( C1 => n27509, C2 => n1795, A => n27496, B => 
                           n27495, ZN => boothmul_pipelined_i_mux_out_7_25_port
                           );
   U2133 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n27506, ZN => n27498);
   U2134 : NAND2_X1 port map( A1 => n9051, A2 => n27505, ZN => n27497);
   U2135 : OAI211_X1 port map( C1 => n27509, C2 => n1794, A => n27498, B => 
                           n27497, ZN => boothmul_pipelined_i_mux_out_7_26_port
                           );
   U2136 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n27507, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n27506, ZN => n27500);
   U2137 : NAND2_X1 port map( A1 => n9048, A2 => n27505, ZN => n27499);
   U2138 : OAI211_X1 port map( C1 => n27509, C2 => n1793, A => n27500, B => 
                           n27499, ZN => n19234);
   U2139 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n27507, B1 => n25894, B2 => n27506, ZN => 
                           n27502);
   U2140 : NAND2_X1 port map( A1 => n9045, A2 => n27505, ZN => n27501);
   U2141 : OAI211_X1 port map( C1 => n27509, C2 => n1792, A => n27502, B => 
                           n27501, ZN => n19233);
   U2142 : AOI22_X1 port map( A1 => n25894, A2 => n27507, B1 => n25896, B2 => 
                           n27506, ZN => n27504);
   U2143 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n27505, ZN => 
                           n27503);
   U2144 : OAI211_X1 port map( C1 => n27509, C2 => n1791, A => n27504, B => 
                           n27503, ZN => n19232);
   U2145 : INV_X1 port map( A => n27505, ZN => n27510);
   U2146 : AOI22_X1 port map( A1 => n25896, A2 => n27507, B1 => n27506, B2 => 
                           n27527, ZN => n27508);
   U2147 : OAI221_X1 port map( B1 => n1790, B2 => n27510, C1 => n1790, C2 => 
                           n27509, A => n27508, ZN => n19231);
   U2148 : INV_X1 port map( A => n27511, ZN => n27530);
   U2149 : OAI222_X1 port map( A1 => n1807, A2 => n27522, B1 => n25899, B2 => 
                           n27524, C1 => n27530, C2 => n1805, ZN => n18839);
   U2150 : OAI222_X1 port map( A1 => n25897, A2 => n27522, B1 => n27512, B2 => 
                           n27524, C1 => n1803, C2 => n27530, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2151 : OAI222_X1 port map( A1 => n1802, A2 => n27530, B1 => n27513, B2 => 
                           n27524, C1 => n27512, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2152 : OAI222_X1 port map( A1 => n1800, A2 => n27530, B1 => n27514, B2 => 
                           n27524, C1 => n27513, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2153 : OAI222_X1 port map( A1 => n1799, A2 => n27530, B1 => n27515, B2 => 
                           n27524, C1 => n27514, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2154 : OAI222_X1 port map( A1 => n1798, A2 => n27530, B1 => n27516, B2 => 
                           n27524, C1 => n27515, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2155 : OAI222_X1 port map( A1 => n1797, A2 => n27530, B1 => n27517, B2 => 
                           n27524, C1 => n27516, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2156 : OAI222_X1 port map( A1 => n1796, A2 => n27530, B1 => n27518, B2 => 
                           n27524, C1 => n27517, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2157 : OAI222_X1 port map( A1 => n1795, A2 => n27530, B1 => n27519, B2 => 
                           n27524, C1 => n27518, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2158 : OAI222_X1 port map( A1 => n1794, A2 => n27530, B1 => n27520, B2 => 
                           n27524, C1 => n27519, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2159 : OAI222_X1 port map( A1 => n1793, A2 => n27530, B1 => n27521, B2 => 
                           n27524, C1 => n27520, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2160 : OAI222_X1 port map( A1 => n1792, A2 => n27530, B1 => n27523, B2 => 
                           n27524, C1 => n27521, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2161 : OAI222_X1 port map( A1 => n1791, A2 => n27530, B1 => n25893, B2 => 
                           n27524, C1 => n27523, C2 => n27522, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2162 : AOI22_X1 port map( A1 => n27528, A2 => n25896, B1 => n27526, B2 => 
                           n25894, ZN => n27525);
   U2163 : OAI21_X1 port map( B1 => n27530, B2 => n1790, A => n27525, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2164 : AOI22_X1 port map( A1 => n27528, A2 => n27527, B1 => n27526, B2 => 
                           n25896, ZN => n27529);
   U2165 : OAI21_X1 port map( B1 => n27530, B2 => n1790, A => n27529, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U2166 : XNOR2_X1 port map( A => n27532, B => n27531, ZN => n19147);
   U2167 : AOI21_X1 port map( B1 => n24178, B2 => n27652, A => n27651, ZN => 
                           n27535);
   U2168 : OAI22_X1 port map( A1 => n27535, A2 => n27534, B1 => n27533, B2 => 
                           n27570, ZN => n27541);
   U2169 : NAND3_X1 port map( A1 => n1831, A2 => n27624, A3 => n27536, ZN => 
                           n27537);
   U2170 : OAI21_X1 port map( B1 => n27539, B2 => n27538, A => n27537, ZN => 
                           n27540);
   U2171 : AOI211_X1 port map( C1 => n27542, C2 => n23618, A => n27541, B => 
                           n27540, ZN => n18882);
   U2172 : OAI22_X1 port map( A1 => n24103, A2 => n27544, B1 => n23966, B2 => 
                           n27543, ZN => n27545);
   U2173 : INV_X1 port map( A => n27545, ZN => n27546);
   U2174 : OAI211_X1 port map( C1 => n24036, C2 => n27546, A => n23896, B => 
                           n24031, ZN => OUTALU(6));
   U2175 : NOR3_X1 port map( A1 => n27549, A2 => n27548, A3 => n27547, ZN => 
                           n27555);
   U2176 : AOI211_X1 port map( C1 => n27553, C2 => n27552, A => n27551, B => 
                           n27550, ZN => n27554);
   U2177 : AOI211_X1 port map( C1 => n27557, C2 => n27556, A => n27555, B => 
                           n27554, ZN => n18878);
   U2178 : AOI22_X1 port map( A1 => n27648, A2 => n27646, B1 => n27649, B2 => 
                           n27558, ZN => n18877);
   U2179 : OAI22_X1 port map( A1 => n27641, A2 => n27596, B1 => n27559, B2 => 
                           n27636, ZN => n27562);
   U2180 : OAI22_X1 port map( A1 => n26425, A2 => n27616, B1 => n27560, B2 => 
                           n27607, ZN => n27561);
   U2181 : AOI211_X1 port map( C1 => n27709, C2 => n27563, A => n27562, B => 
                           n27561, ZN => n1834);
   U2182 : OAI22_X1 port map( A1 => n1842, A2 => n27564, B1 => n1834, B2 => 
                           n1836, ZN => n19419);
   U2183 : NOR2_X1 port map( A1 => n27566, A2 => n27565, ZN => n27569);
   U2184 : NAND2_X1 port map( A1 => n27567, A2 => n23801, ZN => n27568);
   U2185 : OAI21_X1 port map( B1 => n27570, B2 => n27569, A => n27568, ZN => 
                           n19433);
   U2186 : AOI22_X1 port map( A1 => n27575, A2 => DATA2(4), B1 => n27592, B2 =>
                           n27571, ZN => n27572);
   U2187 : NAND3_X1 port map( A1 => n1866, A2 => n27572, A3 => n27583, ZN => 
                           n25859);
   U2188 : NAND4_X1 port map( A1 => DATA2(1), A2 => n27574, A3 => n27594, A4 =>
                           n27573, ZN => n25865);
   U2189 : OAI21_X1 port map( B1 => DATA2(2), B2 => DATA2(1), A => n27581, ZN 
                           => n25866);
   U2190 : INV_X1 port map( A => n27574, ZN => n27576);
   U2191 : NOR3_X1 port map( A1 => DATA2(3), A2 => n27579, A3 => n27576, ZN => 
                           n25867);
   U2192 : NAND2_X1 port map( A1 => DATA2(1), A2 => n27578, ZN => n25868);
   U2193 : NAND3_X1 port map( A1 => n27575, A2 => n27581, A3 => n27592, ZN => 
                           n25869);
   U2194 : NOR4_X1 port map( A1 => DATA2(2), A2 => DATA2(3), A3 => n1863, A4 =>
                           n27579, ZN => n25870);
   U2195 : NOR3_X1 port map( A1 => DATA2(3), A2 => n27591, A3 => n27576, ZN => 
                           n25871);
   U2196 : NOR4_X1 port map( A1 => DATA2(2), A2 => DATA2(3), A3 => n27577, A4 
                           => n27591, ZN => n25873);
   U2197 : INV_X1 port map( A => n27578, ZN => n27582);
   U2198 : NOR2_X1 port map( A1 => n27582, A2 => n27579, ZN => n25874);
   U2199 : NAND3_X1 port map( A1 => n27581, A2 => n27580, A3 => n27592, ZN => 
                           n25875);
   U2200 : NOR2_X1 port map( A1 => n27593, A2 => n27582, ZN => n25876);
   U2201 : NOR2_X1 port map( A1 => n27583, A2 => n1841, ZN => n25879);
   U2202 : NAND2_X1 port map( A1 => n4302, A2 => n27584, ZN => n25881);
   U2203 : OR2_X1 port map( A1 => n22765, A2 => n19293, ZN => n25882);
   U2204 : NOR3_X1 port map( A1 => n14287, A2 => n19292, A3 => n1808, ZN => 
                           n25883);
   U2205 : NOR2_X1 port map( A1 => n27586, A2 => n27585, ZN => n25885);
   U2206 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           A3 => n27587, ZN => n25886);
   U2207 : NOR2_X1 port map( A1 => n4302, A2 => n27588, ZN => n25887);
   U2208 : NOR2_X1 port map( A1 => n27589, A2 => n17932, ZN => n25888);
   U2209 : AOI21_X1 port map( B1 => n27592, B2 => n27591, A => n27590, ZN => 
                           n1870);
   U2210 : NOR2_X1 port map( A1 => DATA2(2), A2 => n27593, ZN => n27595);
   U2211 : AOI21_X1 port map( B1 => n27595, B2 => n27594, A => n1863, ZN => 
                           n1868);
   U2212 : OAI22_X1 port map( A1 => n27636, A2 => n27597, B1 => n27638, B2 => 
                           n27596, ZN => n27598);
   U2213 : INV_X1 port map( A => n27598, ZN => n27602);
   U2214 : AOI22_X1 port map( A1 => n25892, A2 => n27600, B1 => n27645, B2 => 
                           n27599, ZN => n27601);
   U2215 : OAI211_X1 port map( C1 => n27641, C2 => n27603, A => n27602, B => 
                           n27601, ZN => n1839);
   U2216 : AOI22_X1 port map( A1 => n27632, A2 => n27612, B1 => n27624, B2 => 
                           n27610, ZN => n27606);
   U2217 : AOI22_X1 port map( A1 => n27709, A2 => n27611, B1 => n27645, B2 => 
                           n27604, ZN => n27605);
   U2218 : OAI211_X1 port map( C1 => n27608, C2 => n27607, A => n27606, B => 
                           n27605, ZN => n1838);
   U2219 : AOI22_X1 port map( A1 => n25892, A2 => n27610, B1 => n27632, B2 => 
                           n27609, ZN => n27614);
   U2220 : AOI22_X1 port map( A1 => n27709, A2 => n27612, B1 => n27645, B2 => 
                           n27611, ZN => n27613);
   U2221 : OAI211_X1 port map( C1 => n27641, C2 => n27615, A => n27614, B => 
                           n27613, ZN => n1835);
   U2222 : INV_X1 port map( A => n27616, ZN => n27618);
   U2223 : AOI22_X1 port map( A1 => n25892, A2 => n27618, B1 => n27617, B2 => 
                           n27645, ZN => n27622);
   U2224 : AOI22_X1 port map( A1 => n27632, A2 => n27620, B1 => n27709, B2 => 
                           n27619, ZN => n27621);
   U2225 : OAI211_X1 port map( C1 => n27641, C2 => n27623, A => n27622, B => 
                           n27621, ZN => n1833);
   U2226 : INV_X1 port map( A => n27637, ZN => n27629);
   U2227 : AOI22_X1 port map( A1 => n27709, A2 => n27630, B1 => n27624, B2 => 
                           n27629, ZN => n27627);
   U2228 : INV_X1 port map( A => n27639, ZN => n27631);
   U2229 : AOI22_X1 port map( A1 => n25892, A2 => n27631, B1 => n27645, B2 => 
                           n27625, ZN => n27626);
   U2230 : OAI211_X1 port map( C1 => n27628, C2 => n27636, A => n27627, B => 
                           n27626, ZN => n1829);
   U2231 : INV_X1 port map( A => n27628, ZN => n27644);
   U2232 : AOI22_X1 port map( A1 => n25892, A2 => n27629, B1 => n27709, B2 => 
                           n27644, ZN => n27634);
   U2233 : AOI22_X1 port map( A1 => n27632, A2 => n27631, B1 => n27645, B2 => 
                           n27630, ZN => n27633);
   U2234 : OAI211_X1 port map( C1 => n27641, C2 => n27635, A => n27634, B => 
                           n27633, ZN => n1827);
   U2235 : OAI22_X1 port map( A1 => n27637, A2 => n27636, B1 => n27635, B2 => 
                           n27607, ZN => n27643);
   U2236 : OAI22_X1 port map( A1 => n27641, A2 => n27640, B1 => n27639, B2 => 
                           n27638, ZN => n27642);
   U2237 : AOI211_X1 port map( C1 => n27645, C2 => n27644, A => n27643, B => 
                           n27642, ZN => n1818);
   U2238 : INV_X1 port map( A => n27646, ZN => n27647);
   U2239 : AOI22_X1 port map( A1 => n27650, A2 => n27649, B1 => n27648, B2 => 
                           n27647, ZN => n27656);
   U2240 : INV_X1 port map( A => n1809, ZN => n27655);
   U2241 : AOI21_X1 port map( B1 => DATA2(21), B2 => n27652, A => n27651, ZN =>
                           n27654);
   U2242 : OAI22_X1 port map( A1 => n27656, A2 => n27655, B1 => n27654, B2 => 
                           n27653, ZN => n1788);
   U2243 : OAI22_X1 port map( A1 => n27660, A2 => n27659, B1 => n27658, B2 => 
                           n27657, ZN => n1786);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n40552, n40555, n40558, n40561, n40574, n40576, n40577, n40580, 
      n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, 
      n40591, n40592, n40604, n40605, n40606, n40607, n40608, n40609, n40610, 
      n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619, 
      n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628, 
      n40629, n40632, n40633, n40636, n40637, n40638, n40639, n40642, n40643, 
      n40646, n40647, n41686, n41687, n41688, n41689, n41690, n41691, n41692, 
      n47428, n47429, n47430, n47431, n49085, n49086, n49087, n49088, n49089, 
      n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097, n51364, 
      n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373, 
      n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382, 
      n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391, 
      n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400, 
      n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409, 
      n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418, 
      n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427, 
      n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436, 
      n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445, 
      n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454, 
      n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463, 
      n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472, 
      n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481, 
      n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490, 
      n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499, 
      n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508, 
      n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517, 
      n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526, 
      n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535, 
      n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544, 
      n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553, 
      n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562, 
      n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571, 
      n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580, 
      n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589, 
      n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598, 
      n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607, 
      n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616, 
      n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625, 
      n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634, 
      n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643, 
      n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652, 
      n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661, 
      n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670, 
      n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679, 
      n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688, 
      n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697, 
      n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706, 
      n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715, 
      n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724, 
      n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733, 
      n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742, 
      n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751, 
      n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760, 
      n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769, 
      n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778, 
      n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787, 
      n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796, 
      n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805, 
      n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814, 
      n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823, 
      n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832, 
      n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841, 
      n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850, 
      n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859, 
      n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868, 
      n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877, 
      n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886, 
      n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895, 
      n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904, 
      n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913, 
      n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922, 
      n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931, 
      n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940, 
      n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949, 
      n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958, 
      n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967, 
      n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976, 
      n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985, 
      n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994, 
      n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003, 
      n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012, 
      n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021, 
      n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030, 
      n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039, 
      n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048, 
      n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057, 
      n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066, 
      n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075, 
      n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084, 
      n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093, 
      n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102, 
      n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111, 
      n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120, 
      n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129, 
      n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138, 
      n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147, 
      n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156, 
      n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165, 
      n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174, 
      n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183, 
      n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192, 
      n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201, 
      n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210, 
      n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219, 
      n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228, 
      n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237, 
      n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246, 
      n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255, 
      n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264, 
      n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273, 
      n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282, 
      n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291, 
      n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300, 
      n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309, 
      n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318, 
      n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327, 
      n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336, 
      n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345, 
      n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354, 
      n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363, 
      n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372, 
      n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381, 
      n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390, 
      n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399, 
      n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408, 
      n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417, 
      n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426, 
      n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435, 
      n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444, 
      n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453, 
      n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462, 
      n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471, 
      n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480, 
      n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489, 
      n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498, 
      n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507, 
      n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516, 
      n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525, 
      n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534, 
      n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543, 
      n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552, 
      n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561, 
      n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570, 
      n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579, 
      n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588, 
      n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597, 
      n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606, 
      n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615, 
      n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624, 
      n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633, 
      n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642, 
      n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651, 
      n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660, 
      n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669, 
      n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678, 
      n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687, 
      n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696, 
      n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705, 
      n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714, 
      n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723, 
      n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732, 
      n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741, 
      n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750, 
      n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759, 
      n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768, 
      n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777, 
      n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786, 
      n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795, 
      n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804, 
      n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813, 
      n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822, 
      n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831, 
      n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840, 
      n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849, 
      n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858, 
      n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867, 
      n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876, 
      n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885, 
      n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894, 
      n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903, 
      n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912, 
      n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921, 
      n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930, 
      n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939, 
      n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948, 
      n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957, 
      n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966, 
      n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975, 
      n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984, 
      n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993, 
      n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002, 
      n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011, 
      n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020, 
      n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029, 
      n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038, 
      n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047, 
      n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056, 
      n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065, 
      n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074, 
      n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083, 
      n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092, 
      n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101, 
      n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110, 
      n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119, 
      n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128, 
      n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137, 
      n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146, 
      n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155, 
      n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164, 
      n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173, 
      n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182, 
      n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191, 
      n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200, 
      n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209, 
      n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218, 
      n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227, 
      n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236, 
      n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245, 
      n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, 
      n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263, 
      n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272, 
      n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281, 
      n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290, 
      n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299, 
      n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308, 
      n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317, 
      n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326, 
      n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335, 
      n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344, 
      n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353, 
      n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362, 
      n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371, 
      n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380, 
      n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389, 
      n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398, 
      n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407, 
      n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416, 
      n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425, 
      n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434, 
      n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443, 
      n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452, 
      n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461, 
      n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470, 
      n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479, 
      n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488, 
      n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497, 
      n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506, 
      n53509, n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, 
      n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, 
      n53528, n53529, n53530, n53531, n53533, n53534, n53535, n53536, n53537, 
      n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546, 
      n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555, 
      n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564, 
      n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573, 
      n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582, 
      n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591, 
      n53592, n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600, 
      n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609, 
      n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618, 
      n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627, 
      n53629, n58166, n58167, n58168, n58169, n2534, n2535, n2536, n2537, n2538
      , n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
      n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
      n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
      n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
      n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
      n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
      n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
      n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
      n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
      n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
      n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
      n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
      n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
      n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
      n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
      n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
      n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n58170, n58171, n58172, 
      n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180, n58181, 
      n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189, n58190, 
      n58191, n58192, n58193, n58194, n58195, n58196, n58197, n58198, n58199, 
      n58200, n58201, n58202, n58203, n58204, n58205, n58206, n58207, n58208, 
      n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58216, n58217, 
      n58218, n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226, 
      n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234, n58235, 
      n58236, n58237, n58238, n58239, n58240, n58241, n58242, n58243, n58244, 
      n58245, n58246, n58247, n58248, n58249, n58250, n58251, n58252, n58253, 
      n58254, n58255, n58256, n58257, n58258, n58259, n58260, n58261, n58262, 
      n58263, n58264, n58265, n58266, n58267, n58268, n58269, n58270, n58271, 
      n58272, n58273, n58274, n58275, n58276, n58277, n58278, n58279, n58280, 
      n58281, n58282, n58283, n58284, n58285, n58286, n58287, n58288, n58289, 
      n58290, n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298, 
      n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306, n58307, 
      n58308, n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316, 
      n58317, n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325, 
      n58326, n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334, 
      n58335, n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58343, 
      n58344, n58345, n58346, n58347, n58348, n58349, n58350, n58351, n58352, 
      n58353, n58354, n58355, n58356, n58357, n58358, n58359, n58360, n58361, 
      n58362, n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370, 
      n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378, n58379, 
      n58380, n58381, n58382, n58383, n58384, n58385, n58386, n58387, n58388, 
      n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396, n58397, 
      n58398, n58399, n58400, n58401, n58402, n58403, n58404, n58405, n58406, 
      n58407, n58408, n58409, n58410, n58411, n58412, n58413, n58414, n58415, 
      n58416, n58417, n58418, n58419, n58420, n58421, n58422, n58423, n58424, 
      n58425, n58426, n58427, n58428, n58429, n58430, n58431, n58432, n58433, 
      n58434, n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442, 
      n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450, n58451, 
      n58452, n58453, n58454, n58455, n58456, n58457, n58458, n58459, n58460, 
      n58461, n58462, n58463, n58464, n58465, n58466, n58467, n58468, n58469, 
      n58470, n58471, n58472, n58473, n58474, n58475, n58476, n58477, n58478, 
      n58479, n58480, n58481, n58482, n58483, n58484, n58485, n58486, n58487, 
      n58488, n58489, n58490, n58491, n58492, n58493, n58494, n58495, n58496, 
      n58497, n58498, n58499, n58500, n58501, n58502, n58503, n58504, n58505, 
      n58506, n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514, 
      n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522, n58523, 
      n58524, n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532, 
      n58533, n58534, n58535, n58536, n58537, n58538, n58539, n58540, n58541, 
      n58542, n58543, n58544, n58545, n58546, n58547, n58548, n58549, n58550, 
      n58551, n58552, n58553, n58554, n58555, n58556, n58557, n58558, n58559, 
      n58560, n58561, n58562, n58563, n58564, n58565, n58566, n58567, n58568, 
      n58569, n58570, n58571, n58572, n58573, n58574, n58575, n58576, n58577, 
      n58578, n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586, 
      n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594, n58595, 
      n58596, n58597, n58598, n58599, n58600, n58601, n58602, n58603, n58604, 
      n58605, n58606, n58607, n58608, n58609, n58610, n58611, n58612, n58613, 
      n58614, n58615, n58616, n58617, n58618, n58619, n58620, n58621, n58622, 
      n58623, n58624, n58625, n58626, n58627, n58628, n58629, n58630, n58631, 
      n58632, n58633, n58634, n58635, n58636, n58637, n58638, n58639, n58640, 
      n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648, n58649, 
      n58650, n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658, 
      n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666, n58667, 
      n58668, n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676, 
      n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685, 
      n58686, n58687, n58688, n58689, n58690, n58691, n58692, n58693, n58694, 
      n58695, n58696, n58697, n58698, n58699, n58700, n58701, n58702, n58703, 
      n58704, n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712, 
      n58713, n58714, n58715, n58716, n58717, n58718, n58719, n58720, n58721, 
      n58722, n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730, 
      n58731, n58732, n58733, n58734, n58735, n58736, n58737, n58738, n58739, 
      n58740, n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748, 
      n58749, n58750, n58751, n58752, n58753, n58754, n58755, n58756, n58757, 
      n58758, n58759, n58760, n58761, n58762, n58763, n58764, n58765, n58766, 
      n58767, n58768, n58769, n58770, n58771, n58772, n58773, n58774, n58775, 
      n58776, n58777, n58778, n58779, n58780, n58781, n58782, n58783, n58784, 
      n58785, n58786, n58787, n58788, n58789, n58790, n58791, n58792, n58793, 
      n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58801, n58802, 
      n58803, n58804, n58805, n58806, n58807, n58808, n58809, n58810, n58811, 
      n58812, n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58820, 
      n58821, n58822, n58823, n58824, n58825, n58826, n58827, n58828, n58829, 
      n58830, n58831, n58832, n58833, n58834, n58835, n58836, n58837, n58838, 
      n58839, n58840, n58841, n58842, n58843, n58844, n58845, n58846, n58847, 
      n58848, n58849, n58850, n58851, n58852, n58853, n58854, n58855, n58856, 
      n58857, n58858, n58859, n58860, n58861, n58862, n58863, n58864, n58865, 
      n58866, n58867, n58868, n58869, n58870, n58871, n58872, n58873, n58874, 
      n58875, n58876, n58877, n58878, n58879, n58880, n58881, n58882, n58883, 
      n58884, n58885, n58886, n58887, n58888, n58889, n58890, n58891, n58892, 
      n58893, n58894, n58895, n58896, n58897, n58898, n58899, n58900, n58901, 
      n58902, n58903, n58904, n58905, n58906, n58907, n58908, n58909, n58910, 
      n58911, n58912, n58913, n58914, n58915, n58916, n58917, n58918, n58919, 
      n58920, n58921, n58922, n58923, n58924, n58925, n58926, n58927, n58928, 
      n58929, n58930, n58931, n58932, n58933, n58934, n58935, n58936, n58937, 
      n58938, n58939, n58940, n58941, n58942, n58943, n58944, n58945, n58946, 
      n58947, n58948, n58949, n58950, n58951, n58952, n58953, n58954, n58955, 
      n58956, n58957, n58958, n58959, n58960, n58961, n58962, n58963, n58964, 
      n58965, n58966, n58967, n58968, n58969, n58970, n58971, n58972, n58973, 
      n58974, n58975, n58976, n58977, n58978, n58979, n58980, n58981, n58982, 
      n58983, n58984, n58985, n58986, n58987, n58988, n58989, n58990, n58991, 
      n58992, n58993, n58994, n58995, n58996, n58997, n58998, n58999, n59000, 
      n59001, n59002, n59003, n59004, n59005, n59006, n59007, n59008, n59009, 
      n59010, n59011, n59012, n59013, n59014, n59015, n59016, n59017, n59018, 
      n59019, n59020, n59021, n59022, n59023, n59024, n59025, n59026, n59027, 
      n59028, n59029, n59030, n59031, n59032, n59033, n59034, n59035, n59036, 
      n59037, n59038, n59039, n59040, n59041, n59042, n59043, n59044, n59045, 
      n59046, n59047, n59048, n59049, n59050, n59051, n59052, n59053, n59054, 
      n59055, n59056, n59057, n59058, n59059, n59060, n59061, n59062, n59063, 
      n59064, n59065, n59066, n59067, n59068, n59069, n59070, n59071, n59072, 
      n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080, n59081, 
      n59082, n59083, n59084, n59085, n59086, n59087, n59088, n59089, n59090, 
      n59091, n59092, n59093, n59094, n59095, n59096, n59097, n59098, n59099, 
      n59100, n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108, 
      n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116, n59117, 
      n59118, n59119, n59120, n59121, n59122, n59123, n59124, n59125, n59126, 
      n59127, n59128, n59129, n59130, n59131, n59132, n59133, n59134, n59135, 
      n59136, n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144, 
      n59145, n59146, n59147, n59148, n59149, n59150, n59151, n59152, n59153, 
      n59154, n59155, n59156, n59157, n59158, n59159, n59160, n59161, n59162, 
      n59163, n59164, n59165, n59166, n59167, n59168, n59169, n59170, n59171, 
      n59172, n59173, n59174, n59175, n59176, n59177, n59178, n59179, n59180, 
      n59181, n59182, n59183, n59184, n59185, n59186, n59187, n59188, n59189, 
      n59190, n59191, n59192, n59193, n59194, n59195, n59196, n59197, n59198, 
      n59199, n59200, n59201, n59202, n59203, n59204, n59205, n59206, n59207, 
      n59208, n59209, n59210, n59211, n59212, n59213, n59214, n59215, n59216, 
      n59217, n59218, n59219, n59220, n59221, n59222, n59223, n59224, n59225, 
      n59226, n59227, n59228, n59229, n59230, n59231, n59232, n59233, n59234, 
      n59235, n59236, n59237, n59238, n59239, n59240, n59241, n59242, n59243, 
      n59244, n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252, 
      n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260, n59261, 
      n59262, n59263, n59264, n59265, n59266, n59267, n59268, n59269, n59270, 
      n59271, n59272, n59273, n59274, n59275, n59276, n59277, n59278, n59279, 
      n59280, n59281, n59282, n59283, n59284, n59285, n59286, n59287, n59288, 
      n59289, n59290, n59291, n59292, n59293, n59294, n59295, n59296, n59297, 
      n59298, n59299, n59300, n59301, n59302, n59303, n59304, n59305, n59306, 
      n59307, n59308, n59309, n59310, n59311, n59312, n59313, n59314, n59315, 
      n59316, n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324, 
      n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332, n59333, 
      n59334, n59335, n59336, n59337, n59338, n59339, n59340, n59341, n59342, 
      n59343, n59344, n59345, n59346, n59347, n59348, n59349, n59350, n59351, 
      n59352, n59353, n59354, n59355, n59356, n59357, n59358, n59359, n59360, 
      n59361, n59362, n59363, n59364, n59365, n59366, n59367, n59368, n59369, 
      n59370, n59371, n59372, n59373, n59374, n59375, n59376, n59377, n59378, 
      n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386, n59387, 
      n59388, n59389, n59390, n59391, n59392, n59393, n59394, n59395, n59396, 
      n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404, n59405, 
      n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413, n59414, 
      n59415, n59416, n59417, n59418, n59419, n59420, n59421, n59422, n59423, 
      n59424, n59425, n59426, n59427, n59428, n59429, n59430, n59431, n59432, 
      n59433, n59434, n59435, n59436, n59437, n59438, n59439, n59440, n59441, 
      n59442, n59443, n59444, n59445, n59446, n59447, n59448, n59449, n59450, 
      n59451, n59452, n59453, n59454, n59455, n59456, n59457, n59458, n59459, 
      n59460, n59461, n59462, n59463, n59464, n59465, n59466, n59467, n59468, 
      n59469, n59470, n59471, n59472, n59473, n59474, n59475, n59476, n59477, 
      n59478, n59479, n59480, n59481, n59482, n59483, n59484, n59485, n59486, 
      n59487, n59488, n59489, n59490, n59491, n59492, n59493, n59494, n59495, 
      n59496, n59497, n59498, n59499, n59500, n59501, n59502, n59503, n59504, 
      n59505, n59506, n59507, n59508, n59509, n59510, n59511, n59512, n59513, 
      n59514, n59515, n59516, n59517, n59518, n59519, n59520, n59521, n59522, 
      n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530, n59531, 
      n59532, n59533, n59534, n59535, n59536, n59537, n59538, n59539, n59540, 
      n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548, n59549, 
      n59550, n59551, n59552, n59553, n59554, n59555, n59556, n59557, n59558, 
      n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566, n59567, 
      n59568, n59569, n59570, n59571, n59572, n59573, n59574, n59575, n59576, 
      n59577, n59578, n59579, n59580, n59581, n59582, n59583, n59584, n59585, 
      n59586, n59587, n59588, n59589, n59590, n59591, n59592, n59593, n59594, 
      n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602, n59603, 
      n59604, n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612, 
      n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620, n59621, 
      n59622, n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630, 
      n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638, n59639, 
      n59640, n59641, n59642, n59643, n59644, n59645, n59646, n59647, n59648, 
      n59649, n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657, 
      n59658, n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666, 
      n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675, 
      n59676, n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684, 
      n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693, 
      n59694, n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702, 
      n59703, n59704, n59705, n59706, n59707, n59708, n59709, n59710, n59711, 
      n59712, n59713, n59714, n59715, n59716, n59717, n59718, n59719, n59720, 
      n59721, n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729, 
      n59730, n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738, 
      n59739, n59740, n59741, n59742, n59743, n59744, n59745, n59746, n59747, 
      n59748, n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756, 
      n59757, n59758, n59759, n59760, n59761, n59762, n59763, n59764, n59765, 
      n59766, n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774, 
      n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59782, n59783, 
      n59784, n59785, n59786, n59787, n59788, n59789, n59790, n59791, n59792, 
      n59793, n59794, n59795, n59796, n59797, n59798, n59799, n59800, n59801, 
      n59802, n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810, 
      n59811, n59812, n59813, n59814, n59815, n59816, n59817, n59818, n59819, 
      n59820, n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828, 
      n59829, n59830, n59831, n59832, n59833, n59834, n59835, n59836, n59837, 
      n59838, n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846, 
      n59847, n59848, n59849, n59850, n59851, n59852, n59853, n59854, n59855, 
      n59856, n59857, n59858, n59859, n59860, n59861, n59862, n59863, n59864, 
      n59865, n59866, n59867, n59868, n59869, n59870, n59871, n59872, n59873, 
      n59874, n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882, 
      n59883, n59884, n59885, n59886, n59887, n59888, n59889, n59890, n59891, 
      n59892, n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900, 
      n59901, n59902, n59903, n59904, n59905, n59906, n59907, n59908, n59909, 
      n59910, n59911, n59912, n59913, n59914, n59915, n59916, n59917, n59918, 
      n59919, n59920, n59921, n59922, n59923, n59924, n59925, n59926, n59927, 
      n59928, n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936, 
      n59937, n59938, n59939, n59940, n59941, n59942, n59943, n59944, n59945, 
      n59946, n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954, 
      n59955, n59956, n59957, n59958, n59959, n59960, n59961, n59962, n59963, 
      n59964, n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972, 
      n59973, n59974, n59975, n59976, n59977, n59978, n59979, n59980, n59981, 
      n59982, n59983, n59984, n59985, n59986, n59987, n59988, n59989, n59990, 
      n59991, n59992, n59993, n59994, n59995, n59996, n59997, n59998, n59999, 
      n60000, n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008, 
      n60009, n60010, n60011, n60012, n60013, n60014, n60015, n60016, n60017, 
      n60018, n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026, 
      n60027, n60028, n60029, n60030, n60031, n60032, n60033, n60034, n60035, 
      n60036, n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044, 
      n60045, n60046, n60047, n60048, n60049, n60050, n60051, n60052, n60053, 
      n60054, n60055, n60056, n60057, n60058, n60059, n60060, n60061, n60062, 
      n60063, n60064, n60065, n60066, n60067, n60068, n60069, n60070, n60071, 
      n60072, n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080, 
      n60081, n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089, 
      n60090, n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098, 
      n60099, n60100, n60101, n60102, n60103, n60104, n60105, n60106, n60107, 
      n60108, n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116, 
      n60117, n60118, n60119, n60120, n60121, n60122, n60123, n60124, n60125, 
      n60126, n60127, n60128, n60129, n60130, n60131, n60132, n60133, n60134, 
      n60135, n60136, n60137, n60138, n60139, n60140, n60141, n60142, n60143, 
      n60144, n60145, n60146, n60147, n60148, n60149, n60150, n60151, n60152, 
      n60153, n60154, n60155, n60156, n60157, n60158, n60159, n60160, n60161, 
      n60162, n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170, 
      n60171, n60172, n60173, n60174, n60175, n60176, n60177, n60178, n60179, 
      n60180, n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188, 
      n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196, n60197, 
      n60198, n60199, n60200, n60201, n60202, n60203, n60204, n60205, n60206, 
      n60207, n60208, n60209, n60210, n60211, n60212, n60213, n60214, n60215, 
      n60216, n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224, 
      n60225, n60226, n60227, n60228, n60229, n60230, n60231, n60232, n60233, 
      n60234, n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242, 
      n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250, n60251, 
      n60252, n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260, 
      n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268, n60269, 
      n60270, n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278, 
      n60279, n60280, n60281, n60282, n60283, n60284, n60285, n60286, n60287, 
      n60288, n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296, 
      n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304, n60305, 
      n60306, n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314, 
      n60315, n60316, n60317, n60318, n60319, n60320, n60321, n60322, n60323, 
      n60324, n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332, 
      n60333, n60334, n60335, n60336, n60337, n60338, n60339, n60340, n60341, 
      n60342, n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350, 
      n60351, n60352, n60353, n60354, n60355, n60356, n60357, n60358, n60359, 
      n60360, n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368, 
      n60369, n60370, n60371, n60372, n60373, n60374, n60375, n60376, n60377, 
      n60378, n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386, 
      n60387, n60388, n60389, n60390, n60391, n60392, n60393, n60394, n60395, 
      n60396, n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404, 
      n60405, n60406, n60407, n60408, n60409, n60410, n60411, n60412, n60413, 
      n60414, n60415, n60416, n60417, n60418, n60419, n60420, n60421, n60422, 
      n60423, n60424, n60425, n60426, n60427, n60428, n60429, n60430, n60431, 
      n60432, n60433, n60434, n60435, n60436, n60437, n60438, n60439, n60440, 
      n60441, n60442, n60443, n60444, n60445, n60446, n60447, n60448, n60449, 
      n60450, n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458, 
      n60459, n60460, n60461, n60462, n60463, n60464, n60465, n60466, n60467, 
      n60468, n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476, 
      n60477, n60478, n60479, n60480, n60481, n60482, n60483, n60484, n60485, 
      n60486, n60487, n60488, n60489, n60490, n60491, n60492, n60493, n60494, 
      n60495, n60496, n60497, n60498, n60499, n60500, n60501, n60502, n60503, 
      n60504, n60505, n60506, n60507, n60508, n60509, n60510, n60511, n60512, 
      n60513, n60514, n60515, n60516, n60517, n60518, n60519, n60520, n60521, 
      n60522, n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530, 
      n60531, n60532, n60533, n60534, n60535, n60536, n60537, n60538, n60539, 
      n60540, n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548, 
      n60549, n60550, n60551, n60552, n60553, n60554, n60555, n60556, n60557, 
      n60558, n60559, n60560, n60561, n60562, n60563, n60564, n60565, n60566, 
      n60567, n60568, n60569, n60570, n60571, n60572, n60573, n60574, n60575, 
      n60576, n60577, n60578, n60579, n60580, n60581, n60582, n60583, n60584, 
      n60585, n60586, n60587, n60588, n60589, n60590, n60591, n60592, n60593, 
      n60594, n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602, 
      n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610, n60611, 
      n60612, n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620, 
      n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628, n60629, 
      n60630, n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638, 
      n60639, n60640, n60641, n60642, n60643, n60644, n60645, n60646, n60647, 
      n60648, n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656, 
      n60657, n60658, n60659, n60660, n60661, n60662, n60663, n60664, n60665, 
      n60666, n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674, 
      n60675, n60676, n60677, n60678, n60679, n60680, n60681, n60682, n60683, 
      n60684, n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692, 
      n60693, n60694, n60695, n60696, n60697, n60698, n60699, n60700, n60701, 
      n60702, n60703, n60704, n60705, n60706, n60707, n60708, n60709, n60710, 
      n60711, n60712, n60713, n60714, n60715, n60716, n60717, n60718, n60719, 
      n60720, n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728, 
      n60729, n60730, n60731, n60732, n60733, n60734, n60735, n60736, n60737, 
      n60738, n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746, 
      n60747, n60748, n60749, n60750, n60751, n60752, n60753, n60754, n60755, 
      n60756, n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764, 
      n60765, n60766, n60767, n60768, n60769, n60770, n60771, n60772, n60773, 
      n60774, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, 
      n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, 
      n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, 
      n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, 
      n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, 
      n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, 
      n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, 
      n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, 
      n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, 
      n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, 
      n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, 
      n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, 
      n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, 
      n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, 
      n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, 
      n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, 
      n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, 
      n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, 
      n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, 
      n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, 
      n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, 
      n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, 
      n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, 
      n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, 
      n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, 
      n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, 
      n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, 
      n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, 
      n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, 
      n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, 
      n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, 
      n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, 
      n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, 
      n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, 
      n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, 
      n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, 
      n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, 
      n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, 
      n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, 
      n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, 
      n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, 
      n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, 
      n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, 
      n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, 
      n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, 
      n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, 
      n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, 
      n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, 
      n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, 
      n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, 
      n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, 
      n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, 
      n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, 
      n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, 
      n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, 
      n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, 
      n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, 
      n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, 
      n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, 
      n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, 
      n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, 
      n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, 
      n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, 
      n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, 
      n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, 
      n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, 
      n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, 
      n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, 
      n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, 
      n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, 
      n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, 
      n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, 
      n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, 
      n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, 
      n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, 
      n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, 
      n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, 
      n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, 
      n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, 
      n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, 
      n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, 
      n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, 
      n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, 
      n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, 
      n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, 
      n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, 
      n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, 
      n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, 
      n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, 
      n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, 
      n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, 
      n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, 
      n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, 
      n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, 
      n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, 
      n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, 
      n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, 
      n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, 
      n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, 
      n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, 
      n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, 
      n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, 
      n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, 
      n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, 
      n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, 
      n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, 
      n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, 
      n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, 
      n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, 
      n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, 
      n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, 
      n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, 
      n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, 
      n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, 
      n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, 
      n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, 
      n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, 
      n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, 
      n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, 
      n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, 
      n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, 
      n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, 
      n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, 
      n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, 
      n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, 
      n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, 
      n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, 
      n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, 
      n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, 
      n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, 
      n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, 
      n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, 
      n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, 
      n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, 
      n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, 
      n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, 
      n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, 
      n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, 
      n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, 
      n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, 
      n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, 
      n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, 
      n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, 
      n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, 
      n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, 
      n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, 
      n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, 
      n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, 
      n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, 
      n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, 
      n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, 
      n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, 
      n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, 
      n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, 
      n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, 
      n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, 
      n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, 
      n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, 
      n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, 
      n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, 
      n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, 
      n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, 
      n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, 
      n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, 
      n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, 
      n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, 
      n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, 
      n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, 
      n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, 
      n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, 
      n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, 
      n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, 
      n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, 
      n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, 
      n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, 
      n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, 
      n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, 
      n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, 
      n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, 
      n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, 
      n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, 
      n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, 
      n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, 
      n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, 
      n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, 
      n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, 
      n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, 
      n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, 
      n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, 
      n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, 
      n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, 
      n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818 : std_logic;

begin
   
   clk_r_REG16701_S5 : DFFR_X1 port map( D => ENABLE, CK => CLK, RN => 
                           RESET_BAR, Q => n53629, QN => n_1554);
   clk_r_REG16748_S2 : DFFR_X1 port map( D => RD1, CK => CLK, RN => RESET_BAR, 
                           Q => n53627, QN => n_1555);
   clk_r_REG16687_S2 : DFFR_X1 port map( D => RD2, CK => CLK, RN => RESET_BAR, 
                           Q => n53626, QN => n_1556);
   clk_r_REG16996_S7 : DFFR_X1 port map( D => ADD_RD1(4), CK => CLK, RN => 
                           RESET_BAR, Q => n53625, QN => n_1557);
   clk_r_REG16998_S7 : DFFS_X1 port map( D => n3558, CK => CLK, SN => RESET_BAR
                           , Q => n_1558, QN => n53624);
   clk_r_REG16931_S7 : DFFR_X1 port map( D => ADD_RD2(4), CK => CLK, RN => 
                           RESET_BAR, Q => n53623, QN => n_1559);
   clk_r_REG16896_S7 : DFFS_X1 port map( D => n3567, CK => CLK, SN => RESET_BAR
                           , Q => n_1560, QN => n53622);
   clk_r_REG13707_S6 : DFFR_X1 port map( D => DATAIN(31), CK => CLK, RN => 
                           RESET_BAR, Q => n53621, QN => n_1561);
   clk_r_REG13700_S8 : DFFR_X1 port map( D => DATAIN(30), CK => CLK, RN => 
                           RESET_BAR, Q => n53620, QN => n_1562);
   clk_r_REG13777_S5 : DFFR_X1 port map( D => DATAIN(29), CK => CLK, RN => 
                           RESET_BAR, Q => n53619, QN => n_1563);
   clk_r_REG13770_S6 : DFFR_X1 port map( D => DATAIN(28), CK => CLK, RN => 
                           RESET_BAR, Q => n53618, QN => n_1564);
   clk_r_REG13763_S5 : DFFR_X1 port map( D => DATAIN(27), CK => CLK, RN => 
                           RESET_BAR, Q => n53617, QN => n_1565);
   clk_r_REG13756_S8 : DFFR_X1 port map( D => DATAIN(26), CK => CLK, RN => 
                           RESET_BAR, Q => n53616, QN => n_1566);
   clk_r_REG13749_S5 : DFFR_X1 port map( D => DATAIN(25), CK => CLK, RN => 
                           RESET_BAR, Q => n53615, QN => n_1567);
   clk_r_REG13740_S5 : DFFR_X1 port map( D => DATAIN(24), CK => CLK, RN => 
                           RESET_BAR, Q => n53614, QN => n_1568);
   clk_r_REG13733_S5 : DFFR_X1 port map( D => DATAIN(23), CK => CLK, RN => 
                           RESET_BAR, Q => n53613, QN => n_1569);
   clk_r_REG13726_S5 : DFFR_X1 port map( D => DATAIN(22), CK => CLK, RN => 
                           RESET_BAR, Q => n53612, QN => n_1570);
   clk_r_REG13719_S5 : DFFR_X1 port map( D => DATAIN(21), CK => CLK, RN => 
                           RESET_BAR, Q => n53611, QN => n_1571);
   clk_r_REG13823_S5 : DFFR_X1 port map( D => DATAIN(20), CK => CLK, RN => 
                           RESET_BAR, Q => n53610, QN => n_1572);
   clk_r_REG13816_S5 : DFFR_X1 port map( D => DATAIN(19), CK => CLK, RN => 
                           RESET_BAR, Q => n53609, QN => n_1573);
   clk_r_REG13809_S5 : DFFR_X1 port map( D => DATAIN(18), CK => CLK, RN => 
                           RESET_BAR, Q => n53608, QN => n_1574);
   clk_r_REG13802_S5 : DFFR_X1 port map( D => DATAIN(17), CK => CLK, RN => 
                           RESET_BAR, Q => n53607, QN => n_1575);
   clk_r_REG13793_S5 : DFFR_X1 port map( D => DATAIN(16), CK => CLK, RN => 
                           RESET_BAR, Q => n53606, QN => n_1576);
   clk_r_REG13916_S11 : DFFR_X1 port map( D => DATAIN(15), CK => CLK, RN => 
                           RESET_BAR, Q => n53605, QN => n_1577);
   clk_r_REG13686_S8 : DFFR_X1 port map( D => DATAIN(14), CK => CLK, RN => 
                           RESET_BAR, Q => n53604, QN => n_1578);
   clk_r_REG13672_S12 : DFFR_X1 port map( D => DATAIN(13), CK => CLK, RN => 
                           RESET_BAR, Q => n53603, QN => n_1579);
   clk_r_REG13903_S11 : DFFR_X1 port map( D => DATAIN(12), CK => CLK, RN => 
                           RESET_BAR, Q => n53602, QN => n_1580);
   clk_r_REG13867_S11 : DFFR_X1 port map( D => DATAIN(11), CK => CLK, RN => 
                           RESET_BAR, Q => n53601, QN => n_1581);
   clk_r_REG13658_S8 : DFFR_X1 port map( D => DATAIN(10), CK => CLK, RN => 
                           RESET_BAR, Q => n53600, QN => n_1582);
   clk_r_REG13848_S11 : DFFR_X1 port map( D => DATAIN(9), CK => CLK, RN => 
                           RESET_BAR, Q => n53599, QN => n_1583);
   clk_r_REG14030_S11 : DFFR_X1 port map( D => DATAIN(8), CK => CLK, RN => 
                           RESET_BAR, Q => n53598, QN => n_1584);
   clk_r_REG14077_S11 : DFFR_X1 port map( D => DATAIN(7), CK => CLK, RN => 
                           RESET_BAR, Q => n53597, QN => n_1585);
   clk_r_REG13835_S5 : DFFR_X1 port map( D => DATAIN(6), CK => CLK, RN => 
                           RESET_BAR, Q => n53596, QN => n_1586);
   clk_r_REG14139_S11 : DFFR_X1 port map( D => DATAIN(5), CK => CLK, RN => 
                           RESET_BAR, Q => n53595, QN => n_1587);
   clk_r_REG14158_S4 : DFFR_X1 port map( D => DATAIN(4), CK => CLK, RN => 
                           RESET_BAR, Q => n53594, QN => n_1588);
   clk_r_REG14118_S5 : DFFR_X1 port map( D => DATAIN(3), CK => CLK, RN => 
                           RESET_BAR, Q => n53593, QN => n_1589);
   clk_r_REG14064_S5 : DFFR_X1 port map( D => DATAIN(2), CK => CLK, RN => 
                           RESET_BAR, Q => n53592, QN => n_1590);
   clk_r_REG14009_S5 : DFFR_X1 port map( D => DATAIN(1), CK => CLK, RN => 
                           RESET_BAR, Q => n53591, QN => n_1591);
   clk_r_REG13647_S11 : DFFR_X1 port map( D => DATAIN(0), CK => CLK, RN => 
                           RESET_BAR, Q => n53590, QN => n_1592);
   clk_r_REG16916_S7 : DFFR_X1 port map( D => n40589, CK => CLK, RN => 
                           RESET_BAR, Q => n53589, QN => n_1593);
   clk_r_REG16914_S7 : DFFR_X1 port map( D => n40588, CK => CLK, RN => 
                           RESET_BAR, Q => n53588, QN => n_1594);
   clk_r_REG16912_S7 : DFFR_X1 port map( D => n49092, CK => CLK, RN => 
                           RESET_BAR, Q => n53587, QN => n_1595);
   clk_r_REG16928_S7 : DFFR_X1 port map( D => n47429, CK => CLK, RN => 
                           RESET_BAR, Q => n53586, QN => n_1596);
   clk_r_REG16924_S7 : DFFR_X1 port map( D => n49090, CK => CLK, RN => 
                           RESET_BAR, Q => n53585, QN => n_1597);
   clk_r_REG16948_S7 : DFFS_X1 port map( D => n3568, CK => CLK, SN => RESET_BAR
                           , Q => n53584, QN => n_1598);
   clk_r_REG16954_S7 : DFFR_X1 port map( D => n41691, CK => CLK, RN => 
                           RESET_BAR, Q => n53583, QN => n_1599);
   clk_r_REG16957_S7 : DFFR_X1 port map( D => n3571, CK => CLK, RN => RESET_BAR
                           , Q => n53582, QN => n_1600);
   clk_r_REG16941_S7 : DFFR_X1 port map( D => n3570, CK => CLK, RN => RESET_BAR
                           , Q => n53581, QN => n_1601);
   clk_r_REG16938_S7 : DFFR_X1 port map( D => n3569, CK => CLK, RN => RESET_BAR
                           , Q => n53580, QN => n_1602);
   clk_r_REG16936_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR
                           , Q => n53578, QN => n_1603);
   clk_r_REG16945_S7 : DFFR_X1 port map( D => n3574, CK => CLK, RN => RESET_BAR
                           , Q => n53577, QN => n_1604);
   clk_r_REG16902_S7 : DFFR_X1 port map( D => n49088, CK => CLK, RN => 
                           RESET_BAR, Q => n53576, QN => n_1605);
   clk_r_REG16900_S7 : DFFR_X1 port map( D => n47428, CK => CLK, RN => 
                           RESET_BAR, Q => n53575, QN => n_1606);
   clk_r_REG16908_S7 : DFFR_X1 port map( D => n49094, CK => CLK, RN => 
                           RESET_BAR, Q => n53574, QN => n_1607);
   clk_r_REG16906_S7 : DFFR_X1 port map( D => n49089, CK => CLK, RN => 
                           RESET_BAR, Q => n53573, QN => n_1608);
   clk_r_REG16922_S7 : DFFR_X1 port map( D => n49086, CK => CLK, RN => 
                           RESET_BAR, Q => n53572, QN => n_1609);
   clk_r_REG16935_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR
                           , Q => n53571, QN => n_1610);
   clk_r_REG16956_S7 : DFFR_X1 port map( D => n3571, CK => CLK, RN => RESET_BAR
                           , Q => n53570, QN => n_1611);
   clk_r_REG16904_S7 : DFFR_X1 port map( D => n49091, CK => CLK, RN => 
                           RESET_BAR, Q => n53569, QN => n_1612);
   clk_r_REG16898_S7 : DFFR_X1 port map( D => n40592, CK => CLK, RN => 
                           RESET_BAR, Q => n53568, QN => n_1613);
   clk_r_REG16918_S7 : DFFR_X1 port map( D => n49085, CK => CLK, RN => 
                           RESET_BAR, Q => n53567, QN => n_1614);
   clk_r_REG16947_S7 : DFFS_X1 port map( D => n3568, CK => CLK, SN => RESET_BAR
                           , Q => n53565, QN => n_1615);
   clk_r_REG16920_S7 : DFFR_X1 port map( D => n40591, CK => CLK, RN => 
                           RESET_BAR, Q => n53564, QN => n_1616);
   clk_r_REG16926_S7 : DFFR_X1 port map( D => n49087, CK => CLK, RN => 
                           RESET_BAR, Q => n53563, QN => n_1617);
   clk_r_REG16944_S7 : DFFR_X1 port map( D => n3574, CK => CLK, RN => RESET_BAR
                           , Q => n53562, QN => n_1618);
   clk_r_REG16910_S7 : DFFR_X1 port map( D => n49093, CK => CLK, RN => 
                           RESET_BAR, Q => n53561, QN => n_1619);
   clk_r_REG16950_S7 : DFFR_X1 port map( D => n3573, CK => CLK, RN => RESET_BAR
                           , Q => n53560, QN => n_1620);
   clk_r_REG16951_S7 : DFFR_X1 port map( D => n3573, CK => CLK, RN => RESET_BAR
                           , Q => n53559, QN => n_1621);
   clk_r_REG16883_S7 : DFFR_X1 port map( D => n40581, CK => CLK, RN => 
                           RESET_BAR, Q => n53558, QN => n_1622);
   clk_r_REG16876_S7 : DFFR_X1 port map( D => n40582, CK => CLK, RN => 
                           RESET_BAR, Q => n53557, QN => n_1623);
   clk_r_REG16866_S7 : DFFR_X1 port map( D => n40576, CK => CLK, RN => 
                           RESET_BAR, Q => n53556, QN => n_1624);
   clk_r_REG16888_S7 : DFFR_X1 port map( D => n40585, CK => CLK, RN => 
                           RESET_BAR, Q => n53555, QN => n_1625);
   clk_r_REG16881_S7 : DFFR_X1 port map( D => n40574, CK => CLK, RN => 
                           RESET_BAR, Q => n53554, QN => n_1626);
   clk_r_REG16846_S7 : DFFR_X1 port map( D => n47431, CK => CLK, RN => 
                           RESET_BAR, Q => n53553, QN => n_1627);
   clk_r_REG16868_S7 : DFFR_X1 port map( D => n40577, CK => CLK, RN => 
                           RESET_BAR, Q => n53552, QN => n_1628);
   clk_r_REG16864_S7 : DFFR_X1 port map( D => n41692, CK => CLK, RN => 
                           RESET_BAR, Q => n53551, QN => n_1629);
   clk_r_REG16870_S7 : DFFR_X1 port map( D => n3560, CK => CLK, RN => RESET_BAR
                           , Q => n53550, QN => n_1630);
   clk_r_REG16885_S7 : DFFR_X1 port map( D => n41689, CK => CLK, RN => 
                           RESET_BAR, Q => n53549, QN => n_1631);
   clk_r_REG16842_S7 : DFFR_X1 port map( D => n3566, CK => CLK, RN => RESET_BAR
                           , Q => n53548, QN => n_1632);
   clk_r_REG16857_S7 : DFFR_X1 port map( D => n41686, CK => CLK, RN => 
                           RESET_BAR, Q => n53546, QN => n_1633);
   clk_r_REG16860_S7 : DFFR_X1 port map( D => n49097, CK => CLK, RN => 
                           RESET_BAR, Q => n53545, QN => n_1634);
   clk_r_REG16838_S7 : DFFR_X1 port map( D => n49095, CK => CLK, RN => 
                           RESET_BAR, Q => n53544, QN => n_1635);
   clk_r_REG16855_S7 : DFFR_X1 port map( D => n40584, CK => CLK, RN => 
                           RESET_BAR, Q => n53543, QN => n_1636);
   clk_r_REG16840_S7 : DFFR_X1 port map( D => n40586, CK => CLK, RN => 
                           RESET_BAR, Q => n53542, QN => n_1637);
   clk_r_REG16850_S7 : DFFR_X1 port map( D => n41687, CK => CLK, RN => 
                           RESET_BAR, Q => n53541, QN => n_1638);
   clk_r_REG16878_S7 : DFFR_X1 port map( D => n41688, CK => CLK, RN => 
                           RESET_BAR, Q => n53540, QN => n_1639);
   clk_r_REG16892_S7 : DFFS_X1 port map( D => n41690, CK => CLK, SN => 
                           RESET_BAR, Q => n53539, QN => n_1640);
   clk_r_REG16871_S7 : DFFR_X1 port map( D => n3560, CK => CLK, RN => RESET_BAR
                           , Q => n53538, QN => n_1641);
   clk_r_REG16890_S7 : DFFR_X1 port map( D => n40587, CK => CLK, RN => 
                           RESET_BAR, Q => n53537, QN => n_1642);
   clk_r_REG16853_S7 : DFFR_X1 port map( D => n40580, CK => CLK, RN => 
                           RESET_BAR, Q => n53536, QN => n_1643);
   clk_r_REG16848_S7 : DFFR_X1 port map( D => n49096, CK => CLK, RN => 
                           RESET_BAR, Q => n53535, QN => n_1644);
   clk_r_REG16874_S7 : DFFR_X1 port map( D => n47430, CK => CLK, RN => 
                           RESET_BAR, Q => n53534, QN => n_1645);
   clk_r_REG16862_S7 : DFFR_X1 port map( D => n40583, CK => CLK, RN => 
                           RESET_BAR, Q => n53533, QN => n_1646);
   clk_r_REG16783_S3 : DFFS_X1 port map( D => n58169, CK => CLK, SN => 
                           RESET_BAR, Q => n_1647, QN => n58166);
   clk_r_REG16784_S4 : DFFR_X1 port map( D => n58166, CK => CLK, RN => 
                           RESET_BAR, Q => n_1648, QN => n53531);
   clk_r_REG16785_S4 : DFFR_X1 port map( D => n58166, CK => CLK, RN => 
                           RESET_BAR, Q => n53530, QN => n_1649);
   clk_r_REG15349_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n53529, QN 
                           => n_1650);
   clk_r_REG16856_S7 : DFFR_X1 port map( D => n41686, CK => CLK, RN => 
                           RESET_BAR, Q => n53528, QN => n_1651);
   clk_r_REG16849_S7 : DFFR_X1 port map( D => n41687, CK => CLK, RN => 
                           RESET_BAR, Q => n53527, QN => n_1652);
   clk_r_REG16877_S7 : DFFR_X1 port map( D => n41688, CK => CLK, RN => 
                           RESET_BAR, Q => n53526, QN => n_1653);
   clk_r_REG16891_S7 : DFFS_X1 port map( D => n41690, CK => CLK, SN => 
                           RESET_BAR, Q => n53525, QN => n_1654);
   clk_r_REG16884_S7 : DFFR_X1 port map( D => n41689, CK => CLK, RN => 
                           RESET_BAR, Q => n53524, QN => n_1655);
   clk_r_REG16953_S7 : DFFR_X1 port map( D => n41691, CK => CLK, RN => 
                           RESET_BAR, Q => n53523, QN => n_1656);
   clk_r_REG16863_S7 : DFFR_X1 port map( D => n41692, CK => CLK, RN => 
                           RESET_BAR, Q => n53522, QN => n_1657);
   clk_r_REG16649_S1 : DFF_X1 port map( D => n3541, CK => CLK, Q => n53521, QN 
                           => n_1658);
   clk_r_REG16955_S7 : DFFR_X1 port map( D => n3571, CK => CLK, RN => RESET_BAR
                           , Q => n53520, QN => n_1659);
   clk_r_REG16949_S7 : DFFR_X1 port map( D => n3573, CK => CLK, RN => RESET_BAR
                           , Q => n53519, QN => n_1660);
   clk_r_REG16869_S7 : DFFR_X1 port map( D => n3560, CK => CLK, RN => RESET_BAR
                           , Q => n53518, QN => n_1661);
   clk_r_REG16841_S7 : DFFR_X1 port map( D => n3566, CK => CLK, RN => RESET_BAR
                           , Q => n53517, QN => n_1662);
   clk_r_REG16946_S7 : DFFS_X1 port map( D => n3568, CK => CLK, SN => RESET_BAR
                           , Q => n53516, QN => n_1663);
   clk_r_REG16940_S7 : DFFR_X1 port map( D => n3570, CK => CLK, RN => RESET_BAR
                           , Q => n53515, QN => n_1664);
   clk_r_REG16934_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR
                           , Q => n53514, QN => n_1665);
   clk_r_REG16943_S7 : DFFR_X1 port map( D => n3574, CK => CLK, RN => RESET_BAR
                           , Q => n53513, QN => n_1666);
   clk_r_REG16937_S7 : DFFR_X1 port map( D => n3569, CK => CLK, RN => RESET_BAR
                           , Q => n53512, QN => n_1667);
   clk_r_REG16789_S4 : DFFR_X1 port map( D => n58167, CK => CLK, RN => 
                           RESET_BAR, Q => n53511, QN => n_1668);
   clk_r_REG16787_S3 : DFFS_X1 port map( D => n58168, CK => CLK, SN => 
                           RESET_BAR, Q => n_1669, QN => n58167);
   clk_r_REG16788_S4 : DFFR_X1 port map( D => n58167, CK => CLK, RN => 
                           RESET_BAR, Q => n_1670, QN => n53509);
   clk_r_REG16786_S2 : DFFR_X1 port map( D => ADD_WR(4), CK => CLK, RN => 
                           RESET_BAR, Q => n_1671, QN => n58168);
   clk_r_REG16782_S2 : DFFR_X1 port map( D => ADD_WR(3), CK => CLK, RN => 
                           RESET_BAR, Q => n_1672, QN => n58169);
   clk_r_REG15989_S1 : DFF_X1 port map( D => n2735, CK => CLK, Q => n53506, QN 
                           => n_1673);
   clk_r_REG15861_S1 : DFF_X1 port map( D => n2671, CK => CLK, Q => n53505, QN 
                           => n_1674);
   clk_r_REG15733_S1 : DFF_X1 port map( D => n2607, CK => CLK, Q => n53504, QN 
                           => n_1675);
   clk_r_REG16053_S1 : DFF_X1 port map( D => n2767, CK => CLK, Q => n53503, QN 
                           => n_1676);
   clk_r_REG15797_S1 : DFF_X1 port map( D => n2639, CK => CLK, Q => n53502, QN 
                           => n_1677);
   clk_r_REG16055_S1 : DFF_X1 port map( D => n2766, CK => CLK, Q => n53501, QN 
                           => n_1678);
   clk_r_REG16308_S1 : DFF_X1 port map( D => n2543, CK => CLK, Q => n53500, QN 
                           => n_1679);
   clk_r_REG16310_S1 : DFF_X1 port map( D => n2542, CK => CLK, Q => n53499, QN 
                           => n_1680);
   clk_r_REG16372_S1 : DFF_X1 port map( D => n2575, CK => CLK, Q => n53498, QN 
                           => n_1681);
   clk_r_REG15799_S1 : DFF_X1 port map( D => n2638, CK => CLK, Q => n53497, QN 
                           => n_1682);
   clk_r_REG15991_S1 : DFF_X1 port map( D => n2734, CK => CLK, Q => n53496, QN 
                           => n_1683);
   clk_r_REG15993_S1 : DFF_X1 port map( D => n2733, CK => CLK, Q => n53495, QN 
                           => n_1684);
   clk_r_REG15995_S1 : DFF_X1 port map( D => n2732, CK => CLK, Q => n53494, QN 
                           => n_1685);
   clk_r_REG15863_S1 : DFF_X1 port map( D => n2670, CK => CLK, Q => n53493, QN 
                           => n_1686);
   clk_r_REG16057_S1 : DFF_X1 port map( D => n2765, CK => CLK, Q => n53492, QN 
                           => n_1687);
   clk_r_REG15801_S1 : DFF_X1 port map( D => n2637, CK => CLK, Q => n53491, QN 
                           => n_1688);
   clk_r_REG16059_S1 : DFF_X1 port map( D => n2764, CK => CLK, Q => n53490, QN 
                           => n_1689);
   clk_r_REG16374_S1 : DFF_X1 port map( D => n2574, CK => CLK, Q => n53489, QN 
                           => n_1690);
   clk_r_REG16376_S1 : DFF_X1 port map( D => n2573, CK => CLK, Q => n53488, QN 
                           => n_1691);
   clk_r_REG15891_S1 : DFF_X1 port map( D => n2694, CK => CLK, Q => n53487, QN 
                           => n_1692);
   clk_r_REG16061_S1 : DFF_X1 port map( D => n2763, CK => CLK, Q => n53486, QN 
                           => n_1693);
   clk_r_REG15865_S1 : DFF_X1 port map( D => n2669, CK => CLK, Q => n53485, QN 
                           => n_1694);
   clk_r_REG15997_S1 : DFF_X1 port map( D => n2731, CK => CLK, Q => n53484, QN 
                           => n_1695);
   clk_r_REG16312_S1 : DFF_X1 port map( D => n2541, CK => CLK, Q => n53483, QN 
                           => n_1696);
   clk_r_REG15893_S1 : DFF_X1 port map( D => n2695, CK => CLK, Q => n53482, QN 
                           => n_1697);
   clk_r_REG16314_S1 : DFF_X1 port map( D => n2540, CK => CLK, Q => n53481, QN 
                           => n_1698);
   clk_r_REG16316_S1 : DFF_X1 port map( D => n2539, CK => CLK, Q => n53480, QN 
                           => n_1699);
   clk_r_REG16063_S1 : DFF_X1 port map( D => n2762, CK => CLK, Q => n53479, QN 
                           => n_1700);
   clk_r_REG15735_S1 : DFF_X1 port map( D => n2606, CK => CLK, Q => n53478, QN 
                           => n_1701);
   clk_r_REG15999_S1 : DFF_X1 port map( D => n2730, CK => CLK, Q => n53477, QN 
                           => n_1702);
   clk_r_REG16318_S1 : DFF_X1 port map( D => n2538, CK => CLK, Q => n53476, QN 
                           => n_1703);
   clk_r_REG16320_S1 : DFF_X1 port map( D => n2537, CK => CLK, Q => n53475, QN 
                           => n_1704);
   clk_r_REG16065_S1 : DFF_X1 port map( D => n2761, CK => CLK, Q => n53474, QN 
                           => n_1705);
   clk_r_REG16001_S1 : DFF_X1 port map( D => n2729, CK => CLK, Q => n53473, QN 
                           => n_1706);
   clk_r_REG16003_S1 : DFF_X1 port map( D => n2728, CK => CLK, Q => n53472, QN 
                           => n_1707);
   clk_r_REG15895_S1 : DFF_X1 port map( D => n2696, CK => CLK, Q => n53471, QN 
                           => n_1708);
   clk_r_REG15737_S1 : DFF_X1 port map( D => n2605, CK => CLK, Q => n53470, QN 
                           => n_1709);
   clk_r_REG15897_S1 : DFF_X1 port map( D => n2697, CK => CLK, Q => n53469, QN 
                           => n_1710);
   clk_r_REG15867_S1 : DFF_X1 port map( D => n2668, CK => CLK, Q => n53468, QN 
                           => n_1711);
   clk_r_REG15899_S1 : DFF_X1 port map( D => n2698, CK => CLK, Q => n53467, QN 
                           => n_1712);
   clk_r_REG15803_S1 : DFF_X1 port map( D => n2636, CK => CLK, Q => n53466, QN 
                           => n_1713);
   clk_r_REG16322_S1 : DFF_X1 port map( D => n2536, CK => CLK, Q => n53465, QN 
                           => n_1714);
   clk_r_REG15739_S1 : DFF_X1 port map( D => n2604, CK => CLK, Q => n53464, QN 
                           => n_1715);
   clk_r_REG16378_S1 : DFF_X1 port map( D => n2572, CK => CLK, Q => n53463, QN 
                           => n_1716);
   clk_r_REG16067_S1 : DFF_X1 port map( D => n2760, CK => CLK, Q => n53462, QN 
                           => n_1717);
   clk_r_REG13709_S1 : DFF_X1 port map( D => n2565, CK => CLK, Q => n53461, QN 
                           => n_1718);
   clk_r_REG15869_S1 : DFF_X1 port map( D => n2667, CK => CLK, Q => n53460, QN 
                           => n_1719);
   clk_r_REG16380_S1 : DFF_X1 port map( D => n2571, CK => CLK, Q => n53459, QN 
                           => n_1720);
   clk_r_REG13751_S1 : DFF_X1 port map( D => n2757, CK => CLK, Q => n53458, QN 
                           => n_1721);
   clk_r_REG16382_S1 : DFF_X1 port map( D => n2570, CK => CLK, Q => n53457, QN 
                           => n_1722);
   clk_r_REG16384_S1 : DFF_X1 port map( D => n2569, CK => CLK, Q => n53456, QN 
                           => n_1723);
   clk_r_REG15805_S1 : DFF_X1 port map( D => n2635, CK => CLK, Q => n53455, QN 
                           => n_1724);
   clk_r_REG15871_S1 : DFF_X1 port map( D => n2666, CK => CLK, Q => n53454, QN 
                           => n_1725);
   clk_r_REG15873_S1 : DFF_X1 port map( D => n2665, CK => CLK, Q => n53453, QN 
                           => n_1726);
   clk_r_REG15807_S1 : DFF_X1 port map( D => n2634, CK => CLK, Q => n53452, QN 
                           => n_1727);
   clk_r_REG15809_S1 : DFF_X1 port map( D => n2633, CK => CLK, Q => n53451, QN 
                           => n_1728);
   clk_r_REG16386_S1 : DFF_X1 port map( D => n2568, CK => CLK, Q => n53450, QN 
                           => n_1729);
   clk_r_REG13702_S1 : DFF_X1 port map( D => n2597, CK => CLK, Q => n53449, QN 
                           => n_1730);
   clk_r_REG15875_S1 : DFF_X1 port map( D => n2664, CK => CLK, Q => n53448, QN 
                           => n_1731);
   clk_r_REG13765_S1 : DFF_X1 port map( D => n2693, CK => CLK, Q => n53447, QN 
                           => n_1732);
   clk_r_REG15741_S1 : DFF_X1 port map( D => n2603, CK => CLK, Q => n53446, QN 
                           => n_1733);
   clk_r_REG15901_S1 : DFF_X1 port map( D => n2699, CK => CLK, Q => n53445, QN 
                           => n_1734);
   clk_r_REG15811_S1 : DFF_X1 port map( D => n2632, CK => CLK, Q => n53444, QN 
                           => n_1735);
   clk_r_REG15903_S1 : DFF_X1 port map( D => n2700, CK => CLK, Q => n53443, QN 
                           => n_1736);
   clk_r_REG13772_S1 : DFF_X1 port map( D => n2661, CK => CLK, Q => n53442, QN 
                           => n_1737);
   clk_r_REG15905_S1 : DFF_X1 port map( D => n2701, CK => CLK, Q => n53441, QN 
                           => n_1738);
   clk_r_REG13758_S1 : DFF_X1 port map( D => n2725, CK => CLK, Q => n53440, QN 
                           => n_1739);
   clk_r_REG15743_S1 : DFF_X1 port map( D => n2602, CK => CLK, Q => n53439, QN 
                           => n_1740);
   clk_r_REG15745_S1 : DFF_X1 port map( D => n2601, CK => CLK, Q => n53438, QN 
                           => n_1741);
   clk_r_REG15747_S1 : DFF_X1 port map( D => n2600, CK => CLK, Q => n53437, QN 
                           => n_1742);
   clk_r_REG13779_S1 : DFF_X1 port map( D => n2629, CK => CLK, Q => n53436, QN 
                           => n_1743);
   clk_r_REG13742_S1 : DFF_X1 port map( D => n2789, CK => CLK, Q => n53435, QN 
                           => n_1744);
   clk_r_REG16330_S1 : DFF_X1 port map( D => n2596, CK => CLK, Q => n53434, QN 
                           => n_1745);
   clk_r_REG15947_S1 : DFF_X1 port map( D => n2756, CK => CLK, Q => n53433, QN 
                           => n_1746);
   clk_r_REG15819_S1 : DFF_X1 port map( D => n2692, CK => CLK, Q => n53432, QN 
                           => n_1747);
   clk_r_REG15821_S1 : DFF_X1 port map( D => n2691, CK => CLK, Q => n53431, QN 
                           => n_1748);
   clk_r_REG15949_S1 : DFF_X1 port map( D => n2755, CK => CLK, Q => n53430, QN 
                           => n_1749);
   clk_r_REG16332_S1 : DFF_X1 port map( D => n2595, CK => CLK, Q => n53429, QN 
                           => n_1750);
   clk_r_REG15755_S1 : DFF_X1 port map( D => n2660, CK => CLK, Q => n53428, QN 
                           => n_1751);
   clk_r_REG16011_S1 : DFF_X1 port map( D => n2788, CK => CLK, Q => n53427, QN 
                           => n_1752);
   clk_r_REG16334_S1 : DFF_X1 port map( D => n2594, CK => CLK, Q => n53426, QN 
                           => n_1753);
   clk_r_REG16180_S1 : DFF_X1 port map( D => n2832, CK => CLK, Q => n53425, QN 
                           => n_1754);
   clk_r_REG16336_S1 : DFF_X1 port map( D => n2593, CK => CLK, Q => n53424, QN 
                           => n_1755);
   clk_r_REG15757_S1 : DFF_X1 port map( D => n2659, CK => CLK, Q => n53423, QN 
                           => n_1756);
   clk_r_REG15759_S1 : DFF_X1 port map( D => n2658, CK => CLK, Q => n53422, QN 
                           => n_1757);
   clk_r_REG15157_S1 : DFF_X1 port map( D => n3152, CK => CLK, Q => n53421, QN 
                           => n_1758);
   clk_r_REG15761_S1 : DFF_X1 port map( D => n2657, CK => CLK, Q => n53420, QN 
                           => n_1759);
   clk_r_REG15823_S1 : DFF_X1 port map( D => n2690, CK => CLK, Q => n53419, QN 
                           => n_1760);
   clk_r_REG16266_S1 : DFF_X1 port map( D => n2564, CK => CLK, Q => n53418, QN 
                           => n_1761);
   clk_r_REG15825_S1 : DFF_X1 port map( D => n2689, CK => CLK, Q => n53417, QN 
                           => n_1762);
   clk_r_REG15813_S1 : DFF_X1 port map( D => n2631, CK => CLK, Q => n53416, QN 
                           => n_1763);
   clk_r_REG16268_S1 : DFF_X1 port map( D => n2563, CK => CLK, Q => n53415, QN 
                           => n_1764);
   clk_r_REG15951_S1 : DFF_X1 port map( D => n2754, CK => CLK, Q => n53414, QN 
                           => n_1765);
   clk_r_REG15883_S1 : DFF_X1 port map( D => n2724, CK => CLK, Q => n53413, QN 
                           => n_1766);
   clk_r_REG15885_S1 : DFF_X1 port map( D => n2723, CK => CLK, Q => n53412, QN 
                           => n_1767);
   clk_r_REG15691_S1 : DFF_X1 port map( D => n2628, CK => CLK, Q => n53411, QN 
                           => n_1768);
   clk_r_REG15693_S1 : DFF_X1 port map( D => n2627, CK => CLK, Q => n53410, QN 
                           => n_1769);
   clk_r_REG16388_S1 : DFF_X1 port map( D => n2567, CK => CLK, Q => n53409, QN 
                           => n_1770);
   clk_r_REG16390_S1 : DFF_X1 port map( D => n2566, CK => CLK, Q => n53408, QN 
                           => n_1771);
   clk_r_REG16338_S1 : DFF_X1 port map( D => n2592, CK => CLK, Q => n53407, QN 
                           => n_1772);
   clk_r_REG16270_S1 : DFF_X1 port map( D => n2562, CK => CLK, Q => n53406, QN 
                           => n_1773);
   clk_r_REG16272_S1 : DFF_X1 port map( D => n2561, CK => CLK, Q => n53405, QN 
                           => n_1774);
   clk_r_REG15887_S1 : DFF_X1 port map( D => n2722, CK => CLK, Q => n53404, QN 
                           => n_1775);
   clk_r_REG15889_S1 : DFF_X1 port map( D => n2721, CK => CLK, Q => n53403, QN 
                           => n_1776);
   clk_r_REG15953_S1 : DFF_X1 port map( D => n2753, CK => CLK, Q => n53402, QN 
                           => n_1777);
   clk_r_REG15877_S1 : DFF_X1 port map( D => n2663, CK => CLK, Q => n53401, QN 
                           => n_1778);
   clk_r_REG16324_S1 : DFF_X1 port map( D => n2535, CK => CLK, Q => n53400, QN 
                           => n_1779);
   clk_r_REG16005_S1 : DFF_X1 port map( D => n2727, CK => CLK, Q => n53399, QN 
                           => n_1780);
   clk_r_REG15695_S1 : DFF_X1 port map( D => n2626, CK => CLK, Q => n53398, QN 
                           => n_1781);
   clk_r_REG16013_S1 : DFF_X1 port map( D => n2787, CK => CLK, Q => n53397, QN 
                           => n_1782);
   clk_r_REG15879_S1 : DFF_X1 port map( D => n2662, CK => CLK, Q => n53396, QN 
                           => n_1783);
   clk_r_REG15907_S1 : DFF_X1 port map( D => n2702, CK => CLK, Q => n53395, QN 
                           => n_1784);
   clk_r_REG15159_S1 : DFF_X1 port map( D => n3151, CK => CLK, Q => n53394, QN 
                           => n_1785);
   clk_r_REG16007_S1 : DFF_X1 port map( D => n2726, CK => CLK, Q => n53393, QN 
                           => n_1786);
   clk_r_REG16326_S1 : DFF_X1 port map( D => n2534, CK => CLK, Q => n53392, QN 
                           => n_1787);
   clk_r_REG15827_S1 : DFF_X1 port map( D => n2688, CK => CLK, Q => n53391, QN 
                           => n_1788);
   clk_r_REG16116_S1 : DFF_X1 port map( D => n2800, CK => CLK, Q => n53390, QN 
                           => n_1789);
   clk_r_REG16118_S1 : DFF_X1 port map( D => n2799, CK => CLK, Q => n53389, QN 
                           => n_1790);
   clk_r_REG16434_S1 : DFF_X1 port map( D => n3088, CK => CLK, Q => n53388, QN 
                           => n_1791);
   clk_r_REG16436_S1 : DFF_X1 port map( D => n3087, CK => CLK, Q => n53387, QN 
                           => n_1792);
   clk_r_REG16015_S1 : DFF_X1 port map( D => n2786, CK => CLK, Q => n53386, QN 
                           => n_1793);
   clk_r_REG15909_S1 : DFF_X1 port map( D => n2703, CK => CLK, Q => n53385, QN 
                           => n_1794);
   clk_r_REG15697_S1 : DFF_X1 port map( D => n2625, CK => CLK, Q => n53384, QN 
                           => n_1795);
   clk_r_REG15955_S1 : DFF_X1 port map( D => n2752, CK => CLK, Q => n53383, QN 
                           => n_1796);
   clk_r_REG15911_S1 : DFF_X1 port map( D => n2720, CK => CLK, Q => n53382, QN 
                           => n_1797);
   clk_r_REG15699_S1 : DFF_X1 port map( D => n2624, CK => CLK, Q => n53381, QN 
                           => n_1798);
   clk_r_REG15749_S1 : DFF_X1 port map( D => n2599, CK => CLK, Q => n53380, QN 
                           => n_1799);
   clk_r_REG15913_S1 : DFF_X1 port map( D => n2719, CK => CLK, Q => n53379, QN 
                           => n_1800);
   clk_r_REG15751_S1 : DFF_X1 port map( D => n2598, CK => CLK, Q => n53378, QN 
                           => n_1801);
   clk_r_REG16274_S1 : DFF_X1 port map( D => n2560, CK => CLK, Q => n53377, QN 
                           => n_1802);
   clk_r_REG15829_S1 : DFF_X1 port map( D => n2687, CK => CLK, Q => n53376, QN 
                           => n_1803);
   clk_r_REG16182_S1 : DFF_X1 port map( D => n2831, CK => CLK, Q => n53375, QN 
                           => n_1804);
   clk_r_REG16340_S1 : DFF_X1 port map( D => n2591, CK => CLK, Q => n53374, QN 
                           => n_1805);
   clk_r_REG15701_S1 : DFF_X1 port map( D => n2623, CK => CLK, Q => n53373, QN 
                           => n_1806);
   clk_r_REG16120_S1 : DFF_X1 port map( D => n2798, CK => CLK, Q => n53372, QN 
                           => n_1807);
   clk_r_REG16017_S1 : DFF_X1 port map( D => n2785, CK => CLK, Q => n53371, QN 
                           => n_1808);
   clk_r_REG16184_S1 : DFF_X1 port map( D => n2830, CK => CLK, Q => n53370, QN 
                           => n_1809);
   clk_r_REG16019_S1 : DFF_X1 port map( D => n2784, CK => CLK, Q => n53369, QN 
                           => n_1810);
   clk_r_REG15957_S1 : DFF_X1 port map( D => n2751, CK => CLK, Q => n53368, QN 
                           => n_1811);
   clk_r_REG15763_S1 : DFF_X1 port map( D => n2656, CK => CLK, Q => n53367, QN 
                           => n_1812);
   clk_r_REG16069_S1 : DFF_X1 port map( D => n2759, CK => CLK, Q => n53366, QN 
                           => n_1813);
   clk_r_REG15765_S1 : DFF_X1 port map( D => n2655, CK => CLK, Q => n53365, QN 
                           => n_1814);
   clk_r_REG15815_S1 : DFF_X1 port map( D => n2630, CK => CLK, Q => n53364, QN 
                           => n_1815);
   clk_r_REG16071_S1 : DFF_X1 port map( D => n2758, CK => CLK, Q => n53363, QN 
                           => n_1816);
   clk_r_REG15447_S1 : DFF_X1 port map( D => n2918, CK => CLK, Q => n53362, QN 
                           => n_1817);
   clk_r_REG16244_S1 : DFF_X1 port map( D => n2864, CK => CLK, Q => n53361, QN 
                           => n_1818);
   clk_r_REG16499_S1 : DFF_X1 port map( D => n3120, CK => CLK, Q => n53360, QN 
                           => n_1819);
   clk_r_REG16276_S1 : DFF_X1 port map( D => n2559, CK => CLK, Q => n53359, QN 
                           => n_1820);
   clk_r_REG15449_S1 : DFF_X1 port map( D => n2919, CK => CLK, Q => n53358, QN 
                           => n_1821);
   clk_r_REG15161_S1 : DFF_X1 port map( D => n3150, CK => CLK, Q => n53357, QN 
                           => n_1822);
   clk_r_REG15451_S1 : DFF_X1 port map( D => n2920, CK => CLK, Q => n53356, QN 
                           => n_1823);
   clk_r_REG16021_S1 : DFF_X1 port map( D => n2783, CK => CLK, Q => n53355, QN 
                           => n_1824);
   clk_r_REG15453_S1 : DFF_X1 port map( D => n2921, CK => CLK, Q => n53354, QN 
                           => n_1825);
   clk_r_REG15703_S1 : DFF_X1 port map( D => n2622, CK => CLK, Q => n53353, QN 
                           => n_1826);
   clk_r_REG15705_S1 : DFF_X1 port map( D => n2621, CK => CLK, Q => n53352, QN 
                           => n_1827);
   clk_r_REG16342_S1 : DFF_X1 port map( D => n2590, CK => CLK, Q => n53351, QN 
                           => n_1828);
   clk_r_REG15541_S1 : DFF_X1 port map( D => n2960, CK => CLK, Q => n53350, QN 
                           => n_1829);
   clk_r_REG16122_S1 : DFF_X1 port map( D => n2797, CK => CLK, Q => n53349, QN 
                           => n_1830);
   clk_r_REG16344_S1 : DFF_X1 port map( D => n2589, CK => CLK, Q => n53348, QN 
                           => n_1831);
   clk_r_REG15707_S1 : DFF_X1 port map( D => n2620, CK => CLK, Q => n53347, QN 
                           => n_1832);
   clk_r_REG15709_S1 : DFF_X1 port map( D => n2619, CK => CLK, Q => n53346, QN 
                           => n_1833);
   clk_r_REG15831_S1 : DFF_X1 port map( D => n2686, CK => CLK, Q => n53345, QN 
                           => n_1834);
   clk_r_REG16246_S1 : DFF_X1 port map( D => n2863, CK => CLK, Q => n53344, QN 
                           => n_1835);
   clk_r_REG15669_S1 : DFF_X1 port map( D => n3024, CK => CLK, Q => n53343, QN 
                           => n_1836);
   clk_r_REG15833_S1 : DFF_X1 port map( D => n2685, CK => CLK, Q => n53342, QN 
                           => n_1837);
   clk_r_REG15835_S1 : DFF_X1 port map( D => n2684, CK => CLK, Q => n53341, QN 
                           => n_1838);
   clk_r_REG16023_S1 : DFF_X1 port map( D => n2782, CK => CLK, Q => n53340, QN 
                           => n_1839);
   clk_r_REG15915_S1 : DFF_X1 port map( D => n2718, CK => CLK, Q => n53339, QN 
                           => n_1840);
   clk_r_REG15089_S1 : DFF_X1 port map( D => n3056, CK => CLK, Q => n53338, QN 
                           => n_1841);
   clk_r_REG15288_S1 : DFF_X1 port map( D => n3248, CK => CLK, Q => n53337, QN 
                           => n_1842);
   clk_r_REG15711_S1 : DFF_X1 port map( D => n2618, CK => CLK, Q => n53336, QN 
                           => n_1843);
   clk_r_REG16346_S1 : DFF_X1 port map( D => n2588, CK => CLK, Q => n53335, QN 
                           => n_1844);
   clk_r_REG15837_S1 : DFF_X1 port map( D => n2683, CK => CLK, Q => n53334, QN 
                           => n_1845);
   clk_r_REG15455_S1 : DFF_X1 port map( D => n2922, CK => CLK, Q => n53333, QN 
                           => n_1846);
   clk_r_REG16348_S1 : DFF_X1 port map( D => n2587, CK => CLK, Q => n53332, QN 
                           => n_1847);
   clk_r_REG15290_S1 : DFF_X1 port map( D => n3247, CK => CLK, Q => n53331, QN 
                           => n_1848);
   clk_r_REG16350_S1 : DFF_X1 port map( D => n2586, CK => CLK, Q => n53330, QN 
                           => n_1849);
   clk_r_REG15091_S1 : DFF_X1 port map( D => n3055, CK => CLK, Q => n53329, QN 
                           => n_1850);
   clk_r_REG15917_S1 : DFF_X1 port map( D => n2717, CK => CLK, Q => n53328, QN 
                           => n_1851);
   clk_r_REG16025_S1 : DFF_X1 port map( D => n2781, CK => CLK, Q => n53327, QN 
                           => n_1852);
   clk_r_REG15543_S1 : DFF_X1 port map( D => n2959, CK => CLK, Q => n53326, QN 
                           => n_1853);
   clk_r_REG15292_S1 : DFF_X1 port map( D => n3246, CK => CLK, Q => n53325, QN 
                           => n_1854);
   clk_r_REG15919_S1 : DFF_X1 port map( D => n2716, CK => CLK, Q => n53324, QN 
                           => n_1855);
   clk_r_REG15921_S1 : DFF_X1 port map( D => n2715, CK => CLK, Q => n53323, QN 
                           => n_1856);
   clk_r_REG16278_S1 : DFF_X1 port map( D => n2558, CK => CLK, Q => n53322, QN 
                           => n_1857);
   clk_r_REG15767_S1 : DFF_X1 port map( D => n2654, CK => CLK, Q => n53321, QN 
                           => n_1858);
   clk_r_REG15769_S1 : DFF_X1 port map( D => n2653, CK => CLK, Q => n53320, QN 
                           => n_1859);
   clk_r_REG15923_S1 : DFF_X1 port map( D => n2714, CK => CLK, Q => n53319, QN 
                           => n_1860);
   clk_r_REG15294_S1 : DFF_X1 port map( D => n3245, CK => CLK, Q => n53318, QN 
                           => n_1861);
   clk_r_REG15457_S1 : DFF_X1 port map( D => n2923, CK => CLK, Q => n53317, QN 
                           => n_1862);
   clk_r_REG16027_S1 : DFF_X1 port map( D => n2780, CK => CLK, Q => n53316, QN 
                           => n_1863);
   clk_r_REG16280_S1 : DFF_X1 port map( D => n2557, CK => CLK, Q => n53315, QN 
                           => n_1864);
   clk_r_REG16282_S1 : DFF_X1 port map( D => n2556, CK => CLK, Q => n53314, QN 
                           => n_1865);
   clk_r_REG16284_S1 : DFF_X1 port map( D => n2555, CK => CLK, Q => n53313, QN 
                           => n_1866);
   clk_r_REG16029_S1 : DFF_X1 port map( D => n2779, CK => CLK, Q => n53312, QN 
                           => n_1867);
   clk_r_REG15839_S1 : DFF_X1 port map( D => n2682, CK => CLK, Q => n53311, QN 
                           => n_1868);
   clk_r_REG15459_S1 : DFF_X1 port map( D => n2924, CK => CLK, Q => n53310, QN 
                           => n_1869);
   clk_r_REG15771_S1 : DFF_X1 port map( D => n2652, CK => CLK, Q => n53309, QN 
                           => n_1870);
   clk_r_REG16563_S1 : DFF_X1 port map( D => n3216, CK => CLK, Q => n53308, QN 
                           => n_1871);
   clk_r_REG15713_S1 : DFF_X1 port map( D => n2617, CK => CLK, Q => n53307, QN 
                           => n_1872);
   clk_r_REG16352_S1 : DFF_X1 port map( D => n2585, CK => CLK, Q => n53306, QN 
                           => n_1873);
   clk_r_REG16286_S1 : DFF_X1 port map( D => n2554, CK => CLK, Q => n53305, QN 
                           => n_1874);
   clk_r_REG16288_S1 : DFF_X1 port map( D => n2553, CK => CLK, Q => n53304, QN 
                           => n_1875);
   clk_r_REG15925_S1 : DFF_X1 port map( D => n2713, CK => CLK, Q => n53303, QN 
                           => n_1876);
   clk_r_REG15715_S1 : DFF_X1 port map( D => n2616, CK => CLK, Q => n53302, QN 
                           => n_1877);
   clk_r_REG15959_S1 : DFF_X1 port map( D => n2750, CK => CLK, Q => n53301, QN 
                           => n_1878);
   clk_r_REG16290_S1 : DFF_X1 port map( D => n2552, CK => CLK, Q => n53300, QN 
                           => n_1879);
   clk_r_REG15773_S1 : DFF_X1 port map( D => n2651, CK => CLK, Q => n53299, QN 
                           => n_1880);
   clk_r_REG15927_S1 : DFF_X1 port map( D => n2712, CK => CLK, Q => n53298, QN 
                           => n_1881);
   clk_r_REG15961_S1 : DFF_X1 port map( D => n2749, CK => CLK, Q => n53297, QN 
                           => n_1882);
   clk_r_REG15963_S1 : DFF_X1 port map( D => n2748, CK => CLK, Q => n53296, QN 
                           => n_1883);
   clk_r_REG16248_S1 : DFF_X1 port map( D => n2862, CK => CLK, Q => n53295, QN 
                           => n_1884);
   clk_r_REG15965_S1 : DFF_X1 port map( D => n2747, CK => CLK, Q => n53294, QN 
                           => n_1885);
   clk_r_REG15717_S1 : DFF_X1 port map( D => n2615, CK => CLK, Q => n53293, QN 
                           => n_1886);
   clk_r_REG16565_S1 : DFF_X1 port map( D => n3215, CK => CLK, Q => n53292, QN 
                           => n_1887);
   clk_r_REG16567_S1 : DFF_X1 port map( D => n3214, CK => CLK, Q => n53291, QN 
                           => n_1888);
   clk_r_REG16292_S1 : DFF_X1 port map( D => n2551, CK => CLK, Q => n53290, QN 
                           => n_1889);
   clk_r_REG16569_S1 : DFF_X1 port map( D => n3213, CK => CLK, Q => n53289, QN 
                           => n_1890);
   clk_r_REG16571_S1 : DFF_X1 port map( D => n3212, CK => CLK, Q => n53288, QN 
                           => n_1891);
   clk_r_REG16294_S1 : DFF_X1 port map( D => n2550, CK => CLK, Q => n53287, QN 
                           => n_1892);
   clk_r_REG16031_S1 : DFF_X1 port map( D => n2778, CK => CLK, Q => n53286, QN 
                           => n_1893);
   clk_r_REG15605_S1 : DFF_X1 port map( D => n2992, CK => CLK, Q => n53285, QN 
                           => n_1894);
   clk_r_REG15545_S1 : DFF_X1 port map( D => n2958, CK => CLK, Q => n53284, QN 
                           => n_1895);
   clk_r_REG15719_S1 : DFF_X1 port map( D => n2614, CK => CLK, Q => n53283, QN 
                           => n_1896);
   clk_r_REG15721_S1 : DFF_X1 port map( D => n2613, CK => CLK, Q => n53282, QN 
                           => n_1897);
   clk_r_REG15929_S1 : DFF_X1 port map( D => n2711, CK => CLK, Q => n53281, QN 
                           => n_1898);
   clk_r_REG15607_S1 : DFF_X1 port map( D => n2991, CK => CLK, Q => n53280, QN 
                           => n_1899);
   clk_r_REG15931_S1 : DFF_X1 port map( D => n2710, CK => CLK, Q => n53279, QN 
                           => n_1900);
   clk_r_REG15296_S1 : DFF_X1 port map( D => n3244, CK => CLK, Q => n53278, QN 
                           => n_1901);
   clk_r_REG16033_S1 : DFF_X1 port map( D => n2777, CK => CLK, Q => n53277, QN 
                           => n_1902);
   clk_r_REG15723_S1 : DFF_X1 port map( D => n2612, CK => CLK, Q => n53276, QN 
                           => n_1903);
   clk_r_REG16035_S1 : DFF_X1 port map( D => n2776, CK => CLK, Q => n53275, QN 
                           => n_1904);
   clk_r_REG16296_S1 : DFF_X1 port map( D => n2549, CK => CLK, Q => n53274, QN 
                           => n_1905);
   clk_r_REG15775_S1 : DFF_X1 port map( D => n2650, CK => CLK, Q => n53273, QN 
                           => n_1906);
   clk_r_REG15933_S1 : DFF_X1 port map( D => n2709, CK => CLK, Q => n53272, QN 
                           => n_1907);
   clk_r_REG15671_S1 : DFF_X1 port map( D => n3023, CK => CLK, Q => n53271, QN 
                           => n_1908);
   clk_r_REG16037_S1 : DFF_X1 port map( D => n2775, CK => CLK, Q => n53270, QN 
                           => n_1909);
   clk_r_REG16573_S1 : DFF_X1 port map( D => n3211, CK => CLK, Q => n53269, QN 
                           => n_1910);
   clk_r_REG16250_S1 : DFF_X1 port map( D => n2861, CK => CLK, Q => n53268, QN 
                           => n_1911);
   clk_r_REG16039_S1 : DFF_X1 port map( D => n2774, CK => CLK, Q => n53267, QN 
                           => n_1912);
   clk_r_REG16298_S1 : DFF_X1 port map( D => n2548, CK => CLK, Q => n53266, QN 
                           => n_1913);
   clk_r_REG15967_S1 : DFF_X1 port map( D => n2746, CK => CLK, Q => n53265, QN 
                           => n_1914);
   clk_r_REG15725_S1 : DFF_X1 port map( D => n2611, CK => CLK, Q => n53264, QN 
                           => n_1915);
   clk_r_REG16252_S1 : DFF_X1 port map( D => n2860, CK => CLK, Q => n53263, QN 
                           => n_1916);
   clk_r_REG16575_S1 : DFF_X1 port map( D => n3210, CK => CLK, Q => n53262, QN 
                           => n_1917);
   clk_r_REG16041_S1 : DFF_X1 port map( D => n2773, CK => CLK, Q => n53261, QN 
                           => n_1918);
   clk_r_REG15935_S1 : DFF_X1 port map( D => n2708, CK => CLK, Q => n53260, QN 
                           => n_1919);
   clk_r_REG15461_S1 : DFF_X1 port map( D => n2925, CK => CLK, Q => n53259, QN 
                           => n_1920);
   clk_r_REG15937_S1 : DFF_X1 port map( D => n2707, CK => CLK, Q => n53258, QN 
                           => n_1921);
   clk_r_REG15841_S1 : DFF_X1 port map( D => n2681, CK => CLK, Q => n53257, QN 
                           => n_1922);
   clk_r_REG16354_S1 : DFF_X1 port map( D => n2584, CK => CLK, Q => n53256, QN 
                           => n_1923);
   clk_r_REG15413_S1 : DFF_X1 port map( D => n2896, CK => CLK, Q => n53255, QN 
                           => n_1924);
   clk_r_REG16577_S1 : DFF_X1 port map( D => n3209, CK => CLK, Q => n53254, QN 
                           => n_1925);
   clk_r_REG16300_S1 : DFF_X1 port map( D => n2547, CK => CLK, Q => n53253, QN 
                           => n_1926);
   clk_r_REG15969_S1 : DFF_X1 port map( D => n2745, CK => CLK, Q => n53252, QN 
                           => n_1927);
   clk_r_REG15673_S1 : DFF_X1 port map( D => n3022, CK => CLK, Q => n53251, QN 
                           => n_1928);
   clk_r_REG16043_S1 : DFF_X1 port map( D => n2772, CK => CLK, Q => n53250, QN 
                           => n_1929);
   clk_r_REG16254_S1 : DFF_X1 port map( D => n2859, CK => CLK, Q => n53249, QN 
                           => n_1930);
   clk_r_REG16045_S1 : DFF_X1 port map( D => n2771, CK => CLK, Q => n53248, QN 
                           => n_1931);
   clk_r_REG16124_S1 : DFF_X1 port map( D => n2796, CK => CLK, Q => n53247, QN 
                           => n_1932);
   clk_r_REG16356_S1 : DFF_X1 port map( D => n2583, CK => CLK, Q => n53246, QN 
                           => n_1933);
   clk_r_REG16047_S1 : DFF_X1 port map( D => n2770, CK => CLK, Q => n53245, QN 
                           => n_1934);
   clk_r_REG13660_S1 : DFF_X1 port map( D => n3237, CK => CLK, Q => n53244, QN 
                           => n_1935);
   clk_r_REG16302_S1 : DFF_X1 port map( D => n2546, CK => CLK, Q => n53243, QN 
                           => n_1936);
   clk_r_REG15777_S1 : DFF_X1 port map( D => n2649, CK => CLK, Q => n53242, QN 
                           => n_1937);
   clk_r_REG16358_S1 : DFF_X1 port map( D => n2582, CK => CLK, Q => n53241, QN 
                           => n_1938);
   clk_r_REG15843_S1 : DFF_X1 port map( D => n2680, CK => CLK, Q => n53240, QN 
                           => n_1939);
   clk_r_REG15971_S1 : DFF_X1 port map( D => n2744, CK => CLK, Q => n53239, QN 
                           => n_1940);
   clk_r_REG15163_S1 : DFF_X1 port map( D => n3149, CK => CLK, Q => n53238, QN 
                           => n_1941);
   clk_r_REG16360_S1 : DFF_X1 port map( D => n2581, CK => CLK, Q => n53237, QN 
                           => n_1942);
   clk_r_REG15779_S1 : DFF_X1 port map( D => n2648, CK => CLK, Q => n53236, QN 
                           => n_1943);
   clk_r_REG15845_S1 : DFF_X1 port map( D => n2679, CK => CLK, Q => n53235, QN 
                           => n_1944);
   clk_r_REG15973_S1 : DFF_X1 port map( D => n2743, CK => CLK, Q => n53234, QN 
                           => n_1945);
   clk_r_REG15975_S1 : DFF_X1 port map( D => n2742, CK => CLK, Q => n53233, QN 
                           => n_1946);
   clk_r_REG16126_S1 : DFF_X1 port map( D => n2795, CK => CLK, Q => n53232, QN 
                           => n_1947);
   clk_r_REG16362_S1 : DFF_X1 port map( D => n2580, CK => CLK, Q => n53231, QN 
                           => n_1948);
   clk_r_REG15781_S1 : DFF_X1 port map( D => n2647, CK => CLK, Q => n53230, QN 
                           => n_1949);
   clk_r_REG15847_S1 : DFF_X1 port map( D => n2678, CK => CLK, Q => n53229, QN 
                           => n_1950);
   clk_r_REG15849_S1 : DFF_X1 port map( D => n2677, CK => CLK, Q => n53228, QN 
                           => n_1951);
   clk_r_REG15783_S1 : DFF_X1 port map( D => n2646, CK => CLK, Q => n53227, QN 
                           => n_1952);
   clk_r_REG16364_S1 : DFF_X1 port map( D => n2579, CK => CLK, Q => n53226, QN 
                           => n_1953);
   clk_r_REG16304_S1 : DFF_X1 port map( D => n2545, CK => CLK, Q => n53225, QN 
                           => n_1954);
   clk_r_REG15977_S1 : DFF_X1 port map( D => n2741, CK => CLK, Q => n53224, QN 
                           => n_1955);
   clk_r_REG15785_S1 : DFF_X1 port map( D => n2645, CK => CLK, Q => n53223, QN 
                           => n_1956);
   clk_r_REG15727_S1 : DFF_X1 port map( D => n2610, CK => CLK, Q => n53222, QN 
                           => n_1957);
   clk_r_REG15939_S1 : DFF_X1 port map( D => n2706, CK => CLK, Q => n53221, QN 
                           => n_1958);
   clk_r_REG16366_S1 : DFF_X1 port map( D => n2578, CK => CLK, Q => n53220, QN 
                           => n_1959);
   clk_r_REG15787_S1 : DFF_X1 port map( D => n2644, CK => CLK, Q => n53219, QN 
                           => n_1960);
   clk_r_REG15979_S1 : DFF_X1 port map( D => n2740, CK => CLK, Q => n53218, QN 
                           => n_1961);
   clk_r_REG15851_S1 : DFF_X1 port map( D => n2676, CK => CLK, Q => n53217, QN 
                           => n_1962);
   clk_r_REG16049_S1 : DFF_X1 port map( D => n2769, CK => CLK, Q => n53216, QN 
                           => n_1963);
   clk_r_REG15941_S1 : DFF_X1 port map( D => n2705, CK => CLK, Q => n53215, QN 
                           => n_1964);
   clk_r_REG15415_S1 : DFF_X1 port map( D => n2895, CK => CLK, Q => n53214, QN 
                           => n_1965);
   clk_r_REG15729_S1 : DFF_X1 port map( D => n2609, CK => CLK, Q => n53213, QN 
                           => n_1966);
   clk_r_REG15731_S1 : DFF_X1 port map( D => n2608, CK => CLK, Q => n53212, QN 
                           => n_1967);
   clk_r_REG13818_S1 : DFF_X1 port map( D => n2949, CK => CLK, Q => n53211, QN 
                           => n_1968);
   clk_r_REG15943_S1 : DFF_X1 port map( D => n2704, CK => CLK, Q => n53210, QN 
                           => n_1969);
   clk_r_REG15853_S1 : DFF_X1 port map( D => n2675, CK => CLK, Q => n53209, QN 
                           => n_1970);
   clk_r_REG16051_S1 : DFF_X1 port map( D => n2768, CK => CLK, Q => n53208, QN 
                           => n_1971);
   clk_r_REG15855_S1 : DFF_X1 port map( D => n2674, CK => CLK, Q => n53207, QN 
                           => n_1972);
   clk_r_REG15981_S1 : DFF_X1 port map( D => n2739, CK => CLK, Q => n53206, QN 
                           => n_1973);
   clk_r_REG15983_S1 : DFF_X1 port map( D => n2738, CK => CLK, Q => n53205, QN 
                           => n_1974);
   clk_r_REG15985_S1 : DFF_X1 port map( D => n2737, CK => CLK, Q => n53204, QN 
                           => n_1975);
   clk_r_REG15417_S1 : DFF_X1 port map( D => n2894, CK => CLK, Q => n53203, QN 
                           => n_1976);
   clk_r_REG16306_S1 : DFF_X1 port map( D => n2544, CK => CLK, Q => n53202, QN 
                           => n_1977);
   clk_r_REG15165_S1 : DFF_X1 port map( D => n3148, CK => CLK, Q => n53201, QN 
                           => n_1978);
   clk_r_REG16256_S1 : DFF_X1 port map( D => n2858, CK => CLK, Q => n53200, QN 
                           => n_1979);
   clk_r_REG15789_S1 : DFF_X1 port map( D => n2643, CK => CLK, Q => n53199, QN 
                           => n_1980);
   clk_r_REG15791_S1 : DFF_X1 port map( D => n2642, CK => CLK, Q => n53198, QN 
                           => n_1981);
   clk_r_REG15793_S1 : DFF_X1 port map( D => n2641, CK => CLK, Q => n53197, QN 
                           => n_1982);
   clk_r_REG14808_S1 : DFF_X1 port map( D => n3312, CK => CLK, Q => n53196, QN 
                           => n_1983);
   clk_r_REG15795_S1 : DFF_X1 port map( D => n2640, CK => CLK, Q => n53195, QN 
                           => n_1984);
   clk_r_REG15857_S1 : DFF_X1 port map( D => n2673, CK => CLK, Q => n53194, QN 
                           => n_1985);
   clk_r_REG16368_S1 : DFF_X1 port map( D => n2577, CK => CLK, Q => n53193, QN 
                           => n_1986);
   clk_r_REG15987_S1 : DFF_X1 port map( D => n2736, CK => CLK, Q => n53192, QN 
                           => n_1987);
   clk_r_REG15859_S1 : DFF_X1 port map( D => n2672, CK => CLK, Q => n53191, QN 
                           => n_1988);
   clk_r_REG16370_S1 : DFF_X1 port map( D => n2576, CK => CLK, Q => n53190, QN 
                           => n_1989);
   clk_r_REG16659_S1 : DFF_X1 port map( D => n3536, CK => CLK, Q => n53189, QN 
                           => n_1990);
   clk_r_REG16661_S1 : DFF_X1 port map( D => n3535, CK => CLK, Q => n53188, QN 
                           => n_1991);
   clk_r_REG16663_S1 : DFF_X1 port map( D => n3534, CK => CLK, Q => n53187, QN 
                           => n_1992);
   clk_r_REG16665_S1 : DFF_X1 port map( D => n3533, CK => CLK, Q => n53186, QN 
                           => n_1993);
   clk_r_REG16667_S1 : DFF_X1 port map( D => n3532, CK => CLK, Q => n53185, QN 
                           => n_1994);
   clk_r_REG16669_S1 : DFF_X1 port map( D => n3531, CK => CLK, Q => n53184, QN 
                           => n_1995);
   clk_r_REG16671_S1 : DFF_X1 port map( D => n3530, CK => CLK, Q => n53183, QN 
                           => n_1996);
   clk_r_REG16673_S1 : DFF_X1 port map( D => n3529, CK => CLK, Q => n53182, QN 
                           => n_1997);
   clk_r_REG13649_S1 : DFF_X1 port map( D => n3557, CK => CLK, Q => n53181, QN 
                           => n_1998);
   clk_r_REG16619_S1 : DFF_X1 port map( D => n3556, CK => CLK, Q => n53180, QN 
                           => n_1999);
   clk_r_REG15437_S1 : DFF_X1 port map( D => n2948, CK => CLK, Q => n53179, QN 
                           => n_2000);
   clk_r_REG16128_S1 : DFF_X1 port map( D => n2794, CK => CLK, Q => n53178, QN 
                           => n_2001);
   clk_r_REG14740_S1 : DFF_X1 port map( D => n3440, CK => CLK, Q => n53177, QN 
                           => n_2002);
   clk_r_REG16186_S1 : DFF_X1 port map( D => n2829, CK => CLK, Q => n53176, QN 
                           => n_2003);
   clk_r_REG15224_S1 : DFF_X1 port map( D => n3184, CK => CLK, Q => n53175, QN 
                           => n_2004);
   clk_r_REG15675_S1 : DFF_X1 port map( D => n3021, CK => CLK, Q => n53174, QN 
                           => n_2005);
   clk_r_REG15547_S1 : DFF_X1 port map( D => n2957, CK => CLK, Q => n53173, QN 
                           => n_2006);
   clk_r_REG15549_S1 : DFF_X1 port map( D => n2956, CK => CLK, Q => n53172, QN 
                           => n_2007);
   clk_r_REG16130_S1 : DFF_X1 port map( D => n2793, CK => CLK, Q => n53171, QN 
                           => n_2008);
   clk_r_REG15439_S1 : DFF_X1 port map( D => n2947, CK => CLK, Q => n53170, QN 
                           => n_2009);
   clk_r_REG15551_S1 : DFF_X1 port map( D => n2955, CK => CLK, Q => n53169, QN 
                           => n_2010);
   clk_r_REG16258_S1 : DFF_X1 port map( D => n2857, CK => CLK, Q => n53168, QN 
                           => n_2011);
   clk_r_REG16438_S1 : DFF_X1 port map( D => n3086, CK => CLK, Q => n53167, QN 
                           => n_2012);
   clk_r_REG16188_S1 : DFF_X1 port map( D => n2828, CK => CLK, Q => n53166, QN 
                           => n_2013);
   clk_r_REG15167_S1 : DFF_X1 port map( D => n3147, CK => CLK, Q => n53165, QN 
                           => n_2014);
   clk_r_REG15419_S1 : DFF_X1 port map( D => n2893, CK => CLK, Q => n53164, QN 
                           => n_2015);
   clk_r_REG16190_S1 : DFF_X1 port map( D => n2827, CK => CLK, Q => n53163, QN 
                           => n_2016);
   clk_r_REG14664_S1 : DFF_X1 port map( D => n3376, CK => CLK, Q => n53162, QN 
                           => n_2017);
   clk_r_REG13735_S1 : DFF_X1 port map( D => n2821, CK => CLK, Q => n53161, QN 
                           => n_2018);
   clk_r_REG16440_S1 : DFF_X1 port map( D => n3085, CK => CLK, Q => n53160, QN 
                           => n_2019);
   clk_r_REG15441_S1 : DFF_X1 port map( D => n2946, CK => CLK, Q => n53159, QN 
                           => n_2020);
   clk_r_REG16501_S1 : DFF_X1 port map( D => n3119, CK => CLK, Q => n53158, QN 
                           => n_2021);
   clk_r_REG15443_S1 : DFF_X1 port map( D => n2945, CK => CLK, Q => n53157, QN 
                           => n_2022);
   clk_r_REG15421_S1 : DFF_X1 port map( D => n2892, CK => CLK, Q => n53156, QN 
                           => n_2023);
   clk_r_REG15423_S1 : DFF_X1 port map( D => n2891, CK => CLK, Q => n53155, QN 
                           => n_2024);
   clk_r_REG15425_S1 : DFF_X1 port map( D => n2890, CK => CLK, Q => n53154, QN 
                           => n_2025);
   clk_r_REG15553_S1 : DFF_X1 port map( D => n2954, CK => CLK, Q => n53153, QN 
                           => n_2026);
   clk_r_REG15463_S1 : DFF_X1 port map( D => n2926, CK => CLK, Q => n53152, QN 
                           => n_2027);
   clk_r_REG14948_S1 : DFF_X1 port map( D => n3280, CK => CLK, Q => n53151, QN 
                           => n_2028);
   clk_r_REG16442_S1 : DFF_X1 port map( D => n3084, CK => CLK, Q => n53150, QN 
                           => n_2029);
   clk_r_REG15351_S1 : DFF_X1 port map( D => n3344, CK => CLK, Q => n53149, QN 
                           => n_2030);
   clk_r_REG16192_S1 : DFF_X1 port map( D => n2826, CK => CLK, Q => n53148, QN 
                           => n_2031);
   clk_r_REG16076_S1 : DFF_X1 port map( D => n2820, CK => CLK, Q => n53147, QN 
                           => n_2032);
   clk_r_REG14950_S1 : DFF_X1 port map( D => n3279, CK => CLK, Q => n53146, QN 
                           => n_2033);
   clk_r_REG15093_S1 : DFF_X1 port map( D => n3054, CK => CLK, Q => n53145, QN 
                           => n_2034);
   clk_r_REG16523_S1 : DFF_X1 port map( D => n3236, CK => CLK, Q => n53144, QN 
                           => n_2035);
   clk_r_REG14952_S1 : DFF_X1 port map( D => n3278, CK => CLK, Q => n53143, QN 
                           => n_2036);
   clk_r_REG14954_S1 : DFF_X1 port map( D => n3277, CK => CLK, Q => n53142, QN 
                           => n_2037);
   clk_r_REG15298_S1 : DFF_X1 port map( D => n3243, CK => CLK, Q => n53141, QN 
                           => n_2038);
   clk_r_REG15300_S1 : DFF_X1 port map( D => n3242, CK => CLK, Q => n53140, QN 
                           => n_2039);
   clk_r_REG15302_S1 : DFF_X1 port map( D => n3241, CK => CLK, Q => n53139, QN 
                           => n_2040);
   clk_r_REG14410_S1 : DFF_X1 port map( D => n3408, CK => CLK, Q => n53138, QN 
                           => n_2041);
   clk_r_REG16525_S1 : DFF_X1 port map( D => n3235, CK => CLK, Q => n53137, QN 
                           => n_2042);
   clk_r_REG15095_S1 : DFF_X1 port map( D => n3053, CK => CLK, Q => n53136, QN 
                           => n_2043);
   clk_r_REG15555_S1 : DFF_X1 port map( D => n2953, CK => CLK, Q => n53135, QN 
                           => n_2044);
   clk_r_REG15097_S1 : DFF_X1 port map( D => n3052, CK => CLK, Q => n53134, QN 
                           => n_2045);
   clk_r_REG15099_S1 : DFF_X1 port map( D => n3051, CK => CLK, Q => n53133, QN 
                           => n_2046);
   clk_r_REG15101_S1 : DFF_X1 port map( D => n3050, CK => CLK, Q => n53132, QN 
                           => n_2047);
   clk_r_REG16444_S1 : DFF_X1 port map( D => n3083, CK => CLK, Q => n53131, QN 
                           => n_2048);
   clk_r_REG16503_S1 : DFF_X1 port map( D => n3118, CK => CLK, Q => n53130, QN 
                           => n_2049);
   clk_r_REG15169_S1 : DFF_X1 port map( D => n3146, CK => CLK, Q => n53129, QN 
                           => n_2050);
   clk_r_REG15226_S1 : DFF_X1 port map( D => n3183, CK => CLK, Q => n53128, QN 
                           => n_2051);
   clk_r_REG15022_S1 : DFF_X1 port map( D => n3504, CK => CLK, Q => n53127, QN 
                           => n_2052);
   clk_r_REG16527_S1 : DFF_X1 port map( D => n3234, CK => CLK, Q => n53126, QN 
                           => n_2053);
   clk_r_REG13850_S1 : DFF_X1 port map( D => n3269, CK => CLK, Q => n53125, QN 
                           => n_2054);
   clk_r_REG14956_S1 : DFF_X1 port map( D => n3276, CK => CLK, Q => n53124, QN 
                           => n_2055);
   clk_r_REG16446_S1 : DFF_X1 port map( D => n3082, CK => CLK, Q => n53123, QN 
                           => n_2056);
   clk_r_REG15248_S1 : DFF_X1 port map( D => n3268, CK => CLK, Q => n53122, QN 
                           => n_2057);
   clk_r_REG14958_S1 : DFF_X1 port map( D => n3275, CK => CLK, Q => n53121, QN 
                           => n_2058);
   clk_r_REG16505_S1 : DFF_X1 port map( D => n3117, CK => CLK, Q => n53120, QN 
                           => n_2059);
   clk_r_REG15250_S1 : DFF_X1 port map( D => n3267, CK => CLK, Q => n53119, QN 
                           => n_2060);
   clk_r_REG16529_S1 : DFF_X1 port map( D => n3233, CK => CLK, Q => n53118, QN 
                           => n_2061);
   clk_r_REG16507_S1 : DFF_X1 port map( D => n3116, CK => CLK, Q => n53117, QN 
                           => n_2062);
   clk_r_REG16579_S1 : DFF_X1 port map( D => n3208, CK => CLK, Q => n53116, QN 
                           => n_2063);
   clk_r_REG16509_S1 : DFF_X1 port map( D => n3115, CK => CLK, Q => n53115, QN 
                           => n_2064);
   clk_r_REG16078_S1 : DFF_X1 port map( D => n2819, CK => CLK, Q => n53114, QN 
                           => n_2065);
   clk_r_REG15171_S1 : DFF_X1 port map( D => n3145, CK => CLK, Q => n53113, QN 
                           => n_2066);
   clk_r_REG13905_S1 : DFF_X1 port map( D => n3173, CK => CLK, Q => n53112, QN 
                           => n_2067);
   clk_r_REG15117_S1 : DFF_X1 port map( D => n3172, CK => CLK, Q => n53111, QN 
                           => n_2068);
   clk_r_REG16194_S1 : DFF_X1 port map( D => n2825, CK => CLK, Q => n53110, QN 
                           => n_2069);
   clk_r_REG16531_S1 : DFF_X1 port map( D => n3232, CK => CLK, Q => n53109, QN 
                           => n_2070);
   clk_r_REG14880_S1 : DFF_X1 port map( D => n3472, CK => CLK, Q => n53108, QN 
                           => n_2071);
   clk_r_REG15427_S1 : DFF_X1 port map( D => n2889, CK => CLK, Q => n53107, QN 
                           => n_2072);
   clk_r_REG15445_S1 : DFF_X1 port map( D => n2944, CK => CLK, Q => n53106, QN 
                           => n_2073);
   clk_r_REG13811_S1 : DFF_X1 port map( D => n2981, CK => CLK, Q => n53105, QN 
                           => n_2074);
   clk_r_REG15609_S1 : DFF_X1 port map( D => n2990, CK => CLK, Q => n53104, QN 
                           => n_2075);
   clk_r_REG15103_S1 : DFF_X1 port map( D => n3049, CK => CLK, Q => n53103, QN 
                           => n_2076);
   clk_r_REG16448_S1 : DFF_X1 port map( D => n3081, CK => CLK, Q => n53102, QN 
                           => n_2077);
   clk_r_REG16511_S1 : DFF_X1 port map( D => n3114, CK => CLK, Q => n53101, QN 
                           => n_2078);
   clk_r_REG15119_S1 : DFF_X1 port map( D => n3171, CK => CLK, Q => n53100, QN 
                           => n_2079);
   clk_r_REG15228_S1 : DFF_X1 port map( D => n3182, CK => CLK, Q => n53099, QN 
                           => n_2080);
   clk_r_REG15230_S1 : DFF_X1 port map( D => n3181, CK => CLK, Q => n53098, QN 
                           => n_2081);
   clk_r_REG15232_S1 : DFF_X1 port map( D => n3180, CK => CLK, Q => n53097, QN 
                           => n_2082);
   clk_r_REG15234_S1 : DFF_X1 port map( D => n3179, CK => CLK, Q => n53096, QN 
                           => n_2083);
   clk_r_REG15252_S1 : DFF_X1 port map( D => n3266, CK => CLK, Q => n53095, QN 
                           => n_2084);
   clk_r_REG14960_S1 : DFF_X1 port map( D => n3274, CK => CLK, Q => n53094, QN 
                           => n_2085);
   clk_r_REG16080_S1 : DFF_X1 port map( D => n2818, CK => CLK, Q => n53093, QN 
                           => n_2086);
   clk_r_REG15121_S1 : DFF_X1 port map( D => n3170, CK => CLK, Q => n53092, QN 
                           => n_2087);
   clk_r_REG15236_S1 : DFF_X1 port map( D => n3178, CK => CLK, Q => n53091, QN 
                           => n_2088);
   clk_r_REG16581_S1 : DFF_X1 port map( D => n3207, CK => CLK, Q => n53090, QN 
                           => n_2089);
   clk_r_REG15254_S1 : DFF_X1 port map( D => n3265, CK => CLK, Q => n53089, QN 
                           => n_2090);
   clk_r_REG14962_S1 : DFF_X1 port map( D => n3273, CK => CLK, Q => n53088, QN 
                           => n_2091);
   clk_r_REG15465_S1 : DFF_X1 port map( D => n2927, CK => CLK, Q => n53087, QN 
                           => n_2092);
   clk_r_REG15501_S1 : DFF_X1 port map( D => n2980, CK => CLK, Q => n53086, QN 
                           => n_2093);
   clk_r_REG13918_S1 : DFF_X1 port map( D => n3077, CK => CLK, Q => n53085, QN 
                           => n_2094);
   clk_r_REG13688_S1 : DFF_X1 port map( D => n3109, CK => CLK, Q => n53084, QN 
                           => n_2095);
   clk_r_REG16513_S1 : DFF_X1 port map( D => n3113, CK => CLK, Q => n53083, QN 
                           => n_2096);
   clk_r_REG15123_S1 : DFF_X1 port map( D => n3169, CK => CLK, Q => n53082, QN 
                           => n_2097);
   clk_r_REG15238_S1 : DFF_X1 port map( D => n3177, CK => CLK, Q => n53081, QN 
                           => n_2098);
   clk_r_REG14032_S1 : DFF_X1 port map( D => n3301, CK => CLK, Q => n53080, QN 
                           => n_2099);
   clk_r_REG15304_S1 : DFF_X1 port map( D => n3240, CK => CLK, Q => n53079, QN 
                           => n_2100);
   clk_r_REG16583_S1 : DFF_X1 port map( D => n3206, CK => CLK, Q => n53078, QN 
                           => n_2101);
   clk_r_REG13721_S1 : DFF_X1 port map( D => n2885, CK => CLK, Q => n53077, QN 
                           => n_2102);
   clk_r_REG16204_S1 : DFF_X1 port map( D => n2884, CK => CLK, Q => n53076, QN 
                           => n_2103);
   clk_r_REG16206_S1 : DFF_X1 port map( D => n2883, CK => CLK, Q => n53075, QN 
                           => n_2104);
   clk_r_REG16208_S1 : DFF_X1 port map( D => n2882, CK => CLK, Q => n53074, QN 
                           => n_2105);
   clk_r_REG16210_S1 : DFF_X1 port map( D => n2881, CK => CLK, Q => n53073, QN 
                           => n_2106);
   clk_r_REG16260_S1 : DFF_X1 port map( D => n2856, CK => CLK, Q => n53072, QN 
                           => n_2107);
   clk_r_REG16212_S1 : DFF_X1 port map( D => n2880, CK => CLK, Q => n53071, QN 
                           => n_2108);
   clk_r_REG13825_S1 : DFF_X1 port map( D => n2917, CK => CLK, Q => n53070, QN 
                           => n_2109);
   clk_r_REG13869_S1 : DFF_X1 port map( D => n3205, CK => CLK, Q => n53069, QN 
                           => n_2110);
   clk_r_REG15611_S1 : DFF_X1 port map( D => n2989, CK => CLK, Q => n53068, QN 
                           => n_2111);
   clk_r_REG15613_S1 : DFF_X1 port map( D => n2988, CK => CLK, Q => n53067, QN 
                           => n_2112);
   clk_r_REG15615_S1 : DFF_X1 port map( D => n2987, CK => CLK, Q => n53066, QN 
                           => n_2113);
   clk_r_REG15617_S1 : DFF_X1 port map( D => n2986, CK => CLK, Q => n53065, QN 
                           => n_2114);
   clk_r_REG15619_S1 : DFF_X1 port map( D => n2985, CK => CLK, Q => n53064, QN 
                           => n_2115);
   clk_r_REG13804_S1 : DFF_X1 port map( D => n3013, CK => CLK, Q => n53063, QN 
                           => n_2116);
   clk_r_REG15565_S1 : DFF_X1 port map( D => n3012, CK => CLK, Q => n53062, QN 
                           => n_2117);
   clk_r_REG15677_S1 : DFF_X1 port map( D => n3020, CK => CLK, Q => n53061, QN 
                           => n_2118);
   clk_r_REG15679_S1 : DFF_X1 port map( D => n3019, CK => CLK, Q => n53060, QN 
                           => n_2119);
   clk_r_REG15681_S1 : DFF_X1 port map( D => n3018, CK => CLK, Q => n53059, QN 
                           => n_2120);
   clk_r_REG15683_S1 : DFF_X1 port map( D => n3017, CK => CLK, Q => n53058, QN 
                           => n_2121);
   clk_r_REG13795_S1 : DFF_X1 port map( D => n3045, CK => CLK, Q => n53057, QN 
                           => n_2122);
   clk_r_REG15567_S1 : DFF_X1 port map( D => n3011, CK => CLK, Q => n53056, QN 
                           => n_2123);
   clk_r_REG15629_S1 : DFF_X1 port map( D => n3044, CK => CLK, Q => n53055, QN 
                           => n_2124);
   clk_r_REG15631_S1 : DFF_X1 port map( D => n3043, CK => CLK, Q => n53054, QN 
                           => n_2125);
   clk_r_REG16132_S1 : DFF_X1 port map( D => n2792, CK => CLK, Q => n53053, QN 
                           => n_2126);
   clk_r_REG13728_S1 : DFF_X1 port map( D => n2853, CK => CLK, Q => n53052, QN 
                           => n_2127);
   clk_r_REG16262_S1 : DFF_X1 port map( D => n2855, CK => CLK, Q => n53051, QN 
                           => n_2128);
   clk_r_REG15373_S1 : DFF_X1 port map( D => n2916, CK => CLK, Q => n53050, QN 
                           => n_2129);
   clk_r_REG15467_S1 : DFF_X1 port map( D => n2928, CK => CLK, Q => n53049, QN 
                           => n_2130);
   clk_r_REG15503_S1 : DFF_X1 port map( D => n2979, CK => CLK, Q => n53048, QN 
                           => n_2131);
   clk_r_REG15049_S1 : DFF_X1 port map( D => n3076, CK => CLK, Q => n53047, QN 
                           => n_2132);
   clk_r_REG15633_S1 : DFF_X1 port map( D => n3042, CK => CLK, Q => n53046, QN 
                           => n_2133);
   clk_r_REG13674_S1 : DFF_X1 port map( D => n3141, CK => CLK, Q => n53045, QN 
                           => n_2134);
   clk_r_REG16394_S1 : DFF_X1 port map( D => n3108, CK => CLK, Q => n53044, QN 
                           => n_2135);
   clk_r_REG16621_S1 : DFF_X1 port map( D => n3555, CK => CLK, Q => n53043, QN 
                           => n_2136);
   clk_r_REG15353_S1 : DFF_X1 port map( D => n3343, CK => CLK, Q => n53042, QN 
                           => n_2137);
   clk_r_REG15173_S1 : DFF_X1 port map( D => n3144, CK => CLK, Q => n53041, QN 
                           => n_2138);
   clk_r_REG14810_S1 : DFF_X1 port map( D => n3311, CK => CLK, Q => n53040, QN 
                           => n_2139);
   clk_r_REG14412_S1 : DFF_X1 port map( D => n3407, CK => CLK, Q => n53039, QN 
                           => n_2140);
   clk_r_REG14666_S1 : DFF_X1 port map( D => n3375, CK => CLK, Q => n53038, QN 
                           => n_2141);
   clk_r_REG16533_S1 : DFF_X1 port map( D => n3231, CK => CLK, Q => n53037, QN 
                           => n_2142);
   clk_r_REG15024_S1 : DFF_X1 port map( D => n3503, CK => CLK, Q => n53036, QN 
                           => n_2143);
   clk_r_REG14882_S1 : DFF_X1 port map( D => n3471, CK => CLK, Q => n53035, QN 
                           => n_2144);
   clk_r_REG14742_S1 : DFF_X1 port map( D => n3439, CK => CLK, Q => n53034, QN 
                           => n_2145);
   clk_r_REG15026_S1 : DFF_X1 port map( D => n3502, CK => CLK, Q => n53033, QN 
                           => n_2146);
   clk_r_REG14884_S1 : DFF_X1 port map( D => n3470, CK => CLK, Q => n53032, QN 
                           => n_2147);
   clk_r_REG14744_S1 : DFF_X1 port map( D => n3438, CK => CLK, Q => n53031, QN 
                           => n_2148);
   clk_r_REG14746_S1 : DFF_X1 port map( D => n3437, CK => CLK, Q => n53030, QN 
                           => n_2149);
   clk_r_REG15028_S1 : DFF_X1 port map( D => n3501, CK => CLK, Q => n53029, QN 
                           => n_2150);
   clk_r_REG15030_S1 : DFF_X1 port map( D => n3500, CK => CLK, Q => n53028, QN 
                           => n_2151);
   clk_r_REG15032_S1 : DFF_X1 port map( D => n3499, CK => CLK, Q => n53027, QN 
                           => n_2152);
   clk_r_REG14748_S1 : DFF_X1 port map( D => n3436, CK => CLK, Q => n53026, QN 
                           => n_2153);
   clk_r_REG14750_S1 : DFF_X1 port map( D => n3435, CK => CLK, Q => n53025, QN 
                           => n_2154);
   clk_r_REG14414_S1 : DFF_X1 port map( D => n3406, CK => CLK, Q => n53024, QN 
                           => n_2155);
   clk_r_REG14416_S1 : DFF_X1 port map( D => n3405, CK => CLK, Q => n53023, QN 
                           => n_2156);
   clk_r_REG14418_S1 : DFF_X1 port map( D => n3404, CK => CLK, Q => n53022, QN 
                           => n_2157);
   clk_r_REG14420_S1 : DFF_X1 port map( D => n3403, CK => CLK, Q => n53021, QN 
                           => n_2158);
   clk_r_REG14668_S1 : DFF_X1 port map( D => n3374, CK => CLK, Q => n53020, QN 
                           => n_2159);
   clk_r_REG14812_S1 : DFF_X1 port map( D => n3310, CK => CLK, Q => n53019, QN 
                           => n_2160);
   clk_r_REG15375_S1 : DFF_X1 port map( D => n2915, CK => CLK, Q => n53018, QN 
                           => n_2161);
   clk_r_REG15034_S1 : DFF_X1 port map( D => n3498, CK => CLK, Q => n53017, QN 
                           => n_2162);
   clk_r_REG14886_S1 : DFF_X1 port map( D => n3469, CK => CLK, Q => n53016, QN 
                           => n_2163);
   clk_r_REG14752_S1 : DFF_X1 port map( D => n3434, CK => CLK, Q => n53015, QN 
                           => n_2164);
   clk_r_REG14422_S1 : DFF_X1 port map( D => n3402, CK => CLK, Q => n53014, QN 
                           => n_2165);
   clk_r_REG14670_S1 : DFF_X1 port map( D => n3373, CK => CLK, Q => n53013, QN 
                           => n_2166);
   clk_r_REG15036_S1 : DFF_X1 port map( D => n3497, CK => CLK, Q => n53012, QN 
                           => n_2167);
   clk_r_REG14011_S1 : DFF_X1 port map( D => n3525, CK => CLK, Q => n53011, QN 
                           => n_2168);
   clk_r_REG14672_S1 : DFF_X1 port map( D => n3372, CK => CLK, Q => n53010, QN 
                           => n_2169);
   clk_r_REG14674_S1 : DFF_X1 port map( D => n3371, CK => CLK, Q => n53009, QN 
                           => n_2170);
   clk_r_REG14754_S1 : DFF_X1 port map( D => n3433, CK => CLK, Q => n53008, QN 
                           => n_2171);
   clk_r_REG14814_S1 : DFF_X1 port map( D => n3309, CK => CLK, Q => n53007, QN 
                           => n_2172);
   clk_r_REG16082_S1 : DFF_X1 port map( D => n2817, CK => CLK, Q => n53006, QN 
                           => n_2173);
   clk_r_REG14676_S1 : DFF_X1 port map( D => n3370, CK => CLK, Q => n53005, QN 
                           => n_2174);
   clk_r_REG16140_S1 : DFF_X1 port map( D => n2852, CK => CLK, Q => n53004, QN 
                           => n_2175);
   clk_r_REG16084_S1 : DFF_X1 port map( D => n2816, CK => CLK, Q => n53003, QN 
                           => n_2176);
   clk_r_REG15355_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n53002, QN 
                           => n_2177);
   clk_r_REG14424_S1 : DFF_X1 port map( D => n3401, CK => CLK, Q => n53001, QN 
                           => n_2178);
   clk_r_REG14678_S1 : DFF_X1 port map( D => n3369, CK => CLK, Q => n53000, QN 
                           => n_2179);
   clk_r_REG16142_S1 : DFF_X1 port map( D => n2851, CK => CLK, Q => n52999, QN 
                           => n_2180);
   clk_r_REG15357_S1 : DFF_X1 port map( D => n3341, CK => CLK, Q => n52998, QN 
                           => n_2181);
   clk_r_REG15359_S1 : DFF_X1 port map( D => n3340, CK => CLK, Q => n52997, QN 
                           => n_2182);
   clk_r_REG14816_S1 : DFF_X1 port map( D => n3308, CK => CLK, Q => n52996, QN 
                           => n_2183);
   clk_r_REG14141_S1 : DFF_X1 port map( D => n3397, CK => CLK, Q => n52995, QN 
                           => n_2184);
   clk_r_REG14888_S1 : DFF_X1 port map( D => n3468, CK => CLK, Q => n52994, QN 
                           => n_2185);
   clk_r_REG15361_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n52993, QN 
                           => n_2186);
   clk_r_REG15363_S1 : DFF_X1 port map( D => n3338, CK => CLK, Q => n52992, QN 
                           => n_2187);
   clk_r_REG14890_S1 : DFF_X1 port map( D => n3467, CK => CLK, Q => n52991, QN 
                           => n_2188);
   clk_r_REG14892_S1 : DFF_X1 port map( D => n3466, CK => CLK, Q => n52990, QN 
                           => n_2189);
   clk_r_REG14818_S1 : DFF_X1 port map( D => n3307, CK => CLK, Q => n52989, QN 
                           => n_2190);
   clk_r_REG14894_S1 : DFF_X1 port map( D => n3465, CK => CLK, Q => n52988, QN 
                           => n_2191);
   clk_r_REG14066_S1 : DFF_X1 port map( D => n3493, CK => CLK, Q => n52987, QN 
                           => n_2192);
   clk_r_REG15365_S1 : DFF_X1 port map( D => n3337, CK => CLK, Q => n52986, QN 
                           => n_2193);
   clk_r_REG14120_S1 : DFF_X1 port map( D => n3461, CK => CLK, Q => n52985, QN 
                           => n_2194);
   clk_r_REG14160_S1 : DFF_X1 port map( D => n3429, CK => CLK, Q => n52984, QN 
                           => n_2195);
   clk_r_REG14820_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n52983, QN 
                           => n_2196);
   clk_r_REG14822_S1 : DFF_X1 port map( D => n3305, CK => CLK, Q => n52982, QN 
                           => n_2197);
   clk_r_REG13837_S1 : DFF_X1 port map( D => n3365, CK => CLK, Q => n52981, QN 
                           => n_2198);
   clk_r_REG14079_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n52980, QN 
                           => n_2199);
   clk_r_REG14768_S1 : DFF_X1 port map( D => n3332, CK => CLK, Q => n52979, QN 
                           => n_2200);
   clk_r_REG16144_S1 : DFF_X1 port map( D => n2850, CK => CLK, Q => n52978, QN 
                           => n_2201);
   clk_r_REG15377_S1 : DFF_X1 port map( D => n2914, CK => CLK, Q => n52977, QN 
                           => n_2202);
   clk_r_REG15469_S1 : DFF_X1 port map( D => n2943, CK => CLK, Q => n52976, QN 
                           => n_2203);
   clk_r_REG15505_S1 : DFF_X1 port map( D => n2978, CK => CLK, Q => n52975, QN 
                           => n_2204);
   clk_r_REG15051_S1 : DFF_X1 port map( D => n3075, CK => CLK, Q => n52974, QN 
                           => n_2205);
   clk_r_REG16396_S1 : DFF_X1 port map( D => n3107, CK => CLK, Q => n52973, QN 
                           => n_2206);
   clk_r_REG16459_S1 : DFF_X1 port map( D => n3140, CK => CLK, Q => n52972, QN 
                           => n_2207);
   clk_r_REG15053_S1 : DFF_X1 port map( D => n3074, CK => CLK, Q => n52971, QN 
                           => n_2208);
   clk_r_REG16134_S1 : DFF_X1 port map( D => n2791, CK => CLK, Q => n52970, QN 
                           => n_2209);
   clk_r_REG15311_S1 : DFF_X1 port map( D => n3364, CK => CLK, Q => n52969, QN 
                           => n_2210);
   clk_r_REG14624_S1 : DFF_X1 port map( D => n3396, CK => CLK, Q => n52968, QN 
                           => n_2211);
   clk_r_REG16146_S1 : DFF_X1 port map( D => n2849, CK => CLK, Q => n52967, QN 
                           => n_2212);
   clk_r_REG15507_S1 : DFF_X1 port map( D => n2977, CK => CLK, Q => n52966, QN 
                           => n_2213);
   clk_r_REG15557_S1 : DFF_X1 port map( D => n2952, CK => CLK, Q => n52965, QN 
                           => n_2214);
   clk_r_REG16136_S1 : DFF_X1 port map( D => n2790, CK => CLK, Q => n52964, QN 
                           => n_2215);
   clk_r_REG14626_S1 : DFF_X1 port map( D => n3395, CK => CLK, Q => n52963, QN 
                           => n_2216);
   clk_r_REG14628_S1 : DFF_X1 port map( D => n3394, CK => CLK, Q => n52962, QN 
                           => n_2217);
   clk_r_REG16264_S1 : DFF_X1 port map( D => n2854, CK => CLK, Q => n52961, QN 
                           => n_2218);
   clk_r_REG15313_S1 : DFF_X1 port map( D => n3363, CK => CLK, Q => n52960, QN 
                           => n_2219);
   clk_r_REG15315_S1 : DFF_X1 port map( D => n3362, CK => CLK, Q => n52959, QN 
                           => n_2220);
   clk_r_REG15317_S1 : DFF_X1 port map( D => n3361, CK => CLK, Q => n52958, QN 
                           => n_2221);
   clk_r_REG16214_S1 : DFF_X1 port map( D => n2879, CK => CLK, Q => n52957, QN 
                           => n_2222);
   clk_r_REG15055_S1 : DFF_X1 port map( D => n3073, CK => CLK, Q => n52956, QN 
                           => n_2223);
   clk_r_REG15105_S1 : DFF_X1 port map( D => n3048, CK => CLK, Q => n52955, QN 
                           => n_2224);
   clk_r_REG15471_S1 : DFF_X1 port map( D => n2942, CK => CLK, Q => n52954, QN 
                           => n_2225);
   clk_r_REG14630_S1 : DFF_X1 port map( D => n3393, CK => CLK, Q => n52953, QN 
                           => n_2226);
   clk_r_REG16216_S1 : DFF_X1 port map( D => n2878, CK => CLK, Q => n52952, QN 
                           => n_2227);
   clk_r_REG16218_S1 : DFF_X1 port map( D => n2877, CK => CLK, Q => n52951, QN 
                           => n_2228);
   clk_r_REG15379_S1 : DFF_X1 port map( D => n2913, CK => CLK, Q => n52950, QN 
                           => n_2229);
   clk_r_REG15429_S1 : DFF_X1 port map( D => n2888, CK => CLK, Q => n52949, QN 
                           => n_2230);
   clk_r_REG15509_S1 : DFF_X1 port map( D => n2976, CK => CLK, Q => n52948, QN 
                           => n_2231);
   clk_r_REG16086_S1 : DFF_X1 port map( D => n2815, CK => CLK, Q => n52947, QN 
                           => n_2232);
   clk_r_REG15559_S1 : DFF_X1 port map( D => n2951, CK => CLK, Q => n52946, QN 
                           => n_2233);
   clk_r_REG15561_S1 : DFF_X1 port map( D => n2950, CK => CLK, Q => n52945, QN 
                           => n_2234);
   clk_r_REG15473_S1 : DFF_X1 port map( D => n2941, CK => CLK, Q => n52944, QN 
                           => n_2235);
   clk_r_REG16220_S1 : DFF_X1 port map( D => n2876, CK => CLK, Q => n52943, QN 
                           => n_2236);
   clk_r_REG15057_S1 : DFF_X1 port map( D => n3072, CK => CLK, Q => n52942, QN 
                           => n_2237);
   clk_r_REG14680_S1 : DFF_X1 port map( D => n3368, CK => CLK, Q => n52941, QN 
                           => n_2238);
   clk_r_REG14700_S1 : DFF_X1 port map( D => n3460, CK => CLK, Q => n52940, QN 
                           => n_2239);
   clk_r_REG16623_S1 : DFF_X1 port map( D => n3554, CK => CLK, Q => n52939, QN 
                           => n_2240);
   clk_r_REG16625_S1 : DFF_X1 port map( D => n3553, CK => CLK, Q => n52938, QN 
                           => n_2241);
   clk_r_REG14702_S1 : DFF_X1 port map( D => n3459, CK => CLK, Q => n52937, QN 
                           => n_2242);
   clk_r_REG14632_S1 : DFF_X1 port map( D => n3392, CK => CLK, Q => n52936, QN 
                           => n_2243);
   clk_r_REG15367_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n52935, QN 
                           => n_2244);
   clk_r_REG14704_S1 : DFF_X1 port map( D => n3458, CK => CLK, Q => n52934, QN 
                           => n_2245);
   clk_r_REG14840_S1 : DFF_X1 port map( D => n3492, CK => CLK, Q => n52933, QN 
                           => n_2246);
   clk_r_REG15107_S1 : DFF_X1 port map( D => n3047, CK => CLK, Q => n52932, QN 
                           => n_2247);
   clk_r_REG14370_S1 : DFF_X1 port map( D => n3428, CK => CLK, Q => n52931, QN 
                           => n_2248);
   clk_r_REG16088_S1 : DFF_X1 port map( D => n2814, CK => CLK, Q => n52930, QN 
                           => n_2249);
   clk_r_REG14842_S1 : DFF_X1 port map( D => n3491, CK => CLK, Q => n52929, QN 
                           => n_2250);
   clk_r_REG14706_S1 : DFF_X1 port map( D => n3457, CK => CLK, Q => n52928, QN 
                           => n_2251);
   clk_r_REG14756_S1 : DFF_X1 port map( D => n3432, CK => CLK, Q => n52927, QN 
                           => n_2252);
   clk_r_REG14372_S1 : DFF_X1 port map( D => n3427, CK => CLK, Q => n52926, QN 
                           => n_2253);
   clk_r_REG14374_S1 : DFF_X1 port map( D => n3426, CK => CLK, Q => n52925, QN 
                           => n_2254);
   clk_r_REG14844_S1 : DFF_X1 port map( D => n3490, CK => CLK, Q => n52924, QN 
                           => n_2255);
   clk_r_REG14846_S1 : DFF_X1 port map( D => n3489, CK => CLK, Q => n52923, QN 
                           => n_2256);
   clk_r_REG14708_S1 : DFF_X1 port map( D => n3456, CK => CLK, Q => n52922, QN 
                           => n_2257);
   clk_r_REG14376_S1 : DFF_X1 port map( D => n3425, CK => CLK, Q => n52921, QN 
                           => n_2258);
   clk_r_REG15319_S1 : DFF_X1 port map( D => n3360, CK => CLK, Q => n52920, QN 
                           => n_2259);
   clk_r_REG14982_S1 : DFF_X1 port map( D => n3524, CK => CLK, Q => n52919, QN 
                           => n_2260);
   clk_r_REG14984_S1 : DFF_X1 port map( D => n3523, CK => CLK, Q => n52918, QN 
                           => n_2261);
   clk_r_REG14986_S1 : DFF_X1 port map( D => n3522, CK => CLK, Q => n52917, QN 
                           => n_2262);
   clk_r_REG14988_S1 : DFF_X1 port map( D => n3521, CK => CLK, Q => n52916, QN 
                           => n_2263);
   clk_r_REG14896_S1 : DFF_X1 port map( D => n3464, CK => CLK, Q => n52915, QN 
                           => n_2264);
   clk_r_REG16398_S1 : DFF_X1 port map( D => n3106, CK => CLK, Q => n52914, QN 
                           => n_2265);
   clk_r_REG14848_S1 : DFF_X1 port map( D => n3488, CK => CLK, Q => n52913, QN 
                           => n_2266);
   clk_r_REG16196_S1 : DFF_X1 port map( D => n2824, CK => CLK, Q => n52912, QN 
                           => n_2267);
   clk_r_REG14426_S1 : DFF_X1 port map( D => n3400, CK => CLK, Q => n52911, QN 
                           => n_2268);
   clk_r_REG15569_S1 : DFF_X1 port map( D => n3010, CK => CLK, Q => n52910, QN 
                           => n_2269);
   clk_r_REG15038_S1 : DFF_X1 port map( D => n3496, CK => CLK, Q => n52909, QN 
                           => n_2270);
   clk_r_REG15571_S1 : DFF_X1 port map( D => n3009, CK => CLK, Q => n52908, QN 
                           => n_2271);
   clk_r_REG14378_S1 : DFF_X1 port map( D => n3424, CK => CLK, Q => n52907, QN 
                           => n_2272);
   clk_r_REG15635_S1 : DFF_X1 port map( D => n3041, CK => CLK, Q => n52906, QN 
                           => n_2273);
   clk_r_REG15621_S1 : DFF_X1 port map( D => n2984, CK => CLK, Q => n52905, QN 
                           => n_2274);
   clk_r_REG14990_S1 : DFF_X1 port map( D => n3520, CK => CLK, Q => n52904, QN 
                           => n_2275);
   clk_r_REG14770_S1 : DFF_X1 port map( D => n3331, CK => CLK, Q => n52903, QN 
                           => n_2276);
   clk_r_REG14772_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n52902, QN 
                           => n_2277);
   clk_r_REG16535_S1 : DFF_X1 port map( D => n3230, CK => CLK, Q => n52901, QN 
                           => n_2278);
   clk_r_REG15573_S1 : DFF_X1 port map( D => n3008, CK => CLK, Q => n52900, QN 
                           => n_2279);
   clk_r_REG15623_S1 : DFF_X1 port map( D => n2983, CK => CLK, Q => n52899, QN 
                           => n_2280);
   clk_r_REG16537_S1 : DFF_X1 port map( D => n3229, CK => CLK, Q => n52898, QN 
                           => n_2281);
   clk_r_REG16675_S1 : DFF_X1 port map( D => n3528, CK => CLK, Q => n52897, QN 
                           => n_2282);
   clk_r_REG16539_S1 : DFF_X1 port map( D => n3228, CK => CLK, Q => n52896, QN 
                           => n_2283);
   clk_r_REG16627_S1 : DFF_X1 port map( D => n3552, CK => CLK, Q => n52895, QN 
                           => n_2284);
   clk_r_REG16541_S1 : DFF_X1 port map( D => n3227, CK => CLK, Q => n52894, QN 
                           => n_2285);
   clk_r_REG16677_S1 : DFF_X1 port map( D => n3527, CK => CLK, Q => n52893, QN 
                           => n_2286);
   clk_r_REG16543_S1 : DFF_X1 port map( D => n3226, CK => CLK, Q => n52892, QN 
                           => n_2287);
   clk_r_REG16679_S1 : DFF_X1 port map( D => n3526, CK => CLK, Q => n52891, QN 
                           => n_2288);
   clk_r_REG16629_S1 : DFF_X1 port map( D => n3551, CK => CLK, Q => n52890, QN 
                           => n_2289);
   clk_r_REG16545_S1 : DFF_X1 port map( D => n3225, CK => CLK, Q => n52889, QN 
                           => n_2290);
   clk_r_REG15369_S1 : DFF_X1 port map( D => n3335, CK => CLK, Q => n52888, QN 
                           => n_2291);
   clk_r_REG14774_S1 : DFF_X1 port map( D => n3329, CK => CLK, Q => n52887, QN 
                           => n_2292);
   clk_r_REG15040_S1 : DFF_X1 port map( D => n3495, CK => CLK, Q => n52886, QN 
                           => n_2293);
   clk_r_REG14682_S1 : DFF_X1 port map( D => n3367, CK => CLK, Q => n52885, QN 
                           => n_2294);
   clk_r_REG14428_S1 : DFF_X1 port map( D => n3399, CK => CLK, Q => n52884, QN 
                           => n_2295);
   clk_r_REG14758_S1 : DFF_X1 port map( D => n3431, CK => CLK, Q => n52883, QN 
                           => n_2296);
   clk_r_REG14898_S1 : DFF_X1 port map( D => n3463, CK => CLK, Q => n52882, QN 
                           => n_2297);
   clk_r_REG15042_S1 : DFF_X1 port map( D => n3494, CK => CLK, Q => n52881, QN 
                           => n_2298);
   clk_r_REG14900_S1 : DFF_X1 port map( D => n3462, CK => CLK, Q => n52880, QN 
                           => n_2299);
   clk_r_REG14760_S1 : DFF_X1 port map( D => n3430, CK => CLK, Q => n52879, QN 
                           => n_2300);
   clk_r_REG14430_S1 : DFF_X1 port map( D => n3398, CK => CLK, Q => n52878, QN 
                           => n_2301);
   clk_r_REG14684_S1 : DFF_X1 port map( D => n3366, CK => CLK, Q => n52877, QN 
                           => n_2302);
   clk_r_REG14824_S1 : DFF_X1 port map( D => n3304, CK => CLK, Q => n52876, QN 
                           => n_2303);
   clk_r_REG15371_S1 : DFF_X1 port map( D => n3334, CK => CLK, Q => n52875, QN 
                           => n_2304);
   clk_r_REG14776_S1 : DFF_X1 port map( D => n3328, CK => CLK, Q => n52874, QN 
                           => n_2305);
   clk_r_REG16547_S1 : DFF_X1 port map( D => n3224, CK => CLK, Q => n52873, QN 
                           => n_2306);
   clk_r_REG16549_S1 : DFF_X1 port map( D => n3223, CK => CLK, Q => n52872, QN 
                           => n_2307);
   clk_r_REG15381_S1 : DFF_X1 port map( D => n2912, CK => CLK, Q => n52871, QN 
                           => n_2308);
   clk_r_REG15431_S1 : DFF_X1 port map( D => n2887, CK => CLK, Q => n52870, QN 
                           => n_2309);
   clk_r_REG15433_S1 : DFF_X1 port map( D => n2886, CK => CLK, Q => n52869, QN 
                           => n_2310);
   clk_r_REG16148_S1 : DFF_X1 port map( D => n2848, CK => CLK, Q => n52868, QN 
                           => n_2311);
   clk_r_REG14826_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n52867, QN 
                           => n_2312);
   clk_r_REG14828_S1 : DFF_X1 port map( D => n3302, CK => CLK, Q => n52866, QN 
                           => n_2313);
   clk_r_REG15383_S1 : DFF_X1 port map( D => n2911, CK => CLK, Q => n52865, QN 
                           => n_2314);
   clk_r_REG15385_S1 : DFF_X1 port map( D => n2910, CK => CLK, Q => n52864, QN 
                           => n_2315);
   clk_r_REG16198_S1 : DFF_X1 port map( D => n2823, CK => CLK, Q => n52863, QN 
                           => n_2316);
   clk_r_REG14778_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n52862, QN 
                           => n_2317);
   clk_r_REG15387_S1 : DFF_X1 port map( D => n2909, CK => CLK, Q => n52861, QN 
                           => n_2318);
   clk_r_REG16200_S1 : DFF_X1 port map( D => n2822, CK => CLK, Q => n52860, QN 
                           => n_2319);
   clk_r_REG16090_S1 : DFF_X1 port map( D => n2813, CK => CLK, Q => n52859, QN 
                           => n_2320);
   clk_r_REG15109_S1 : DFF_X1 port map( D => n3046, CK => CLK, Q => n52858, QN 
                           => n_2321);
   clk_r_REG15625_S1 : DFF_X1 port map( D => n2982, CK => CLK, Q => n52857, QN 
                           => n_2322);
   clk_r_REG15511_S1 : DFF_X1 port map( D => n2975, CK => CLK, Q => n52856, QN 
                           => n_2323);
   clk_r_REG15475_S1 : DFF_X1 port map( D => n2940, CK => CLK, Q => n52855, QN 
                           => n_2324);
   clk_r_REG16222_S1 : DFF_X1 port map( D => n2875, CK => CLK, Q => n52854, QN 
                           => n_2325);
   clk_r_REG14908_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n52853, QN 
                           => n_2326);
   clk_r_REG15256_S1 : DFF_X1 port map( D => n3264, CK => CLK, Q => n52852, QN 
                           => n_2327);
   clk_r_REG15184_S1 : DFF_X1 port map( D => n3204, CK => CLK, Q => n52851, QN 
                           => n_2328);
   clk_r_REG16461_S1 : DFF_X1 port map( D => n3139, CK => CLK, Q => n52850, QN 
                           => n_2329);
   clk_r_REG16400_S1 : DFF_X1 port map( D => n3105, CK => CLK, Q => n52849, QN 
                           => n_2330);
   clk_r_REG15059_S1 : DFF_X1 port map( D => n3071, CK => CLK, Q => n52848, QN 
                           => n_2331);
   clk_r_REG15685_S1 : DFF_X1 port map( D => n3016, CK => CLK, Q => n52847, QN 
                           => n_2332);
   clk_r_REG15575_S1 : DFF_X1 port map( D => n3007, CK => CLK, Q => n52846, QN 
                           => n_2333);
   clk_r_REG15637_S1 : DFF_X1 port map( D => n3040, CK => CLK, Q => n52845, QN 
                           => n_2334);
   clk_r_REG15513_S1 : DFF_X1 port map( D => n2974, CK => CLK, Q => n52844, QN 
                           => n_2335);
   clk_r_REG15477_S1 : DFF_X1 port map( D => n2939, CK => CLK, Q => n52843, QN 
                           => n_2336);
   clk_r_REG16224_S1 : DFF_X1 port map( D => n2874, CK => CLK, Q => n52842, QN 
                           => n_2337);
   clk_r_REG16463_S1 : DFF_X1 port map( D => n3138, CK => CLK, Q => n52841, QN 
                           => n_2338);
   clk_r_REG15186_S1 : DFF_X1 port map( D => n3203, CK => CLK, Q => n52840, QN 
                           => n_2339);
   clk_r_REG15306_S1 : DFF_X1 port map( D => n3239, CK => CLK, Q => n52839, QN 
                           => n_2340);
   clk_r_REG14910_S1 : DFF_X1 port map( D => n3299, CK => CLK, Q => n52838, QN 
                           => n_2341);
   clk_r_REG15308_S1 : DFF_X1 port map( D => n3238, CK => CLK, Q => n52837, QN 
                           => n_2342);
   clk_r_REG15258_S1 : DFF_X1 port map( D => n3263, CK => CLK, Q => n52836, QN 
                           => n_2343);
   clk_r_REG15260_S1 : DFF_X1 port map( D => n3262, CK => CLK, Q => n52835, QN 
                           => n_2344);
   clk_r_REG15262_S1 : DFF_X1 port map( D => n3261, CK => CLK, Q => n52834, QN 
                           => n_2345);
   clk_r_REG15264_S1 : DFF_X1 port map( D => n3260, CK => CLK, Q => n52833, QN 
                           => n_2346);
   clk_r_REG15266_S1 : DFF_X1 port map( D => n3259, CK => CLK, Q => n52832, QN 
                           => n_2347);
   clk_r_REG14912_S1 : DFF_X1 port map( D => n3298, CK => CLK, Q => n52831, QN 
                           => n_2348);
   clk_r_REG14914_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n52830, QN 
                           => n_2349);
   clk_r_REG14964_S1 : DFF_X1 port map( D => n3272, CK => CLK, Q => n52829, QN 
                           => n_2350);
   clk_r_REG14916_S1 : DFF_X1 port map( D => n3296, CK => CLK, Q => n52828, QN 
                           => n_2351);
   clk_r_REG14966_S1 : DFF_X1 port map( D => n3271, CK => CLK, Q => n52827, QN 
                           => n_2352);
   clk_r_REG14968_S1 : DFF_X1 port map( D => n3270, CK => CLK, Q => n52826, QN 
                           => n_2353);
   clk_r_REG16450_S1 : DFF_X1 port map( D => n3080, CK => CLK, Q => n52825, QN 
                           => n_2354);
   clk_r_REG16402_S1 : DFF_X1 port map( D => n3104, CK => CLK, Q => n52824, QN 
                           => n_2355);
   clk_r_REG15061_S1 : DFF_X1 port map( D => n3070, CK => CLK, Q => n52823, QN 
                           => n_2356);
   clk_r_REG16452_S1 : DFF_X1 port map( D => n3079, CK => CLK, Q => n52822, QN 
                           => n_2357);
   clk_r_REG16454_S1 : DFF_X1 port map( D => n3078, CK => CLK, Q => n52821, QN 
                           => n_2358);
   clk_r_REG16465_S1 : DFF_X1 port map( D => n3137, CK => CLK, Q => n52820, QN 
                           => n_2359);
   clk_r_REG16515_S1 : DFF_X1 port map( D => n3112, CK => CLK, Q => n52819, QN 
                           => n_2360);
   clk_r_REG16467_S1 : DFF_X1 port map( D => n3136, CK => CLK, Q => n52818, QN 
                           => n_2361);
   clk_r_REG16517_S1 : DFF_X1 port map( D => n3111, CK => CLK, Q => n52817, QN 
                           => n_2362);
   clk_r_REG16519_S1 : DFF_X1 port map( D => n3110, CK => CLK, Q => n52816, QN 
                           => n_2363);
   clk_r_REG15125_S1 : DFF_X1 port map( D => n3168, CK => CLK, Q => n52815, QN 
                           => n_2364);
   clk_r_REG15515_S1 : DFF_X1 port map( D => n2973, CK => CLK, Q => n52814, QN 
                           => n_2365);
   clk_r_REG15175_S1 : DFF_X1 port map( D => n3143, CK => CLK, Q => n52813, QN 
                           => n_2366);
   clk_r_REG15177_S1 : DFF_X1 port map( D => n3142, CK => CLK, Q => n52812, QN 
                           => n_2367);
   clk_r_REG15127_S1 : DFF_X1 port map( D => n3167, CK => CLK, Q => n52811, QN 
                           => n_2368);
   clk_r_REG15129_S1 : DFF_X1 port map( D => n3166, CK => CLK, Q => n52810, QN 
                           => n_2369);
   clk_r_REG15577_S1 : DFF_X1 port map( D => n3006, CK => CLK, Q => n52809, QN 
                           => n_2370);
   clk_r_REG15188_S1 : DFF_X1 port map( D => n3202, CK => CLK, Q => n52808, QN 
                           => n_2371);
   clk_r_REG15190_S1 : DFF_X1 port map( D => n3201, CK => CLK, Q => n52807, QN 
                           => n_2372);
   clk_r_REG15240_S1 : DFF_X1 port map( D => n3176, CK => CLK, Q => n52806, QN 
                           => n_2373);
   clk_r_REG15192_S1 : DFF_X1 port map( D => n3200, CK => CLK, Q => n52805, QN 
                           => n_2374);
   clk_r_REG15242_S1 : DFF_X1 port map( D => n3175, CK => CLK, Q => n52804, QN 
                           => n_2375);
   clk_r_REG15479_S1 : DFF_X1 port map( D => n2938, CK => CLK, Q => n52803, QN 
                           => n_2376);
   clk_r_REG15244_S1 : DFF_X1 port map( D => n3174, CK => CLK, Q => n52802, QN 
                           => n_2377);
   clk_r_REG15687_S1 : DFF_X1 port map( D => n3015, CK => CLK, Q => n52801, QN 
                           => n_2378);
   clk_r_REG15689_S1 : DFF_X1 port map( D => n3014, CK => CLK, Q => n52800, QN 
                           => n_2379);
   clk_r_REG15639_S1 : DFF_X1 port map( D => n3039, CK => CLK, Q => n52799, QN 
                           => n_2380);
   clk_r_REG15641_S1 : DFF_X1 port map( D => n3038, CK => CLK, Q => n52798, QN 
                           => n_2381);
   clk_r_REG15643_S1 : DFF_X1 port map( D => n3037, CK => CLK, Q => n52797, QN 
                           => n_2382);
   clk_r_REG15321_S1 : DFF_X1 port map( D => n3359, CK => CLK, Q => n52796, QN 
                           => n_2383);
   clk_r_REG14850_S1 : DFF_X1 port map( D => n3487, CK => CLK, Q => n52795, QN 
                           => n_2384);
   clk_r_REG16469_S1 : DFF_X1 port map( D => n3135, CK => CLK, Q => n52794, QN 
                           => n_2385);
   clk_r_REG14380_S1 : DFF_X1 port map( D => n3423, CK => CLK, Q => n52793, QN 
                           => n_2386);
   clk_r_REG15323_S1 : DFF_X1 port map( D => n3358, CK => CLK, Q => n52792, QN 
                           => n_2387);
   clk_r_REG14710_S1 : DFF_X1 port map( D => n3455, CK => CLK, Q => n52791, QN 
                           => n_2388);
   clk_r_REG16471_S1 : DFF_X1 port map( D => n3134, CK => CLK, Q => n52790, QN 
                           => n_2389);
   clk_r_REG14382_S1 : DFF_X1 port map( D => n3422, CK => CLK, Q => n52789, QN 
                           => n_2390);
   clk_r_REG14852_S1 : DFF_X1 port map( D => n3486, CK => CLK, Q => n52788, QN 
                           => n_2391);
   clk_r_REG14780_S1 : DFF_X1 port map( D => n3326, CK => CLK, Q => n52787, QN 
                           => n_2392);
   clk_r_REG15325_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n52786, QN 
                           => n_2393);
   clk_r_REG15131_S1 : DFF_X1 port map( D => n3165, CK => CLK, Q => n52785, QN 
                           => n_2394);
   clk_r_REG14634_S1 : DFF_X1 port map( D => n3391, CK => CLK, Q => n52784, QN 
                           => n_2395);
   clk_r_REG15327_S1 : DFF_X1 port map( D => n3356, CK => CLK, Q => n52783, QN 
                           => n_2396);
   clk_r_REG16473_S1 : DFF_X1 port map( D => n3133, CK => CLK, Q => n52782, QN 
                           => n_2397);
   clk_r_REG14636_S1 : DFF_X1 port map( D => n3390, CK => CLK, Q => n52781, QN 
                           => n_2398);
   clk_r_REG15133_S1 : DFF_X1 port map( D => n3164, CK => CLK, Q => n52780, QN 
                           => n_2399);
   clk_r_REG14782_S1 : DFF_X1 port map( D => n3325, CK => CLK, Q => n52779, QN 
                           => n_2400);
   clk_r_REG15135_S1 : DFF_X1 port map( D => n3163, CK => CLK, Q => n52778, QN 
                           => n_2401);
   clk_r_REG14638_S1 : DFF_X1 port map( D => n3389, CK => CLK, Q => n52777, QN 
                           => n_2402);
   clk_r_REG14992_S1 : DFF_X1 port map( D => n3519, CK => CLK, Q => n52776, QN 
                           => n_2403);
   clk_r_REG15194_S1 : DFF_X1 port map( D => n3199, CK => CLK, Q => n52775, QN 
                           => n_2404);
   clk_r_REG14994_S1 : DFF_X1 port map( D => n3518, CK => CLK, Q => n52774, QN 
                           => n_2405);
   clk_r_REG16631_S1 : DFF_X1 port map( D => n3550, CK => CLK, Q => n52773, QN 
                           => n_2406);
   clk_r_REG15196_S1 : DFF_X1 port map( D => n3198, CK => CLK, Q => n52772, QN 
                           => n_2407);
   clk_r_REG14854_S1 : DFF_X1 port map( D => n3485, CK => CLK, Q => n52771, QN 
                           => n_2408);
   clk_r_REG14712_S1 : DFF_X1 port map( D => n3454, CK => CLK, Q => n52770, QN 
                           => n_2409);
   clk_r_REG16633_S1 : DFF_X1 port map( D => n3549, CK => CLK, Q => n52769, QN 
                           => n_2410);
   clk_r_REG14384_S1 : DFF_X1 port map( D => n3421, CK => CLK, Q => n52768, QN 
                           => n_2411);
   clk_r_REG14856_S1 : DFF_X1 port map( D => n3484, CK => CLK, Q => n52767, QN 
                           => n_2412);
   clk_r_REG15389_S1 : DFF_X1 port map( D => n2908, CK => CLK, Q => n52766, QN 
                           => n_2413);
   clk_r_REG14640_S1 : DFF_X1 port map( D => n3388, CK => CLK, Q => n52765, QN 
                           => n_2414);
   clk_r_REG14714_S1 : DFF_X1 port map( D => n3453, CK => CLK, Q => n52764, QN 
                           => n_2415);
   clk_r_REG14716_S1 : DFF_X1 port map( D => n3452, CK => CLK, Q => n52763, QN 
                           => n_2416);
   clk_r_REG14718_S1 : DFF_X1 port map( D => n3451, CK => CLK, Q => n52762, QN 
                           => n_2417);
   clk_r_REG15198_S1 : DFF_X1 port map( D => n3197, CK => CLK, Q => n52761, QN 
                           => n_2418);
   clk_r_REG14642_S1 : DFF_X1 port map( D => n3387, CK => CLK, Q => n52760, QN 
                           => n_2419);
   clk_r_REG15063_S1 : DFF_X1 port map( D => n3069, CK => CLK, Q => n52759, QN 
                           => n_2420);
   clk_r_REG16551_S1 : DFF_X1 port map( D => n3222, CK => CLK, Q => n52758, QN 
                           => n_2421);
   clk_r_REG14996_S1 : DFF_X1 port map( D => n3517, CK => CLK, Q => n52757, QN 
                           => n_2422);
   clk_r_REG14386_S1 : DFF_X1 port map( D => n3420, CK => CLK, Q => n52756, QN 
                           => n_2423);
   clk_r_REG14998_S1 : DFF_X1 port map( D => n3516, CK => CLK, Q => n52755, QN 
                           => n_2424);
   clk_r_REG14858_S1 : DFF_X1 port map( D => n3483, CK => CLK, Q => n52754, QN 
                           => n_2425);
   clk_r_REG14784_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n52753, QN 
                           => n_2426);
   clk_r_REG15000_S1 : DFF_X1 port map( D => n3515, CK => CLK, Q => n52752, QN 
                           => n_2427);
   clk_r_REG14388_S1 : DFF_X1 port map( D => n3419, CK => CLK, Q => n52751, QN 
                           => n_2428);
   clk_r_REG16635_S1 : DFF_X1 port map( D => n3548, CK => CLK, Q => n52750, QN 
                           => n_2429);
   clk_r_REG15065_S1 : DFF_X1 port map( D => n3068, CK => CLK, Q => n52749, QN 
                           => n_2430);
   clk_r_REG15329_S1 : DFF_X1 port map( D => n3355, CK => CLK, Q => n52748, QN 
                           => n_2431);
   clk_r_REG14786_S1 : DFF_X1 port map( D => n3323, CK => CLK, Q => n52747, QN 
                           => n_2432);
   clk_r_REG16150_S1 : DFF_X1 port map( D => n2847, CK => CLK, Q => n52746, QN 
                           => n_2433);
   clk_r_REG15067_S1 : DFF_X1 port map( D => n3067, CK => CLK, Q => n52745, QN 
                           => n_2434);
   clk_r_REG15268_S1 : DFF_X1 port map( D => n3258, CK => CLK, Q => n52744, QN 
                           => n_2435);
   clk_r_REG16152_S1 : DFF_X1 port map( D => n2846, CK => CLK, Q => n52743, QN 
                           => n_2436);
   clk_r_REG15391_S1 : DFF_X1 port map( D => n2907, CK => CLK, Q => n52742, QN 
                           => n_2437);
   clk_r_REG15517_S1 : DFF_X1 port map( D => n2972, CK => CLK, Q => n52741, QN 
                           => n_2438);
   clk_r_REG14918_S1 : DFF_X1 port map( D => n3295, CK => CLK, Q => n52740, QN 
                           => n_2439);
   clk_r_REG16404_S1 : DFF_X1 port map( D => n3103, CK => CLK, Q => n52739, QN 
                           => n_2440);
   clk_r_REG14920_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n52738, QN 
                           => n_2441);
   clk_r_REG15645_S1 : DFF_X1 port map( D => n3036, CK => CLK, Q => n52737, QN 
                           => n_2442);
   clk_r_REG14922_S1 : DFF_X1 port map( D => n3293, CK => CLK, Q => n52736, QN 
                           => n_2443);
   clk_r_REG15519_S1 : DFF_X1 port map( D => n2971, CK => CLK, Q => n52735, QN 
                           => n_2444);
   clk_r_REG16154_S1 : DFF_X1 port map( D => n2845, CK => CLK, Q => n52734, QN 
                           => n_2445);
   clk_r_REG16156_S1 : DFF_X1 port map( D => n2844, CK => CLK, Q => n52733, QN 
                           => n_2446);
   clk_r_REG16092_S1 : DFF_X1 port map( D => n2812, CK => CLK, Q => n52732, QN 
                           => n_2447);
   clk_r_REG16158_S1 : DFF_X1 port map( D => n2843, CK => CLK, Q => n52731, QN 
                           => n_2448);
   clk_r_REG16094_S1 : DFF_X1 port map( D => n2811, CK => CLK, Q => n52730, QN 
                           => n_2449);
   clk_r_REG16096_S1 : DFF_X1 port map( D => n2810, CK => CLK, Q => n52729, QN 
                           => n_2450);
   clk_r_REG16098_S1 : DFF_X1 port map( D => n2809, CK => CLK, Q => n52728, QN 
                           => n_2451);
   clk_r_REG15393_S1 : DFF_X1 port map( D => n2906, CK => CLK, Q => n52727, QN 
                           => n_2452);
   clk_r_REG16406_S1 : DFF_X1 port map( D => n3102, CK => CLK, Q => n52726, QN 
                           => n_2453);
   clk_r_REG15395_S1 : DFF_X1 port map( D => n2905, CK => CLK, Q => n52725, QN 
                           => n_2454);
   clk_r_REG16408_S1 : DFF_X1 port map( D => n3101, CK => CLK, Q => n52724, QN 
                           => n_2455);
   clk_r_REG16410_S1 : DFF_X1 port map( D => n3100, CK => CLK, Q => n52723, QN 
                           => n_2456);
   clk_r_REG15270_S1 : DFF_X1 port map( D => n3257, CK => CLK, Q => n52722, QN 
                           => n_2457);
   clk_r_REG16100_S1 : DFF_X1 port map( D => n2808, CK => CLK, Q => n52721, QN 
                           => n_2458);
   clk_r_REG14924_S1 : DFF_X1 port map( D => n3292, CK => CLK, Q => n52720, QN 
                           => n_2459);
   clk_r_REG15521_S1 : DFF_X1 port map( D => n2970, CK => CLK, Q => n52719, QN 
                           => n_2460);
   clk_r_REG15397_S1 : DFF_X1 port map( D => n2904, CK => CLK, Q => n52718, QN 
                           => n_2461);
   clk_r_REG16475_S1 : DFF_X1 port map( D => n3132, CK => CLK, Q => n52717, QN 
                           => n_2462);
   clk_r_REG15647_S1 : DFF_X1 port map( D => n3035, CK => CLK, Q => n52716, QN 
                           => n_2463);
   clk_r_REG16160_S1 : DFF_X1 port map( D => n2842, CK => CLK, Q => n52715, QN 
                           => n_2464);
   clk_r_REG14788_S1 : DFF_X1 port map( D => n3322, CK => CLK, Q => n52714, QN 
                           => n_2465);
   clk_r_REG15200_S1 : DFF_X1 port map( D => n3196, CK => CLK, Q => n52713, QN 
                           => n_2466);
   clk_r_REG16637_S1 : DFF_X1 port map( D => n3547, CK => CLK, Q => n52712, QN 
                           => n_2467);
   clk_r_REG15137_S1 : DFF_X1 port map( D => n3162, CK => CLK, Q => n52711, QN 
                           => n_2468);
   clk_r_REG16553_S1 : DFF_X1 port map( D => n3221, CK => CLK, Q => n52710, QN 
                           => n_2469);
   clk_r_REG16102_S1 : DFF_X1 port map( D => n2807, CK => CLK, Q => n52709, QN 
                           => n_2470);
   clk_r_REG16555_S1 : DFF_X1 port map( D => n3220, CK => CLK, Q => n52708, QN 
                           => n_2471);
   clk_r_REG16557_S1 : DFF_X1 port map( D => n3219, CK => CLK, Q => n52707, QN 
                           => n_2472);
   clk_r_REG15399_S1 : DFF_X1 port map( D => n2903, CK => CLK, Q => n52706, QN 
                           => n_2473);
   clk_r_REG16639_S1 : DFF_X1 port map( D => n3546, CK => CLK, Q => n52705, QN 
                           => n_2474);
   clk_r_REG16641_S1 : DFF_X1 port map( D => n3545, CK => CLK, Q => n52704, QN 
                           => n_2475);
   clk_r_REG16643_S1 : DFF_X1 port map( D => n3544, CK => CLK, Q => n52703, QN 
                           => n_2476);
   clk_r_REG15401_S1 : DFF_X1 port map( D => n2902, CK => CLK, Q => n52702, QN 
                           => n_2477);
   clk_r_REG15649_S1 : DFF_X1 port map( D => n3034, CK => CLK, Q => n52701, QN 
                           => n_2478);
   clk_r_REG15651_S1 : DFF_X1 port map( D => n3033, CK => CLK, Q => n52700, QN 
                           => n_2479);
   clk_r_REG16162_S1 : DFF_X1 port map( D => n2841, CK => CLK, Q => n52699, QN 
                           => n_2480);
   clk_r_REG16164_S1 : DFF_X1 port map( D => n2840, CK => CLK, Q => n52698, QN 
                           => n_2481);
   clk_r_REG15403_S1 : DFF_X1 port map( D => n2901, CK => CLK, Q => n52697, QN 
                           => n_2482);
   clk_r_REG16166_S1 : DFF_X1 port map( D => n2839, CK => CLK, Q => n52696, QN 
                           => n_2483);
   clk_r_REG16168_S1 : DFF_X1 port map( D => n2838, CK => CLK, Q => n52695, QN 
                           => n_2484);
   clk_r_REG16104_S1 : DFF_X1 port map( D => n2806, CK => CLK, Q => n52694, QN 
                           => n_2485);
   clk_r_REG16170_S1 : DFF_X1 port map( D => n2837, CK => CLK, Q => n52693, QN 
                           => n_2486);
   clk_r_REG16106_S1 : DFF_X1 port map( D => n2805, CK => CLK, Q => n52692, QN 
                           => n_2487);
   clk_r_REG16172_S1 : DFF_X1 port map( D => n2836, CK => CLK, Q => n52691, QN 
                           => n_2488);
   clk_r_REG16108_S1 : DFF_X1 port map( D => n2804, CK => CLK, Q => n52690, QN 
                           => n_2489);
   clk_r_REG16174_S1 : DFF_X1 port map( D => n2835, CK => CLK, Q => n52689, QN 
                           => n_2490);
   clk_r_REG16110_S1 : DFF_X1 port map( D => n2803, CK => CLK, Q => n52688, QN 
                           => n_2491);
   clk_r_REG14790_S1 : DFF_X1 port map( D => n3321, CK => CLK, Q => n52687, QN 
                           => n_2492);
   clk_r_REG14792_S1 : DFF_X1 port map( D => n3320, CK => CLK, Q => n52686, QN 
                           => n_2493);
   clk_r_REG15653_S1 : DFF_X1 port map( D => n3032, CK => CLK, Q => n52685, QN 
                           => n_2494);
   clk_r_REG14794_S1 : DFF_X1 port map( D => n3319, CK => CLK, Q => n52684, QN 
                           => n_2495);
   clk_r_REG14796_S1 : DFF_X1 port map( D => n3318, CK => CLK, Q => n52683, QN 
                           => n_2496);
   clk_r_REG15139_S1 : DFF_X1 port map( D => n3161, CK => CLK, Q => n52682, QN 
                           => n_2497);
   clk_r_REG15141_S1 : DFF_X1 port map( D => n3160, CK => CLK, Q => n52681, QN 
                           => n_2498);
   clk_r_REG16412_S1 : DFF_X1 port map( D => n3099, CK => CLK, Q => n52680, QN 
                           => n_2499);
   clk_r_REG14926_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n52679, QN 
                           => n_2500);
   clk_r_REG16414_S1 : DFF_X1 port map( D => n3098, CK => CLK, Q => n52678, QN 
                           => n_2501);
   clk_r_REG15272_S1 : DFF_X1 port map( D => n3256, CK => CLK, Q => n52677, QN 
                           => n_2502);
   clk_r_REG14928_S1 : DFF_X1 port map( D => n3290, CK => CLK, Q => n52676, QN 
                           => n_2503);
   clk_r_REG15655_S1 : DFF_X1 port map( D => n3031, CK => CLK, Q => n52675, QN 
                           => n_2504);
   clk_r_REG15523_S1 : DFF_X1 port map( D => n2969, CK => CLK, Q => n52674, QN 
                           => n_2505);
   clk_r_REG15657_S1 : DFF_X1 port map( D => n3030, CK => CLK, Q => n52673, QN 
                           => n_2506);
   clk_r_REG14860_S1 : DFF_X1 port map( D => n3482, CK => CLK, Q => n52672, QN 
                           => n_2507);
   clk_r_REG14862_S1 : DFF_X1 port map( D => n3481, CK => CLK, Q => n52671, QN 
                           => n_2508);
   clk_r_REG15579_S1 : DFF_X1 port map( D => n3005, CK => CLK, Q => n52670, QN 
                           => n_2509);
   clk_r_REG15069_S1 : DFF_X1 port map( D => n3066, CK => CLK, Q => n52669, QN 
                           => n_2510);
   clk_r_REG14390_S1 : DFF_X1 port map( D => n3418, CK => CLK, Q => n52668, QN 
                           => n_2511);
   clk_r_REG15002_S1 : DFF_X1 port map( D => n3514, CK => CLK, Q => n52667, QN 
                           => n_2512);
   clk_r_REG15331_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n52666, QN 
                           => n_2513);
   clk_r_REG14720_S1 : DFF_X1 port map( D => n3450, CK => CLK, Q => n52665, QN 
                           => n_2514);
   clk_r_REG15405_S1 : DFF_X1 port map( D => n2900, CK => CLK, Q => n52664, QN 
                           => n_2515);
   clk_r_REG14644_S1 : DFF_X1 port map( D => n3386, CK => CLK, Q => n52663, QN 
                           => n_2516);
   clk_r_REG14798_S1 : DFF_X1 port map( D => n3317, CK => CLK, Q => n52662, QN 
                           => n_2517);
   clk_r_REG15581_S1 : DFF_X1 port map( D => n3004, CK => CLK, Q => n52661, QN 
                           => n_2518);
   clk_r_REG14864_S1 : DFF_X1 port map( D => n3480, CK => CLK, Q => n52660, QN 
                           => n_2519);
   clk_r_REG15004_S1 : DFF_X1 port map( D => n3513, CK => CLK, Q => n52659, QN 
                           => n_2520);
   clk_r_REG14392_S1 : DFF_X1 port map( D => n3417, CK => CLK, Q => n52658, QN 
                           => n_2521);
   clk_r_REG15583_S1 : DFF_X1 port map( D => n3003, CK => CLK, Q => n52657, QN 
                           => n_2522);
   clk_r_REG15407_S1 : DFF_X1 port map( D => n2899, CK => CLK, Q => n52656, QN 
                           => n_2523);
   clk_r_REG15333_S1 : DFF_X1 port map( D => n3353, CK => CLK, Q => n52655, QN 
                           => n_2524);
   clk_r_REG14646_S1 : DFF_X1 port map( D => n3385, CK => CLK, Q => n52654, QN 
                           => n_2525);
   clk_r_REG15071_S1 : DFF_X1 port map( D => n3065, CK => CLK, Q => n52653, QN 
                           => n_2526);
   clk_r_REG14866_S1 : DFF_X1 port map( D => n3479, CK => CLK, Q => n52652, QN 
                           => n_2527);
   clk_r_REG14800_S1 : DFF_X1 port map( D => n3316, CK => CLK, Q => n52651, QN 
                           => n_2528);
   clk_r_REG14722_S1 : DFF_X1 port map( D => n3449, CK => CLK, Q => n52650, QN 
                           => n_2529);
   clk_r_REG15585_S1 : DFF_X1 port map( D => n3002, CK => CLK, Q => n52649, QN 
                           => n_2530);
   clk_r_REG14930_S1 : DFF_X1 port map( D => n3289, CK => CLK, Q => n52648, QN 
                           => n_2531);
   clk_r_REG15274_S1 : DFF_X1 port map( D => n3255, CK => CLK, Q => n52647, QN 
                           => n_2532);
   clk_r_REG15587_S1 : DFF_X1 port map( D => n3001, CK => CLK, Q => n52646, QN 
                           => n_2533);
   clk_r_REG15589_S1 : DFF_X1 port map( D => n3000, CK => CLK, Q => n52645, QN 
                           => n_2534);
   clk_r_REG16645_S1 : DFF_X1 port map( D => n3543, CK => CLK, Q => n52644, QN 
                           => n_2535);
   clk_r_REG16647_S1 : DFF_X1 port map( D => n3542, CK => CLK, Q => n52643, QN 
                           => n_2536);
   clk_r_REG14868_S1 : DFF_X1 port map( D => n3478, CK => CLK, Q => n52642, QN 
                           => n_2537);
   clk_r_REG14648_S1 : DFF_X1 port map( D => n3384, CK => CLK, Q => n52641, QN 
                           => n_2538);
   clk_r_REG14724_S1 : DFF_X1 port map( D => n3448, CK => CLK, Q => n52640, QN 
                           => n_2539);
   clk_r_REG15335_S1 : DFF_X1 port map( D => n3352, CK => CLK, Q => n52639, QN 
                           => n_2540);
   clk_r_REG14650_S1 : DFF_X1 port map( D => n3383, CK => CLK, Q => n52638, QN 
                           => n_2541);
   clk_r_REG15006_S1 : DFF_X1 port map( D => n3512, CK => CLK, Q => n52637, QN 
                           => n_2542);
   clk_r_REG15337_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n52636, QN 
                           => n_2543);
   clk_r_REG15339_S1 : DFF_X1 port map( D => n3350, CK => CLK, Q => n52635, QN 
                           => n_2544);
   clk_r_REG14394_S1 : DFF_X1 port map( D => n3416, CK => CLK, Q => n52634, QN 
                           => n_2545);
   clk_r_REG15008_S1 : DFF_X1 port map( D => n3511, CK => CLK, Q => n52633, QN 
                           => n_2546);
   clk_r_REG14396_S1 : DFF_X1 port map( D => n3415, CK => CLK, Q => n52632, QN 
                           => n_2547);
   clk_r_REG15591_S1 : DFF_X1 port map( D => n2999, CK => CLK, Q => n52631, QN 
                           => n_2548);
   clk_r_REG15073_S1 : DFF_X1 port map( D => n3064, CK => CLK, Q => n52630, QN 
                           => n_2549);
   clk_r_REG14726_S1 : DFF_X1 port map( D => n3447, CK => CLK, Q => n52629, QN 
                           => n_2550);
   clk_r_REG15075_S1 : DFF_X1 port map( D => n3063, CK => CLK, Q => n52628, QN 
                           => n_2551);
   clk_r_REG15010_S1 : DFF_X1 port map( D => n3510, CK => CLK, Q => n52627, QN 
                           => n_2552);
   clk_r_REG14802_S1 : DFF_X1 port map( D => n3315, CK => CLK, Q => n52626, QN 
                           => n_2553);
   clk_r_REG14652_S1 : DFF_X1 port map( D => n3382, CK => CLK, Q => n52625, QN 
                           => n_2554);
   clk_r_REG14804_S1 : DFF_X1 port map( D => n3314, CK => CLK, Q => n52624, QN 
                           => n_2555);
   clk_r_REG14728_S1 : DFF_X1 port map( D => n3446, CK => CLK, Q => n52623, QN 
                           => n_2556);
   clk_r_REG14806_S1 : DFF_X1 port map( D => n3313, CK => CLK, Q => n52622, QN 
                           => n_2557);
   clk_r_REG14398_S1 : DFF_X1 port map( D => n3414, CK => CLK, Q => n52621, QN 
                           => n_2558);
   clk_r_REG15593_S1 : DFF_X1 port map( D => n2998, CK => CLK, Q => n52620, QN 
                           => n_2559);
   clk_r_REG15202_S1 : DFF_X1 port map( D => n3195, CK => CLK, Q => n52619, QN 
                           => n_2560);
   clk_r_REG15143_S1 : DFF_X1 port map( D => n3159, CK => CLK, Q => n52618, QN 
                           => n_2561);
   clk_r_REG16477_S1 : DFF_X1 port map( D => n3131, CK => CLK, Q => n52617, QN 
                           => n_2562);
   clk_r_REG16416_S1 : DFF_X1 port map( D => n3097, CK => CLK, Q => n52616, QN 
                           => n_2563);
   clk_r_REG15077_S1 : DFF_X1 port map( D => n3062, CK => CLK, Q => n52615, QN 
                           => n_2564);
   clk_r_REG15525_S1 : DFF_X1 port map( D => n2968, CK => CLK, Q => n52614, QN 
                           => n_2565);
   clk_r_REG16226_S1 : DFF_X1 port map( D => n2873, CK => CLK, Q => n52613, QN 
                           => n_2566);
   clk_r_REG16228_S1 : DFF_X1 port map( D => n2872, CK => CLK, Q => n52612, QN 
                           => n_2567);
   clk_r_REG16230_S1 : DFF_X1 port map( D => n2871, CK => CLK, Q => n52611, QN 
                           => n_2568);
   clk_r_REG16232_S1 : DFF_X1 port map( D => n2870, CK => CLK, Q => n52610, QN 
                           => n_2569);
   clk_r_REG15481_S1 : DFF_X1 port map( D => n2937, CK => CLK, Q => n52609, QN 
                           => n_2570);
   clk_r_REG15409_S1 : DFF_X1 port map( D => n2898, CK => CLK, Q => n52608, QN 
                           => n_2571);
   clk_r_REG16176_S1 : DFF_X1 port map( D => n2834, CK => CLK, Q => n52607, QN 
                           => n_2572);
   clk_r_REG16112_S1 : DFF_X1 port map( D => n2802, CK => CLK, Q => n52606, QN 
                           => n_2573);
   clk_r_REG16234_S1 : DFF_X1 port map( D => n2869, CK => CLK, Q => n52605, QN 
                           => n_2574);
   clk_r_REG16114_S1 : DFF_X1 port map( D => n2801, CK => CLK, Q => n52604, QN 
                           => n_2575);
   clk_r_REG16178_S1 : DFF_X1 port map( D => n2833, CK => CLK, Q => n52603, QN 
                           => n_2576);
   clk_r_REG15411_S1 : DFF_X1 port map( D => n2897, CK => CLK, Q => n52602, QN 
                           => n_2577);
   clk_r_REG15483_S1 : DFF_X1 port map( D => n2936, CK => CLK, Q => n52601, QN 
                           => n_2578);
   clk_r_REG15527_S1 : DFF_X1 port map( D => n2967, CK => CLK, Q => n52600, QN 
                           => n_2579);
   clk_r_REG16418_S1 : DFF_X1 port map( D => n3096, CK => CLK, Q => n52599, QN 
                           => n_2580);
   clk_r_REG16479_S1 : DFF_X1 port map( D => n3130, CK => CLK, Q => n52598, QN 
                           => n_2581);
   clk_r_REG15145_S1 : DFF_X1 port map( D => n3158, CK => CLK, Q => n52597, QN 
                           => n_2582);
   clk_r_REG15204_S1 : DFF_X1 port map( D => n3194, CK => CLK, Q => n52596, QN 
                           => n_2583);
   clk_r_REG14932_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n52595, QN 
                           => n_2584);
   clk_r_REG15276_S1 : DFF_X1 port map( D => n3254, CK => CLK, Q => n52594, QN 
                           => n_2585);
   clk_r_REG15206_S1 : DFF_X1 port map( D => n3193, CK => CLK, Q => n52593, QN 
                           => n_2586);
   clk_r_REG15278_S1 : DFF_X1 port map( D => n3253, CK => CLK, Q => n52592, QN 
                           => n_2587);
   clk_r_REG14934_S1 : DFF_X1 port map( D => n3287, CK => CLK, Q => n52591, QN 
                           => n_2588);
   clk_r_REG15147_S1 : DFF_X1 port map( D => n3157, CK => CLK, Q => n52590, QN 
                           => n_2589);
   clk_r_REG16481_S1 : DFF_X1 port map( D => n3129, CK => CLK, Q => n52589, QN 
                           => n_2590);
   clk_r_REG16420_S1 : DFF_X1 port map( D => n3095, CK => CLK, Q => n52588, QN 
                           => n_2591);
   clk_r_REG15079_S1 : DFF_X1 port map( D => n3061, CK => CLK, Q => n52587, QN 
                           => n_2592);
   clk_r_REG16651_S1 : DFF_X1 port map( D => n3540, CK => CLK, Q => n52586, QN 
                           => n_2593);
   clk_r_REG16236_S1 : DFF_X1 port map( D => n2868, CK => CLK, Q => n52585, QN 
                           => n_2594);
   clk_r_REG15280_S1 : DFF_X1 port map( D => n3252, CK => CLK, Q => n52584, QN 
                           => n_2595);
   clk_r_REG15529_S1 : DFF_X1 port map( D => n2966, CK => CLK, Q => n52583, QN 
                           => n_2596);
   clk_r_REG15208_S1 : DFF_X1 port map( D => n3192, CK => CLK, Q => n52582, QN 
                           => n_2597);
   clk_r_REG16483_S1 : DFF_X1 port map( D => n3128, CK => CLK, Q => n52581, QN 
                           => n_2598);
   clk_r_REG16422_S1 : DFF_X1 port map( D => n3094, CK => CLK, Q => n52580, QN 
                           => n_2599);
   clk_r_REG15595_S1 : DFF_X1 port map( D => n2997, CK => CLK, Q => n52579, QN 
                           => n_2600);
   clk_r_REG15081_S1 : DFF_X1 port map( D => n3060, CK => CLK, Q => n52578, QN 
                           => n_2601);
   clk_r_REG15485_S1 : DFF_X1 port map( D => n2935, CK => CLK, Q => n52577, QN 
                           => n_2602);
   clk_r_REG15531_S1 : DFF_X1 port map( D => n2965, CK => CLK, Q => n52576, QN 
                           => n_2603);
   clk_r_REG15597_S1 : DFF_X1 port map( D => n2996, CK => CLK, Q => n52575, QN 
                           => n_2604);
   clk_r_REG15659_S1 : DFF_X1 port map( D => n3029, CK => CLK, Q => n52574, QN 
                           => n_2605);
   clk_r_REG15083_S1 : DFF_X1 port map( D => n3059, CK => CLK, Q => n52573, QN 
                           => n_2606);
   clk_r_REG15599_S1 : DFF_X1 port map( D => n2995, CK => CLK, Q => n52572, QN 
                           => n_2607);
   clk_r_REG16424_S1 : DFF_X1 port map( D => n3093, CK => CLK, Q => n52571, QN 
                           => n_2608);
   clk_r_REG16485_S1 : DFF_X1 port map( D => n3127, CK => CLK, Q => n52570, QN 
                           => n_2609);
   clk_r_REG15149_S1 : DFF_X1 port map( D => n3156, CK => CLK, Q => n52569, QN 
                           => n_2610);
   clk_r_REG15210_S1 : DFF_X1 port map( D => n3191, CK => CLK, Q => n52568, QN 
                           => n_2611);
   clk_r_REG15282_S1 : DFF_X1 port map( D => n3251, CK => CLK, Q => n52567, QN 
                           => n_2612);
   clk_r_REG14936_S1 : DFF_X1 port map( D => n3286, CK => CLK, Q => n52566, QN 
                           => n_2613);
   clk_r_REG15085_S1 : DFF_X1 port map( D => n3058, CK => CLK, Q => n52565, QN 
                           => n_2614);
   clk_r_REG14938_S1 : DFF_X1 port map( D => n3285, CK => CLK, Q => n52564, QN 
                           => n_2615);
   clk_r_REG14400_S1 : DFF_X1 port map( D => n3413, CK => CLK, Q => n52563, QN 
                           => n_2616);
   clk_r_REG15661_S1 : DFF_X1 port map( D => n3028, CK => CLK, Q => n52562, QN 
                           => n_2617);
   clk_r_REG14870_S1 : DFF_X1 port map( D => n3477, CK => CLK, Q => n52561, QN 
                           => n_2618);
   clk_r_REG16487_S1 : DFF_X1 port map( D => n3126, CK => CLK, Q => n52560, QN 
                           => n_2619);
   clk_r_REG16426_S1 : DFF_X1 port map( D => n3092, CK => CLK, Q => n52559, QN 
                           => n_2620);
   clk_r_REG15212_S1 : DFF_X1 port map( D => n3190, CK => CLK, Q => n52558, QN 
                           => n_2621);
   clk_r_REG16238_S1 : DFF_X1 port map( D => n2867, CK => CLK, Q => n52557, QN 
                           => n_2622);
   clk_r_REG14730_S1 : DFF_X1 port map( D => n3445, CK => CLK, Q => n52556, QN 
                           => n_2623);
   clk_r_REG15151_S1 : DFF_X1 port map( D => n3155, CK => CLK, Q => n52555, QN 
                           => n_2624);
   clk_r_REG15012_S1 : DFF_X1 port map( D => n3509, CK => CLK, Q => n52554, QN 
                           => n_2625);
   clk_r_REG15487_S1 : DFF_X1 port map( D => n2934, CK => CLK, Q => n52553, QN 
                           => n_2626);
   clk_r_REG15087_S1 : DFF_X1 port map( D => n3057, CK => CLK, Q => n52552, QN 
                           => n_2627);
   clk_r_REG15533_S1 : DFF_X1 port map( D => n2964, CK => CLK, Q => n52551, QN 
                           => n_2628);
   clk_r_REG15153_S1 : DFF_X1 port map( D => n3154, CK => CLK, Q => n52550, QN 
                           => n_2629);
   clk_r_REG16489_S1 : DFF_X1 port map( D => n3125, CK => CLK, Q => n52549, QN 
                           => n_2630);
   clk_r_REG16428_S1 : DFF_X1 port map( D => n3091, CK => CLK, Q => n52548, QN 
                           => n_2631);
   clk_r_REG15663_S1 : DFF_X1 port map( D => n3027, CK => CLK, Q => n52547, QN 
                           => n_2632);
   clk_r_REG14940_S1 : DFF_X1 port map( D => n3284, CK => CLK, Q => n52546, QN 
                           => n_2633);
   clk_r_REG15601_S1 : DFF_X1 port map( D => n2994, CK => CLK, Q => n52545, QN 
                           => n_2634);
   clk_r_REG15284_S1 : DFF_X1 port map( D => n3250, CK => CLK, Q => n52544, QN 
                           => n_2635);
   clk_r_REG15214_S1 : DFF_X1 port map( D => n3189, CK => CLK, Q => n52543, QN 
                           => n_2636);
   clk_r_REG14942_S1 : DFF_X1 port map( D => n3283, CK => CLK, Q => n52542, QN 
                           => n_2637);
   clk_r_REG15603_S1 : DFF_X1 port map( D => n2993, CK => CLK, Q => n52541, QN 
                           => n_2638);
   clk_r_REG15535_S1 : DFF_X1 port map( D => n2963, CK => CLK, Q => n52540, QN 
                           => n_2639);
   clk_r_REG15489_S1 : DFF_X1 port map( D => n2933, CK => CLK, Q => n52539, QN 
                           => n_2640);
   clk_r_REG16240_S1 : DFF_X1 port map( D => n2866, CK => CLK, Q => n52538, QN 
                           => n_2641);
   clk_r_REG14944_S1 : DFF_X1 port map( D => n3282, CK => CLK, Q => n52537, QN 
                           => n_2642);
   clk_r_REG16653_S1 : DFF_X1 port map( D => n3539, CK => CLK, Q => n52536, QN 
                           => n_2643);
   clk_r_REG15341_S1 : DFF_X1 port map( D => n3349, CK => CLK, Q => n52535, QN 
                           => n_2644);
   clk_r_REG15665_S1 : DFF_X1 port map( D => n3026, CK => CLK, Q => n52534, QN 
                           => n_2645);
   clk_r_REG14732_S1 : DFF_X1 port map( D => n3444, CK => CLK, Q => n52533, QN 
                           => n_2646);
   clk_r_REG15216_S1 : DFF_X1 port map( D => n3188, CK => CLK, Q => n52532, QN 
                           => n_2647);
   clk_r_REG15491_S1 : DFF_X1 port map( D => n2932, CK => CLK, Q => n52531, QN 
                           => n_2648);
   clk_r_REG14654_S1 : DFF_X1 port map( D => n3381, CK => CLK, Q => n52530, QN 
                           => n_2649);
   clk_r_REG15343_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n52529, QN 
                           => n_2650);
   clk_r_REG15493_S1 : DFF_X1 port map( D => n2931, CK => CLK, Q => n52528, QN 
                           => n_2651);
   clk_r_REG15537_S1 : DFF_X1 port map( D => n2962, CK => CLK, Q => n52527, QN 
                           => n_2652);
   clk_r_REG15495_S1 : DFF_X1 port map( D => n2930, CK => CLK, Q => n52526, QN 
                           => n_2653);
   clk_r_REG16491_S1 : DFF_X1 port map( D => n3124, CK => CLK, Q => n52525, QN 
                           => n_2654);
   clk_r_REG16493_S1 : DFF_X1 port map( D => n3123, CK => CLK, Q => n52524, QN 
                           => n_2655);
   clk_r_REG16430_S1 : DFF_X1 port map( D => n3090, CK => CLK, Q => n52523, QN 
                           => n_2656);
   clk_r_REG15667_S1 : DFF_X1 port map( D => n3025, CK => CLK, Q => n52522, QN 
                           => n_2657);
   clk_r_REG16242_S1 : DFF_X1 port map( D => n2865, CK => CLK, Q => n52521, QN 
                           => n_2658);
   clk_r_REG15155_S1 : DFF_X1 port map( D => n3153, CK => CLK, Q => n52520, QN 
                           => n_2659);
   clk_r_REG15218_S1 : DFF_X1 port map( D => n3187, CK => CLK, Q => n52519, QN 
                           => n_2660);
   clk_r_REG16495_S1 : DFF_X1 port map( D => n3122, CK => CLK, Q => n52518, QN 
                           => n_2661);
   clk_r_REG14656_S1 : DFF_X1 port map( D => n3380, CK => CLK, Q => n52517, QN 
                           => n_2662);
   clk_r_REG15220_S1 : DFF_X1 port map( D => n3186, CK => CLK, Q => n52516, QN 
                           => n_2663);
   clk_r_REG14946_S1 : DFF_X1 port map( D => n3281, CK => CLK, Q => n52515, QN 
                           => n_2664);
   clk_r_REG16497_S1 : DFF_X1 port map( D => n3121, CK => CLK, Q => n52514, QN 
                           => n_2665);
   clk_r_REG16559_S1 : DFF_X1 port map( D => n3218, CK => CLK, Q => n52513, QN 
                           => n_2666);
   clk_r_REG15286_S1 : DFF_X1 port map( D => n3249, CK => CLK, Q => n52512, QN 
                           => n_2667);
   clk_r_REG16561_S1 : DFF_X1 port map( D => n3217, CK => CLK, Q => n52511, QN 
                           => n_2668);
   clk_r_REG16655_S1 : DFF_X1 port map( D => n3538, CK => CLK, Q => n52510, QN 
                           => n_2669);
   clk_r_REG15539_S1 : DFF_X1 port map( D => n2961, CK => CLK, Q => n52509, QN 
                           => n_2670);
   clk_r_REG14872_S1 : DFF_X1 port map( D => n3476, CK => CLK, Q => n52508, QN 
                           => n_2671);
   clk_r_REG14734_S1 : DFF_X1 port map( D => n3443, CK => CLK, Q => n52507, QN 
                           => n_2672);
   clk_r_REG15014_S1 : DFF_X1 port map( D => n3508, CK => CLK, Q => n52506, QN 
                           => n_2673);
   clk_r_REG14658_S1 : DFF_X1 port map( D => n3379, CK => CLK, Q => n52505, QN 
                           => n_2674);
   clk_r_REG16657_S1 : DFF_X1 port map( D => n3537, CK => CLK, Q => n52504, QN 
                           => n_2675);
   clk_r_REG14736_S1 : DFF_X1 port map( D => n3442, CK => CLK, Q => n52503, QN 
                           => n_2676);
   clk_r_REG14874_S1 : DFF_X1 port map( D => n3475, CK => CLK, Q => n52502, QN 
                           => n_2677);
   clk_r_REG15345_S1 : DFF_X1 port map( D => n3347, CK => CLK, Q => n52501, QN 
                           => n_2678);
   clk_r_REG15497_S1 : DFF_X1 port map( D => n2929, CK => CLK, Q => n52500, QN 
                           => n_2679);
   clk_r_REG14738_S1 : DFF_X1 port map( D => n3441, CK => CLK, Q => n52499, QN 
                           => n_2680);
   clk_r_REG15347_S1 : DFF_X1 port map( D => n3346, CK => CLK, Q => n52498, QN 
                           => n_2681);
   clk_r_REG14402_S1 : DFF_X1 port map( D => n3412, CK => CLK, Q => n52497, QN 
                           => n_2682);
   clk_r_REG14404_S1 : DFF_X1 port map( D => n3411, CK => CLK, Q => n52496, QN 
                           => n_2683);
   clk_r_REG14876_S1 : DFF_X1 port map( D => n3474, CK => CLK, Q => n52495, QN 
                           => n_2684);
   clk_r_REG14660_S1 : DFF_X1 port map( D => n3378, CK => CLK, Q => n52494, QN 
                           => n_2685);
   clk_r_REG14406_S1 : DFF_X1 port map( D => n3410, CK => CLK, Q => n52493, QN 
                           => n_2686);
   clk_r_REG14662_S1 : DFF_X1 port map( D => n3377, CK => CLK, Q => n52492, QN 
                           => n_2687);
   clk_r_REG14408_S1 : DFF_X1 port map( D => n3409, CK => CLK, Q => n52491, QN 
                           => n_2688);
   clk_r_REG15016_S1 : DFF_X1 port map( D => n3507, CK => CLK, Q => n52490, QN 
                           => n_2689);
   clk_r_REG15222_S1 : DFF_X1 port map( D => n3185, CK => CLK, Q => n52489, QN 
                           => n_2690);
   clk_r_REG15018_S1 : DFF_X1 port map( D => n3506, CK => CLK, Q => n52488, QN 
                           => n_2691);
   clk_r_REG14878_S1 : DFF_X1 port map( D => n3473, CK => CLK, Q => n52487, QN 
                           => n_2692);
   clk_r_REG15020_S1 : DFF_X1 port map( D => n3505, CK => CLK, Q => n52486, QN 
                           => n_2693);
   clk_r_REG16432_S1 : DFF_X1 port map( D => n3089, CK => CLK, Q => n52485, QN 
                           => n_2694);
   clk_r_REG16929_S7 : DFFS_X1 port map( D => n3567, CK => CLK, SN => RESET_BAR
                           , Q => n52484, QN => n_2695);
   clk_r_REG16999_S7 : DFFS_X1 port map( D => n3558, CK => CLK, SN => RESET_BAR
                           , Q => n52483, QN => n_2696);
   clk_r_REG16773_S2 : DFFR_X1 port map( D => n40643, CK => CLK, RN => 
                           RESET_BAR, Q => n52476, QN => n_2697);
   clk_r_REG16774_S3 : DFFR_X1 port map( D => n52476, CK => CLK, RN => 
                           RESET_BAR, Q => n52475, QN => n_2698);
   clk_r_REG16775_S4 : DFFR_X1 port map( D => n52475, CK => CLK, RN => 
                           RESET_BAR, Q => n52474, QN => n_2699);
   clk_r_REG16770_S2 : DFFR_X1 port map( D => n40639, CK => CLK, RN => 
                           RESET_BAR, Q => n52472, QN => n_2700);
   clk_r_REG16771_S3 : DFFR_X1 port map( D => n52472, CK => CLK, RN => 
                           RESET_BAR, Q => n52471, QN => n_2701);
   clk_r_REG16772_S4 : DFFR_X1 port map( D => n52471, CK => CLK, RN => 
                           RESET_BAR, Q => n52470, QN => n_2702);
   clk_r_REG16761_S2 : DFFR_X1 port map( D => n40633, CK => CLK, RN => 
                           RESET_BAR, Q => n52466, QN => n_2703);
   clk_r_REG16762_S3 : DFFR_X1 port map( D => n52466, CK => CLK, RN => 
                           RESET_BAR, Q => n52465, QN => n_2704);
   clk_r_REG16763_S4 : DFFR_X1 port map( D => n52465, CK => CLK, RN => 
                           RESET_BAR, Q => n52464, QN => n_2705);
   clk_r_REG16758_S2 : DFFR_X1 port map( D => n40629, CK => CLK, RN => 
                           RESET_BAR, Q => n52462, QN => n_2706);
   clk_r_REG16759_S3 : DFFR_X1 port map( D => n52462, CK => CLK, RN => 
                           RESET_BAR, Q => n52461, QN => n_2707);
   clk_r_REG16760_S4 : DFFR_X1 port map( D => n52461, CK => CLK, RN => 
                           RESET_BAR, Q => n52460, QN => n_2708);
   clk_r_REG16927_S7 : DFFR_X1 port map( D => n47429, CK => CLK, RN => 
                           RESET_BAR, Q => n52434, QN => n_2709);
   clk_r_REG16911_S7 : DFFR_X1 port map( D => n49092, CK => CLK, RN => 
                           RESET_BAR, Q => n52433, QN => n_2710);
   clk_r_REG16909_S7 : DFFR_X1 port map( D => n49093, CK => CLK, RN => 
                           RESET_BAR, Q => n52432, QN => n_2711);
   clk_r_REG16907_S7 : DFFR_X1 port map( D => n49094, CK => CLK, RN => 
                           RESET_BAR, Q => n52431, QN => n_2712);
   clk_r_REG16925_S7 : DFFR_X1 port map( D => n49087, CK => CLK, RN => 
                           RESET_BAR, Q => n52430, QN => n_2713);
   clk_r_REG16905_S7 : DFFR_X1 port map( D => n49089, CK => CLK, RN => 
                           RESET_BAR, Q => n52429, QN => n_2714);
   clk_r_REG16903_S7 : DFFR_X1 port map( D => n49091, CK => CLK, RN => 
                           RESET_BAR, Q => n52428, QN => n_2715);
   clk_r_REG16921_S7 : DFFR_X1 port map( D => n49086, CK => CLK, RN => 
                           RESET_BAR, Q => n52426, QN => n_2716);
   clk_r_REG16899_S7 : DFFR_X1 port map( D => n47428, CK => CLK, RN => 
                           RESET_BAR, Q => n52424, QN => n_2717);
   clk_r_REG16897_S7 : DFFR_X1 port map( D => n40592, CK => CLK, RN => 
                           RESET_BAR, Q => n52423, QN => n_2718);
   clk_r_REG16919_S7 : DFFR_X1 port map( D => n40591, CK => CLK, RN => 
                           RESET_BAR, Q => n52422, QN => n_2719);
   clk_r_REG16917_S7 : DFFR_X1 port map( D => n49085, CK => CLK, RN => 
                           RESET_BAR, Q => n52421, QN => n_2720);
   clk_r_REG16915_S7 : DFFR_X1 port map( D => n40589, CK => CLK, RN => 
                           RESET_BAR, Q => n52420, QN => n_2721);
   clk_r_REG16913_S7 : DFFR_X1 port map( D => n40588, CK => CLK, RN => 
                           RESET_BAR, Q => n52419, QN => n_2722);
   clk_r_REG16889_S7 : DFFR_X1 port map( D => n40587, CK => CLK, RN => 
                           RESET_BAR, Q => n52418, QN => n_2723);
   clk_r_REG16839_S7 : DFFR_X1 port map( D => n40586, CK => CLK, RN => 
                           RESET_BAR, Q => n52417, QN => n_2724);
   clk_r_REG16887_S7 : DFFR_X1 port map( D => n40585, CK => CLK, RN => 
                           RESET_BAR, Q => n52416, QN => n_2725);
   clk_r_REG16854_S7 : DFFR_X1 port map( D => n40584, CK => CLK, RN => 
                           RESET_BAR, Q => n52415, QN => n_2726);
   clk_r_REG16861_S7 : DFFR_X1 port map( D => n40583, CK => CLK, RN => 
                           RESET_BAR, Q => n52414, QN => n_2727);
   clk_r_REG16875_S7 : DFFR_X1 port map( D => n40582, CK => CLK, RN => 
                           RESET_BAR, Q => n52413, QN => n_2728);
   clk_r_REG16882_S7 : DFFR_X1 port map( D => n40581, CK => CLK, RN => 
                           RESET_BAR, Q => n52412, QN => n_2729);
   clk_r_REG16852_S7 : DFFR_X1 port map( D => n40580, CK => CLK, RN => 
                           RESET_BAR, Q => n52411, QN => n_2730);
   clk_r_REG16837_S7 : DFFR_X1 port map( D => n49095, CK => CLK, RN => 
                           RESET_BAR, Q => n52410, QN => n_2731);
   clk_r_REG16873_S7 : DFFR_X1 port map( D => n47430, CK => CLK, RN => 
                           RESET_BAR, Q => n52409, QN => n_2732);
   clk_r_REG16867_S7 : DFFR_X1 port map( D => n40577, CK => CLK, RN => 
                           RESET_BAR, Q => n52408, QN => n_2733);
   clk_r_REG16865_S7 : DFFR_X1 port map( D => n40576, CK => CLK, RN => 
                           RESET_BAR, Q => n52407, QN => n_2734);
   clk_r_REG16847_S7 : DFFR_X1 port map( D => n49096, CK => CLK, RN => 
                           RESET_BAR, Q => n52406, QN => n_2735);
   clk_r_REG16880_S7 : DFFR_X1 port map( D => n40574, CK => CLK, RN => 
                           RESET_BAR, Q => n52405, QN => n_2736);
   clk_r_REG16859_S7 : DFFR_X1 port map( D => n49097, CK => CLK, RN => 
                           RESET_BAR, Q => n52404, QN => n_2737);
   clk_r_REG16845_S7 : DFFR_X1 port map( D => n47431, CK => CLK, RN => 
                           RESET_BAR, Q => n52403, QN => n_2738);
   clk_r_REG16779_S2 : DFFS_X1 port map( D => n40561, CK => CLK, SN => 
                           RESET_BAR, Q => n52399, QN => n_2739);
   clk_r_REG16780_S3 : DFFS_X1 port map( D => n52399, CK => CLK, SN => 
                           RESET_BAR, Q => n52398, QN => n_2740);
   clk_r_REG16781_S4 : DFFS_X1 port map( D => n52398, CK => CLK, SN => 
                           RESET_BAR, Q => n52397, QN => n_2741);
   clk_r_REG16776_S2 : DFFR_X1 port map( D => n40558, CK => CLK, RN => 
                           RESET_BAR, Q => n52396, QN => n_2742);
   clk_r_REG16777_S3 : DFFR_X1 port map( D => n52396, CK => CLK, RN => 
                           RESET_BAR, Q => n52395, QN => n_2743);
   clk_r_REG16778_S4 : DFFR_X1 port map( D => n52395, CK => CLK, RN => 
                           RESET_BAR, Q => n52394, QN => n_2744);
   clk_r_REG16767_S2 : DFFR_X1 port map( D => n40555, CK => CLK, RN => 
                           RESET_BAR, Q => n52393, QN => n_2745);
   clk_r_REG16768_S3 : DFFR_X1 port map( D => n52393, CK => CLK, RN => 
                           RESET_BAR, Q => n52392, QN => n_2746);
   clk_r_REG16769_S4 : DFFR_X1 port map( D => n52392, CK => CLK, RN => 
                           RESET_BAR, Q => n52391, QN => n_2747);
   clk_r_REG16764_S2 : DFFR_X1 port map( D => n40552, CK => CLK, RN => 
                           RESET_BAR, Q => n52390, QN => n_2748);
   clk_r_REG16765_S3 : DFFR_X1 port map( D => n52390, CK => CLK, RN => 
                           RESET_BAR, Q => n52389, QN => n_2749);
   clk_r_REG16766_S4 : DFFR_X1 port map( D => n52389, CK => CLK, RN => 
                           RESET_BAR, Q => n52388, QN => n_2750);
   clk_r_REG16431_S1 : DFF_X1 port map( D => n3089, CK => CLK, Q => n_2751, QN 
                           => n52387);
   clk_r_REG15019_S1 : DFF_X1 port map( D => n3505, CK => CLK, Q => n_2752, QN 
                           => n52386);
   clk_r_REG15348_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n_2753, QN 
                           => n52385);
   clk_r_REG14877_S1 : DFF_X1 port map( D => n3473, CK => CLK, Q => n_2754, QN 
                           => n52384);
   clk_r_REG15017_S1 : DFF_X1 port map( D => n3506, CK => CLK, Q => n_2755, QN 
                           => n52383);
   clk_r_REG15221_S1 : DFF_X1 port map( D => n3185, CK => CLK, Q => n_2756, QN 
                           => n52382);
   clk_r_REG15015_S1 : DFF_X1 port map( D => n3507, CK => CLK, Q => n_2757, QN 
                           => n52381);
   clk_r_REG14407_S1 : DFF_X1 port map( D => n3409, CK => CLK, Q => n_2758, QN 
                           => n52380);
   clk_r_REG14661_S1 : DFF_X1 port map( D => n3377, CK => CLK, Q => n_2759, QN 
                           => n52379);
   clk_r_REG14405_S1 : DFF_X1 port map( D => n3410, CK => CLK, Q => n_2760, QN 
                           => n52378);
   clk_r_REG14659_S1 : DFF_X1 port map( D => n3378, CK => CLK, Q => n_2761, QN 
                           => n52377);
   clk_r_REG14875_S1 : DFF_X1 port map( D => n3474, CK => CLK, Q => n_2762, QN 
                           => n52376);
   clk_r_REG14403_S1 : DFF_X1 port map( D => n3411, CK => CLK, Q => n_2763, QN 
                           => n52375);
   clk_r_REG14401_S1 : DFF_X1 port map( D => n3412, CK => CLK, Q => n_2764, QN 
                           => n52374);
   clk_r_REG15346_S1 : DFF_X1 port map( D => n3346, CK => CLK, Q => n_2765, QN 
                           => n52373);
   clk_r_REG14737_S1 : DFF_X1 port map( D => n3441, CK => CLK, Q => n_2766, QN 
                           => n52372);
   clk_r_REG15496_S1 : DFF_X1 port map( D => n2929, CK => CLK, Q => n_2767, QN 
                           => n52371);
   clk_r_REG15344_S1 : DFF_X1 port map( D => n3347, CK => CLK, Q => n_2768, QN 
                           => n52370);
   clk_r_REG14873_S1 : DFF_X1 port map( D => n3475, CK => CLK, Q => n_2769, QN 
                           => n52369);
   clk_r_REG14735_S1 : DFF_X1 port map( D => n3442, CK => CLK, Q => n_2770, QN 
                           => n52368);
   clk_r_REG16656_S1 : DFF_X1 port map( D => n3537, CK => CLK, Q => n_2771, QN 
                           => n52367);
   clk_r_REG14657_S1 : DFF_X1 port map( D => n3379, CK => CLK, Q => n_2772, QN 
                           => n52366);
   clk_r_REG15013_S1 : DFF_X1 port map( D => n3508, CK => CLK, Q => n_2773, QN 
                           => n52365);
   clk_r_REG14733_S1 : DFF_X1 port map( D => n3443, CK => CLK, Q => n_2774, QN 
                           => n52364);
   clk_r_REG14871_S1 : DFF_X1 port map( D => n3476, CK => CLK, Q => n_2775, QN 
                           => n52363);
   clk_r_REG15538_S1 : DFF_X1 port map( D => n2961, CK => CLK, Q => n_2776, QN 
                           => n52362);
   clk_r_REG16654_S1 : DFF_X1 port map( D => n3538, CK => CLK, Q => n_2777, QN 
                           => n52361);
   clk_r_REG16560_S1 : DFF_X1 port map( D => n3217, CK => CLK, Q => n_2778, QN 
                           => n52360);
   clk_r_REG15285_S1 : DFF_X1 port map( D => n3249, CK => CLK, Q => n_2779, QN 
                           => n52359);
   clk_r_REG16558_S1 : DFF_X1 port map( D => n3218, CK => CLK, Q => n_2780, QN 
                           => n52358);
   clk_r_REG16496_S1 : DFF_X1 port map( D => n3121, CK => CLK, Q => n_2781, QN 
                           => n52357);
   clk_r_REG14945_S1 : DFF_X1 port map( D => n3281, CK => CLK, Q => n_2782, QN 
                           => n52356);
   clk_r_REG15219_S1 : DFF_X1 port map( D => n3186, CK => CLK, Q => n_2783, QN 
                           => n52355);
   clk_r_REG14655_S1 : DFF_X1 port map( D => n3380, CK => CLK, Q => n_2784, QN 
                           => n52354);
   clk_r_REG16494_S1 : DFF_X1 port map( D => n3122, CK => CLK, Q => n_2785, QN 
                           => n52353);
   clk_r_REG15217_S1 : DFF_X1 port map( D => n3187, CK => CLK, Q => n_2786, QN 
                           => n52352);
   clk_r_REG15154_S1 : DFF_X1 port map( D => n3153, CK => CLK, Q => n_2787, QN 
                           => n52351);
   clk_r_REG16241_S1 : DFF_X1 port map( D => n2865, CK => CLK, Q => n_2788, QN 
                           => n52350);
   clk_r_REG15666_S1 : DFF_X1 port map( D => n3025, CK => CLK, Q => n_2789, QN 
                           => n52349);
   clk_r_REG16429_S1 : DFF_X1 port map( D => n3090, CK => CLK, Q => n_2790, QN 
                           => n52348);
   clk_r_REG16492_S1 : DFF_X1 port map( D => n3123, CK => CLK, Q => n_2791, QN 
                           => n52347);
   clk_r_REG16490_S1 : DFF_X1 port map( D => n3124, CK => CLK, Q => n_2792, QN 
                           => n52346);
   clk_r_REG15494_S1 : DFF_X1 port map( D => n2930, CK => CLK, Q => n_2793, QN 
                           => n52345);
   clk_r_REG15536_S1 : DFF_X1 port map( D => n2962, CK => CLK, Q => n_2794, QN 
                           => n52344);
   clk_r_REG15492_S1 : DFF_X1 port map( D => n2931, CK => CLK, Q => n_2795, QN 
                           => n52343);
   clk_r_REG15342_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n_2796, QN 
                           => n52342);
   clk_r_REG14653_S1 : DFF_X1 port map( D => n3381, CK => CLK, Q => n_2797, QN 
                           => n52341);
   clk_r_REG15490_S1 : DFF_X1 port map( D => n2932, CK => CLK, Q => n_2798, QN 
                           => n52340);
   clk_r_REG15215_S1 : DFF_X1 port map( D => n3188, CK => CLK, Q => n_2799, QN 
                           => n52339);
   clk_r_REG14731_S1 : DFF_X1 port map( D => n3444, CK => CLK, Q => n_2800, QN 
                           => n52338);
   clk_r_REG15664_S1 : DFF_X1 port map( D => n3026, CK => CLK, Q => n_2801, QN 
                           => n52337);
   clk_r_REG15340_S1 : DFF_X1 port map( D => n3349, CK => CLK, Q => n_2802, QN 
                           => n52336);
   clk_r_REG16652_S1 : DFF_X1 port map( D => n3539, CK => CLK, Q => n_2803, QN 
                           => n52335);
   clk_r_REG14943_S1 : DFF_X1 port map( D => n3282, CK => CLK, Q => n_2804, QN 
                           => n52334);
   clk_r_REG16239_S1 : DFF_X1 port map( D => n2866, CK => CLK, Q => n_2805, QN 
                           => n52333);
   clk_r_REG15488_S1 : DFF_X1 port map( D => n2933, CK => CLK, Q => n_2806, QN 
                           => n52332);
   clk_r_REG15534_S1 : DFF_X1 port map( D => n2963, CK => CLK, Q => n_2807, QN 
                           => n52331);
   clk_r_REG15602_S1 : DFF_X1 port map( D => n2993, CK => CLK, Q => n_2808, QN 
                           => n52330);
   clk_r_REG14941_S1 : DFF_X1 port map( D => n3283, CK => CLK, Q => n_2809, QN 
                           => n52329);
   clk_r_REG15213_S1 : DFF_X1 port map( D => n3189, CK => CLK, Q => n_2810, QN 
                           => n52328);
   clk_r_REG15283_S1 : DFF_X1 port map( D => n3250, CK => CLK, Q => n_2811, QN 
                           => n52327);
   clk_r_REG15600_S1 : DFF_X1 port map( D => n2994, CK => CLK, Q => n_2812, QN 
                           => n52326);
   clk_r_REG14939_S1 : DFF_X1 port map( D => n3284, CK => CLK, Q => n_2813, QN 
                           => n52325);
   clk_r_REG15662_S1 : DFF_X1 port map( D => n3027, CK => CLK, Q => n_2814, QN 
                           => n52324);
   clk_r_REG16427_S1 : DFF_X1 port map( D => n3091, CK => CLK, Q => n_2815, QN 
                           => n52323);
   clk_r_REG16488_S1 : DFF_X1 port map( D => n3125, CK => CLK, Q => n_2816, QN 
                           => n52322);
   clk_r_REG15152_S1 : DFF_X1 port map( D => n3154, CK => CLK, Q => n_2817, QN 
                           => n52321);
   clk_r_REG15532_S1 : DFF_X1 port map( D => n2964, CK => CLK, Q => n_2818, QN 
                           => n52320);
   clk_r_REG15086_S1 : DFF_X1 port map( D => n3057, CK => CLK, Q => n_2819, QN 
                           => n52319);
   clk_r_REG15486_S1 : DFF_X1 port map( D => n2934, CK => CLK, Q => n_2820, QN 
                           => n52318);
   clk_r_REG15011_S1 : DFF_X1 port map( D => n3509, CK => CLK, Q => n_2821, QN 
                           => n52317);
   clk_r_REG15150_S1 : DFF_X1 port map( D => n3155, CK => CLK, Q => n_2822, QN 
                           => n52316);
   clk_r_REG14729_S1 : DFF_X1 port map( D => n3445, CK => CLK, Q => n_2823, QN 
                           => n52315);
   clk_r_REG16237_S1 : DFF_X1 port map( D => n2867, CK => CLK, Q => n_2824, QN 
                           => n52314);
   clk_r_REG15211_S1 : DFF_X1 port map( D => n3190, CK => CLK, Q => n_2825, QN 
                           => n52313);
   clk_r_REG16425_S1 : DFF_X1 port map( D => n3092, CK => CLK, Q => n_2826, QN 
                           => n52312);
   clk_r_REG16486_S1 : DFF_X1 port map( D => n3126, CK => CLK, Q => n_2827, QN 
                           => n52311);
   clk_r_REG14869_S1 : DFF_X1 port map( D => n3477, CK => CLK, Q => n_2828, QN 
                           => n52310);
   clk_r_REG15660_S1 : DFF_X1 port map( D => n3028, CK => CLK, Q => n_2829, QN 
                           => n52309);
   clk_r_REG14399_S1 : DFF_X1 port map( D => n3413, CK => CLK, Q => n_2830, QN 
                           => n52308);
   clk_r_REG14937_S1 : DFF_X1 port map( D => n3285, CK => CLK, Q => n_2831, QN 
                           => n52307);
   clk_r_REG15084_S1 : DFF_X1 port map( D => n3058, CK => CLK, Q => n_2832, QN 
                           => n52306);
   clk_r_REG14935_S1 : DFF_X1 port map( D => n3286, CK => CLK, Q => n_2833, QN 
                           => n52305);
   clk_r_REG15281_S1 : DFF_X1 port map( D => n3251, CK => CLK, Q => n_2834, QN 
                           => n52304);
   clk_r_REG15209_S1 : DFF_X1 port map( D => n3191, CK => CLK, Q => n_2835, QN 
                           => n52303);
   clk_r_REG15148_S1 : DFF_X1 port map( D => n3156, CK => CLK, Q => n_2836, QN 
                           => n52302);
   clk_r_REG16484_S1 : DFF_X1 port map( D => n3127, CK => CLK, Q => n_2837, QN 
                           => n52301);
   clk_r_REG16423_S1 : DFF_X1 port map( D => n3093, CK => CLK, Q => n_2838, QN 
                           => n52300);
   clk_r_REG15598_S1 : DFF_X1 port map( D => n2995, CK => CLK, Q => n_2839, QN 
                           => n52299);
   clk_r_REG15082_S1 : DFF_X1 port map( D => n3059, CK => CLK, Q => n_2840, QN 
                           => n52298);
   clk_r_REG15658_S1 : DFF_X1 port map( D => n3029, CK => CLK, Q => n_2841, QN 
                           => n52297);
   clk_r_REG15596_S1 : DFF_X1 port map( D => n2996, CK => CLK, Q => n_2842, QN 
                           => n52296);
   clk_r_REG15530_S1 : DFF_X1 port map( D => n2965, CK => CLK, Q => n_2843, QN 
                           => n52295);
   clk_r_REG15484_S1 : DFF_X1 port map( D => n2935, CK => CLK, Q => n_2844, QN 
                           => n52294);
   clk_r_REG15080_S1 : DFF_X1 port map( D => n3060, CK => CLK, Q => n_2845, QN 
                           => n52293);
   clk_r_REG15594_S1 : DFF_X1 port map( D => n2997, CK => CLK, Q => n_2846, QN 
                           => n52292);
   clk_r_REG16421_S1 : DFF_X1 port map( D => n3094, CK => CLK, Q => n_2847, QN 
                           => n52291);
   clk_r_REG16482_S1 : DFF_X1 port map( D => n3128, CK => CLK, Q => n_2848, QN 
                           => n52290);
   clk_r_REG15207_S1 : DFF_X1 port map( D => n3192, CK => CLK, Q => n_2849, QN 
                           => n52289);
   clk_r_REG15528_S1 : DFF_X1 port map( D => n2966, CK => CLK, Q => n_2850, QN 
                           => n52288);
   clk_r_REG15279_S1 : DFF_X1 port map( D => n3252, CK => CLK, Q => n_2851, QN 
                           => n52287);
   clk_r_REG16235_S1 : DFF_X1 port map( D => n2868, CK => CLK, Q => n_2852, QN 
                           => n52286);
   clk_r_REG16650_S1 : DFF_X1 port map( D => n3540, CK => CLK, Q => n_2853, QN 
                           => n52285);
   clk_r_REG15078_S1 : DFF_X1 port map( D => n3061, CK => CLK, Q => n_2854, QN 
                           => n52284);
   clk_r_REG16419_S1 : DFF_X1 port map( D => n3095, CK => CLK, Q => n_2855, QN 
                           => n52283);
   clk_r_REG16480_S1 : DFF_X1 port map( D => n3129, CK => CLK, Q => n_2856, QN 
                           => n52282);
   clk_r_REG15146_S1 : DFF_X1 port map( D => n3157, CK => CLK, Q => n_2857, QN 
                           => n52281);
   clk_r_REG14933_S1 : DFF_X1 port map( D => n3287, CK => CLK, Q => n_2858, QN 
                           => n52280);
   clk_r_REG15277_S1 : DFF_X1 port map( D => n3253, CK => CLK, Q => n_2859, QN 
                           => n52279);
   clk_r_REG15205_S1 : DFF_X1 port map( D => n3193, CK => CLK, Q => n_2860, QN 
                           => n52278);
   clk_r_REG15275_S1 : DFF_X1 port map( D => n3254, CK => CLK, Q => n_2861, QN 
                           => n52277);
   clk_r_REG14931_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n_2862, QN 
                           => n52276);
   clk_r_REG15203_S1 : DFF_X1 port map( D => n3194, CK => CLK, Q => n_2863, QN 
                           => n52275);
   clk_r_REG15144_S1 : DFF_X1 port map( D => n3158, CK => CLK, Q => n_2864, QN 
                           => n52274);
   clk_r_REG16478_S1 : DFF_X1 port map( D => n3130, CK => CLK, Q => n_2865, QN 
                           => n52273);
   clk_r_REG16417_S1 : DFF_X1 port map( D => n3096, CK => CLK, Q => n_2866, QN 
                           => n52272);
   clk_r_REG15526_S1 : DFF_X1 port map( D => n2967, CK => CLK, Q => n_2867, QN 
                           => n52271);
   clk_r_REG15482_S1 : DFF_X1 port map( D => n2936, CK => CLK, Q => n_2868, QN 
                           => n52270);
   clk_r_REG15410_S1 : DFF_X1 port map( D => n2897, CK => CLK, Q => n_2869, QN 
                           => n52269);
   clk_r_REG16177_S1 : DFF_X1 port map( D => n2833, CK => CLK, Q => n_2870, QN 
                           => n52268);
   clk_r_REG16113_S1 : DFF_X1 port map( D => n2801, CK => CLK, Q => n_2871, QN 
                           => n52267);
   clk_r_REG16233_S1 : DFF_X1 port map( D => n2869, CK => CLK, Q => n_2872, QN 
                           => n52266);
   clk_r_REG16111_S1 : DFF_X1 port map( D => n2802, CK => CLK, Q => n_2873, QN 
                           => n52265);
   clk_r_REG16175_S1 : DFF_X1 port map( D => n2834, CK => CLK, Q => n_2874, QN 
                           => n52264);
   clk_r_REG15408_S1 : DFF_X1 port map( D => n2898, CK => CLK, Q => n_2875, QN 
                           => n52263);
   clk_r_REG15480_S1 : DFF_X1 port map( D => n2937, CK => CLK, Q => n_2876, QN 
                           => n52262);
   clk_r_REG16231_S1 : DFF_X1 port map( D => n2870, CK => CLK, Q => n_2877, QN 
                           => n52261);
   clk_r_REG16229_S1 : DFF_X1 port map( D => n2871, CK => CLK, Q => n_2878, QN 
                           => n52260);
   clk_r_REG16227_S1 : DFF_X1 port map( D => n2872, CK => CLK, Q => n_2879, QN 
                           => n52259);
   clk_r_REG16225_S1 : DFF_X1 port map( D => n2873, CK => CLK, Q => n_2880, QN 
                           => n52258);
   clk_r_REG15524_S1 : DFF_X1 port map( D => n2968, CK => CLK, Q => n_2881, QN 
                           => n52257);
   clk_r_REG15076_S1 : DFF_X1 port map( D => n3062, CK => CLK, Q => n_2882, QN 
                           => n52256);
   clk_r_REG16415_S1 : DFF_X1 port map( D => n3097, CK => CLK, Q => n_2883, QN 
                           => n52255);
   clk_r_REG16476_S1 : DFF_X1 port map( D => n3131, CK => CLK, Q => n_2884, QN 
                           => n52254);
   clk_r_REG15142_S1 : DFF_X1 port map( D => n3159, CK => CLK, Q => n_2885, QN 
                           => n52253);
   clk_r_REG15201_S1 : DFF_X1 port map( D => n3195, CK => CLK, Q => n_2886, QN 
                           => n52252);
   clk_r_REG15592_S1 : DFF_X1 port map( D => n2998, CK => CLK, Q => n_2887, QN 
                           => n52251);
   clk_r_REG14397_S1 : DFF_X1 port map( D => n3414, CK => CLK, Q => n_2888, QN 
                           => n52250);
   clk_r_REG14805_S1 : DFF_X1 port map( D => n3313, CK => CLK, Q => n_2889, QN 
                           => n52249);
   clk_r_REG14727_S1 : DFF_X1 port map( D => n3446, CK => CLK, Q => n_2890, QN 
                           => n52248);
   clk_r_REG14803_S1 : DFF_X1 port map( D => n3314, CK => CLK, Q => n_2891, QN 
                           => n52247);
   clk_r_REG14651_S1 : DFF_X1 port map( D => n3382, CK => CLK, Q => n_2892, QN 
                           => n52246);
   clk_r_REG14801_S1 : DFF_X1 port map( D => n3315, CK => CLK, Q => n_2893, QN 
                           => n52245);
   clk_r_REG15009_S1 : DFF_X1 port map( D => n3510, CK => CLK, Q => n_2894, QN 
                           => n52244);
   clk_r_REG15074_S1 : DFF_X1 port map( D => n3063, CK => CLK, Q => n_2895, QN 
                           => n52243);
   clk_r_REG14725_S1 : DFF_X1 port map( D => n3447, CK => CLK, Q => n_2896, QN 
                           => n52242);
   clk_r_REG15072_S1 : DFF_X1 port map( D => n3064, CK => CLK, Q => n_2897, QN 
                           => n52241);
   clk_r_REG15590_S1 : DFF_X1 port map( D => n2999, CK => CLK, Q => n_2898, QN 
                           => n52240);
   clk_r_REG14395_S1 : DFF_X1 port map( D => n3415, CK => CLK, Q => n_2899, QN 
                           => n52239);
   clk_r_REG15007_S1 : DFF_X1 port map( D => n3511, CK => CLK, Q => n_2900, QN 
                           => n52238);
   clk_r_REG14393_S1 : DFF_X1 port map( D => n3416, CK => CLK, Q => n_2901, QN 
                           => n52237);
   clk_r_REG15338_S1 : DFF_X1 port map( D => n3350, CK => CLK, Q => n_2902, QN 
                           => n52236);
   clk_r_REG15336_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n_2903, QN 
                           => n52235);
   clk_r_REG15005_S1 : DFF_X1 port map( D => n3512, CK => CLK, Q => n_2904, QN 
                           => n52234);
   clk_r_REG14649_S1 : DFF_X1 port map( D => n3383, CK => CLK, Q => n_2905, QN 
                           => n52233);
   clk_r_REG15334_S1 : DFF_X1 port map( D => n3352, CK => CLK, Q => n_2906, QN 
                           => n52232);
   clk_r_REG14723_S1 : DFF_X1 port map( D => n3448, CK => CLK, Q => n_2907, QN 
                           => n52231);
   clk_r_REG14647_S1 : DFF_X1 port map( D => n3384, CK => CLK, Q => n_2908, QN 
                           => n52230);
   clk_r_REG16648_S1 : DFF_X1 port map( D => n3541, CK => CLK, Q => n_2909, QN 
                           => n52229);
   clk_r_REG14867_S1 : DFF_X1 port map( D => n3478, CK => CLK, Q => n_2910, QN 
                           => n52228);
   clk_r_REG16646_S1 : DFF_X1 port map( D => n3542, CK => CLK, Q => n_2911, QN 
                           => n52227);
   clk_r_REG16644_S1 : DFF_X1 port map( D => n3543, CK => CLK, Q => n_2912, QN 
                           => n52226);
   clk_r_REG15588_S1 : DFF_X1 port map( D => n3000, CK => CLK, Q => n_2913, QN 
                           => n52225);
   clk_r_REG15586_S1 : DFF_X1 port map( D => n3001, CK => CLK, Q => n_2914, QN 
                           => n52224);
   clk_r_REG15273_S1 : DFF_X1 port map( D => n3255, CK => CLK, Q => n_2915, QN 
                           => n52223);
   clk_r_REG14929_S1 : DFF_X1 port map( D => n3289, CK => CLK, Q => n_2916, QN 
                           => n52222);
   clk_r_REG15584_S1 : DFF_X1 port map( D => n3002, CK => CLK, Q => n_2917, QN 
                           => n52221);
   clk_r_REG14721_S1 : DFF_X1 port map( D => n3449, CK => CLK, Q => n_2918, QN 
                           => n52220);
   clk_r_REG14799_S1 : DFF_X1 port map( D => n3316, CK => CLK, Q => n_2919, QN 
                           => n52219);
   clk_r_REG14865_S1 : DFF_X1 port map( D => n3479, CK => CLK, Q => n_2920, QN 
                           => n52218);
   clk_r_REG15070_S1 : DFF_X1 port map( D => n3065, CK => CLK, Q => n_2921, QN 
                           => n52217);
   clk_r_REG14645_S1 : DFF_X1 port map( D => n3385, CK => CLK, Q => n_2922, QN 
                           => n52216);
   clk_r_REG15332_S1 : DFF_X1 port map( D => n3353, CK => CLK, Q => n_2923, QN 
                           => n52215);
   clk_r_REG15406_S1 : DFF_X1 port map( D => n2899, CK => CLK, Q => n_2924, QN 
                           => n52214);
   clk_r_REG15582_S1 : DFF_X1 port map( D => n3003, CK => CLK, Q => n_2925, QN 
                           => n52213);
   clk_r_REG14391_S1 : DFF_X1 port map( D => n3417, CK => CLK, Q => n_2926, QN 
                           => n52212);
   clk_r_REG15003_S1 : DFF_X1 port map( D => n3513, CK => CLK, Q => n_2927, QN 
                           => n52211);
   clk_r_REG14863_S1 : DFF_X1 port map( D => n3480, CK => CLK, Q => n_2928, QN 
                           => n52210);
   clk_r_REG15580_S1 : DFF_X1 port map( D => n3004, CK => CLK, Q => n_2929, QN 
                           => n52209);
   clk_r_REG14797_S1 : DFF_X1 port map( D => n3317, CK => CLK, Q => n_2930, QN 
                           => n52208);
   clk_r_REG14643_S1 : DFF_X1 port map( D => n3386, CK => CLK, Q => n_2931, QN 
                           => n52207);
   clk_r_REG15404_S1 : DFF_X1 port map( D => n2900, CK => CLK, Q => n_2932, QN 
                           => n52206);
   clk_r_REG14719_S1 : DFF_X1 port map( D => n3450, CK => CLK, Q => n_2933, QN 
                           => n52205);
   clk_r_REG15330_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n_2934, QN 
                           => n52204);
   clk_r_REG15001_S1 : DFF_X1 port map( D => n3514, CK => CLK, Q => n_2935, QN 
                           => n52203);
   clk_r_REG14389_S1 : DFF_X1 port map( D => n3418, CK => CLK, Q => n_2936, QN 
                           => n52202);
   clk_r_REG15068_S1 : DFF_X1 port map( D => n3066, CK => CLK, Q => n_2937, QN 
                           => n52201);
   clk_r_REG15578_S1 : DFF_X1 port map( D => n3005, CK => CLK, Q => n_2938, QN 
                           => n52200);
   clk_r_REG14861_S1 : DFF_X1 port map( D => n3481, CK => CLK, Q => n_2939, QN 
                           => n52199);
   clk_r_REG14859_S1 : DFF_X1 port map( D => n3482, CK => CLK, Q => n_2940, QN 
                           => n52198);
   clk_r_REG15656_S1 : DFF_X1 port map( D => n3030, CK => CLK, Q => n_2941, QN 
                           => n52197);
   clk_r_REG15522_S1 : DFF_X1 port map( D => n2969, CK => CLK, Q => n_2942, QN 
                           => n52196);
   clk_r_REG15654_S1 : DFF_X1 port map( D => n3031, CK => CLK, Q => n_2943, QN 
                           => n52195);
   clk_r_REG14927_S1 : DFF_X1 port map( D => n3290, CK => CLK, Q => n_2944, QN 
                           => n52194);
   clk_r_REG15271_S1 : DFF_X1 port map( D => n3256, CK => CLK, Q => n_2945, QN 
                           => n52193);
   clk_r_REG16413_S1 : DFF_X1 port map( D => n3098, CK => CLK, Q => n_2946, QN 
                           => n52192);
   clk_r_REG14925_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n_2947, QN 
                           => n52191);
   clk_r_REG16411_S1 : DFF_X1 port map( D => n3099, CK => CLK, Q => n_2948, QN 
                           => n52190);
   clk_r_REG15140_S1 : DFF_X1 port map( D => n3160, CK => CLK, Q => n_2949, QN 
                           => n52189);
   clk_r_REG15138_S1 : DFF_X1 port map( D => n3161, CK => CLK, Q => n_2950, QN 
                           => n52188);
   clk_r_REG14795_S1 : DFF_X1 port map( D => n3318, CK => CLK, Q => n_2951, QN 
                           => n52187);
   clk_r_REG14793_S1 : DFF_X1 port map( D => n3319, CK => CLK, Q => n_2952, QN 
                           => n52186);
   clk_r_REG15652_S1 : DFF_X1 port map( D => n3032, CK => CLK, Q => n_2953, QN 
                           => n52185);
   clk_r_REG14791_S1 : DFF_X1 port map( D => n3320, CK => CLK, Q => n_2954, QN 
                           => n52184);
   clk_r_REG14789_S1 : DFF_X1 port map( D => n3321, CK => CLK, Q => n_2955, QN 
                           => n52183);
   clk_r_REG16109_S1 : DFF_X1 port map( D => n2803, CK => CLK, Q => n_2956, QN 
                           => n52182);
   clk_r_REG16173_S1 : DFF_X1 port map( D => n2835, CK => CLK, Q => n_2957, QN 
                           => n52181);
   clk_r_REG16107_S1 : DFF_X1 port map( D => n2804, CK => CLK, Q => n_2958, QN 
                           => n52180);
   clk_r_REG16171_S1 : DFF_X1 port map( D => n2836, CK => CLK, Q => n_2959, QN 
                           => n52179);
   clk_r_REG16105_S1 : DFF_X1 port map( D => n2805, CK => CLK, Q => n_2960, QN 
                           => n52178);
   clk_r_REG16169_S1 : DFF_X1 port map( D => n2837, CK => CLK, Q => n_2961, QN 
                           => n52177);
   clk_r_REG16103_S1 : DFF_X1 port map( D => n2806, CK => CLK, Q => n_2962, QN 
                           => n52176);
   clk_r_REG16167_S1 : DFF_X1 port map( D => n2838, CK => CLK, Q => n_2963, QN 
                           => n52175);
   clk_r_REG16165_S1 : DFF_X1 port map( D => n2839, CK => CLK, Q => n_2964, QN 
                           => n52174);
   clk_r_REG15402_S1 : DFF_X1 port map( D => n2901, CK => CLK, Q => n_2965, QN 
                           => n52173);
   clk_r_REG16163_S1 : DFF_X1 port map( D => n2840, CK => CLK, Q => n_2966, QN 
                           => n52172);
   clk_r_REG16161_S1 : DFF_X1 port map( D => n2841, CK => CLK, Q => n_2967, QN 
                           => n52171);
   clk_r_REG15650_S1 : DFF_X1 port map( D => n3033, CK => CLK, Q => n_2968, QN 
                           => n52170);
   clk_r_REG15648_S1 : DFF_X1 port map( D => n3034, CK => CLK, Q => n_2969, QN 
                           => n52169);
   clk_r_REG15400_S1 : DFF_X1 port map( D => n2902, CK => CLK, Q => n_2970, QN 
                           => n52168);
   clk_r_REG16642_S1 : DFF_X1 port map( D => n3544, CK => CLK, Q => n_2971, QN 
                           => n52167);
   clk_r_REG16640_S1 : DFF_X1 port map( D => n3545, CK => CLK, Q => n_2972, QN 
                           => n52166);
   clk_r_REG16638_S1 : DFF_X1 port map( D => n3546, CK => CLK, Q => n_2973, QN 
                           => n52165);
   clk_r_REG15398_S1 : DFF_X1 port map( D => n2903, CK => CLK, Q => n_2974, QN 
                           => n52164);
   clk_r_REG16556_S1 : DFF_X1 port map( D => n3219, CK => CLK, Q => n_2975, QN 
                           => n52163);
   clk_r_REG16554_S1 : DFF_X1 port map( D => n3220, CK => CLK, Q => n_2976, QN 
                           => n52162);
   clk_r_REG16101_S1 : DFF_X1 port map( D => n2807, CK => CLK, Q => n_2977, QN 
                           => n52161);
   clk_r_REG16552_S1 : DFF_X1 port map( D => n3221, CK => CLK, Q => n_2978, QN 
                           => n52160);
   clk_r_REG15136_S1 : DFF_X1 port map( D => n3162, CK => CLK, Q => n_2979, QN 
                           => n52159);
   clk_r_REG16636_S1 : DFF_X1 port map( D => n3547, CK => CLK, Q => n_2980, QN 
                           => n52158);
   clk_r_REG15199_S1 : DFF_X1 port map( D => n3196, CK => CLK, Q => n_2981, QN 
                           => n52157);
   clk_r_REG14787_S1 : DFF_X1 port map( D => n3322, CK => CLK, Q => n_2982, QN 
                           => n52156);
   clk_r_REG16159_S1 : DFF_X1 port map( D => n2842, CK => CLK, Q => n_2983, QN 
                           => n52155);
   clk_r_REG15646_S1 : DFF_X1 port map( D => n3035, CK => CLK, Q => n_2984, QN 
                           => n52154);
   clk_r_REG16474_S1 : DFF_X1 port map( D => n3132, CK => CLK, Q => n_2985, QN 
                           => n52153);
   clk_r_REG15396_S1 : DFF_X1 port map( D => n2904, CK => CLK, Q => n_2986, QN 
                           => n52152);
   clk_r_REG15520_S1 : DFF_X1 port map( D => n2970, CK => CLK, Q => n_2987, QN 
                           => n52151);
   clk_r_REG14923_S1 : DFF_X1 port map( D => n3292, CK => CLK, Q => n_2988, QN 
                           => n52150);
   clk_r_REG16099_S1 : DFF_X1 port map( D => n2808, CK => CLK, Q => n_2989, QN 
                           => n52149);
   clk_r_REG15269_S1 : DFF_X1 port map( D => n3257, CK => CLK, Q => n_2990, QN 
                           => n52148);
   clk_r_REG16409_S1 : DFF_X1 port map( D => n3100, CK => CLK, Q => n_2991, QN 
                           => n52147);
   clk_r_REG16407_S1 : DFF_X1 port map( D => n3101, CK => CLK, Q => n_2992, QN 
                           => n52146);
   clk_r_REG15394_S1 : DFF_X1 port map( D => n2905, CK => CLK, Q => n_2993, QN 
                           => n52145);
   clk_r_REG16405_S1 : DFF_X1 port map( D => n3102, CK => CLK, Q => n_2994, QN 
                           => n52144);
   clk_r_REG15392_S1 : DFF_X1 port map( D => n2906, CK => CLK, Q => n_2995, QN 
                           => n52143);
   clk_r_REG16097_S1 : DFF_X1 port map( D => n2809, CK => CLK, Q => n_2996, QN 
                           => n52142);
   clk_r_REG16095_S1 : DFF_X1 port map( D => n2810, CK => CLK, Q => n_2997, QN 
                           => n52141);
   clk_r_REG16093_S1 : DFF_X1 port map( D => n2811, CK => CLK, Q => n_2998, QN 
                           => n52140);
   clk_r_REG16157_S1 : DFF_X1 port map( D => n2843, CK => CLK, Q => n_2999, QN 
                           => n52139);
   clk_r_REG16091_S1 : DFF_X1 port map( D => n2812, CK => CLK, Q => n_3000, QN 
                           => n52138);
   clk_r_REG16155_S1 : DFF_X1 port map( D => n2844, CK => CLK, Q => n_3001, QN 
                           => n52137);
   clk_r_REG16153_S1 : DFF_X1 port map( D => n2845, CK => CLK, Q => n_3002, QN 
                           => n52136);
   clk_r_REG15518_S1 : DFF_X1 port map( D => n2971, CK => CLK, Q => n_3003, QN 
                           => n52135);
   clk_r_REG14921_S1 : DFF_X1 port map( D => n3293, CK => CLK, Q => n_3004, QN 
                           => n52134);
   clk_r_REG15644_S1 : DFF_X1 port map( D => n3036, CK => CLK, Q => n_3005, QN 
                           => n52133);
   clk_r_REG14919_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n_3006, QN 
                           => n52132);
   clk_r_REG16403_S1 : DFF_X1 port map( D => n3103, CK => CLK, Q => n_3007, QN 
                           => n52131);
   clk_r_REG14917_S1 : DFF_X1 port map( D => n3295, CK => CLK, Q => n_3008, QN 
                           => n52130);
   clk_r_REG15516_S1 : DFF_X1 port map( D => n2972, CK => CLK, Q => n_3009, QN 
                           => n52129);
   clk_r_REG15390_S1 : DFF_X1 port map( D => n2907, CK => CLK, Q => n_3010, QN 
                           => n52128);
   clk_r_REG16151_S1 : DFF_X1 port map( D => n2846, CK => CLK, Q => n_3011, QN 
                           => n52127);
   clk_r_REG15267_S1 : DFF_X1 port map( D => n3258, CK => CLK, Q => n_3012, QN 
                           => n52126);
   clk_r_REG15066_S1 : DFF_X1 port map( D => n3067, CK => CLK, Q => n_3013, QN 
                           => n52125);
   clk_r_REG16149_S1 : DFF_X1 port map( D => n2847, CK => CLK, Q => n_3014, QN 
                           => n52124);
   clk_r_REG14785_S1 : DFF_X1 port map( D => n3323, CK => CLK, Q => n_3015, QN 
                           => n52123);
   clk_r_REG15328_S1 : DFF_X1 port map( D => n3355, CK => CLK, Q => n_3016, QN 
                           => n52122);
   clk_r_REG15064_S1 : DFF_X1 port map( D => n3068, CK => CLK, Q => n_3017, QN 
                           => n52121);
   clk_r_REG16634_S1 : DFF_X1 port map( D => n3548, CK => CLK, Q => n_3018, QN 
                           => n52120);
   clk_r_REG14387_S1 : DFF_X1 port map( D => n3419, CK => CLK, Q => n_3019, QN 
                           => n52119);
   clk_r_REG14999_S1 : DFF_X1 port map( D => n3515, CK => CLK, Q => n_3020, QN 
                           => n52118);
   clk_r_REG14783_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n_3021, QN 
                           => n52117);
   clk_r_REG14857_S1 : DFF_X1 port map( D => n3483, CK => CLK, Q => n_3022, QN 
                           => n52116);
   clk_r_REG14997_S1 : DFF_X1 port map( D => n3516, CK => CLK, Q => n_3023, QN 
                           => n52115);
   clk_r_REG14385_S1 : DFF_X1 port map( D => n3420, CK => CLK, Q => n_3024, QN 
                           => n52114);
   clk_r_REG14995_S1 : DFF_X1 port map( D => n3517, CK => CLK, Q => n_3025, QN 
                           => n52113);
   clk_r_REG16550_S1 : DFF_X1 port map( D => n3222, CK => CLK, Q => n_3026, QN 
                           => n52112);
   clk_r_REG15062_S1 : DFF_X1 port map( D => n3069, CK => CLK, Q => n_3027, QN 
                           => n52111);
   clk_r_REG14641_S1 : DFF_X1 port map( D => n3387, CK => CLK, Q => n_3028, QN 
                           => n52110);
   clk_r_REG15197_S1 : DFF_X1 port map( D => n3197, CK => CLK, Q => n_3029, QN 
                           => n52109);
   clk_r_REG14717_S1 : DFF_X1 port map( D => n3451, CK => CLK, Q => n_3030, QN 
                           => n52108);
   clk_r_REG14715_S1 : DFF_X1 port map( D => n3452, CK => CLK, Q => n_3031, QN 
                           => n52107);
   clk_r_REG14713_S1 : DFF_X1 port map( D => n3453, CK => CLK, Q => n_3032, QN 
                           => n52106);
   clk_r_REG14639_S1 : DFF_X1 port map( D => n3388, CK => CLK, Q => n_3033, QN 
                           => n52105);
   clk_r_REG15388_S1 : DFF_X1 port map( D => n2908, CK => CLK, Q => n_3034, QN 
                           => n52104);
   clk_r_REG14855_S1 : DFF_X1 port map( D => n3484, CK => CLK, Q => n_3035, QN 
                           => n52103);
   clk_r_REG14383_S1 : DFF_X1 port map( D => n3421, CK => CLK, Q => n_3036, QN 
                           => n52102);
   clk_r_REG16632_S1 : DFF_X1 port map( D => n3549, CK => CLK, Q => n_3037, QN 
                           => n52101);
   clk_r_REG14711_S1 : DFF_X1 port map( D => n3454, CK => CLK, Q => n_3038, QN 
                           => n52100);
   clk_r_REG14853_S1 : DFF_X1 port map( D => n3485, CK => CLK, Q => n_3039, QN 
                           => n52099);
   clk_r_REG15195_S1 : DFF_X1 port map( D => n3198, CK => CLK, Q => n_3040, QN 
                           => n52098);
   clk_r_REG16630_S1 : DFF_X1 port map( D => n3550, CK => CLK, Q => n_3041, QN 
                           => n52097);
   clk_r_REG14993_S1 : DFF_X1 port map( D => n3518, CK => CLK, Q => n_3042, QN 
                           => n52096);
   clk_r_REG15193_S1 : DFF_X1 port map( D => n3199, CK => CLK, Q => n_3043, QN 
                           => n52095);
   clk_r_REG14991_S1 : DFF_X1 port map( D => n3519, CK => CLK, Q => n_3044, QN 
                           => n52094);
   clk_r_REG14637_S1 : DFF_X1 port map( D => n3389, CK => CLK, Q => n_3045, QN 
                           => n52093);
   clk_r_REG15134_S1 : DFF_X1 port map( D => n3163, CK => CLK, Q => n_3046, QN 
                           => n52092);
   clk_r_REG14781_S1 : DFF_X1 port map( D => n3325, CK => CLK, Q => n_3047, QN 
                           => n52091);
   clk_r_REG15132_S1 : DFF_X1 port map( D => n3164, CK => CLK, Q => n_3048, QN 
                           => n52090);
   clk_r_REG14635_S1 : DFF_X1 port map( D => n3390, CK => CLK, Q => n_3049, QN 
                           => n52089);
   clk_r_REG16472_S1 : DFF_X1 port map( D => n3133, CK => CLK, Q => n_3050, QN 
                           => n52088);
   clk_r_REG15326_S1 : DFF_X1 port map( D => n3356, CK => CLK, Q => n_3051, QN 
                           => n52087);
   clk_r_REG14633_S1 : DFF_X1 port map( D => n3391, CK => CLK, Q => n_3052, QN 
                           => n52086);
   clk_r_REG15130_S1 : DFF_X1 port map( D => n3165, CK => CLK, Q => n_3053, QN 
                           => n52085);
   clk_r_REG15324_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n_3054, QN 
                           => n52084);
   clk_r_REG14779_S1 : DFF_X1 port map( D => n3326, CK => CLK, Q => n_3055, QN 
                           => n52083);
   clk_r_REG14851_S1 : DFF_X1 port map( D => n3486, CK => CLK, Q => n_3056, QN 
                           => n52082);
   clk_r_REG14381_S1 : DFF_X1 port map( D => n3422, CK => CLK, Q => n_3057, QN 
                           => n52081);
   clk_r_REG16470_S1 : DFF_X1 port map( D => n3134, CK => CLK, Q => n_3058, QN 
                           => n52080);
   clk_r_REG14709_S1 : DFF_X1 port map( D => n3455, CK => CLK, Q => n_3059, QN 
                           => n52079);
   clk_r_REG15322_S1 : DFF_X1 port map( D => n3358, CK => CLK, Q => n_3060, QN 
                           => n52078);
   clk_r_REG14379_S1 : DFF_X1 port map( D => n3423, CK => CLK, Q => n_3061, QN 
                           => n52077);
   clk_r_REG16468_S1 : DFF_X1 port map( D => n3135, CK => CLK, Q => n_3062, QN 
                           => n52076);
   clk_r_REG14849_S1 : DFF_X1 port map( D => n3487, CK => CLK, Q => n_3063, QN 
                           => n52075);
   clk_r_REG15320_S1 : DFF_X1 port map( D => n3359, CK => CLK, Q => n_3064, QN 
                           => n52074);
   clk_r_REG15642_S1 : DFF_X1 port map( D => n3037, CK => CLK, Q => n_3065, QN 
                           => n52073);
   clk_r_REG15640_S1 : DFF_X1 port map( D => n3038, CK => CLK, Q => n_3066, QN 
                           => n52072);
   clk_r_REG15638_S1 : DFF_X1 port map( D => n3039, CK => CLK, Q => n_3067, QN 
                           => n52071);
   clk_r_REG15688_S1 : DFF_X1 port map( D => n3014, CK => CLK, Q => n_3068, QN 
                           => n52070);
   clk_r_REG15686_S1 : DFF_X1 port map( D => n3015, CK => CLK, Q => n_3069, QN 
                           => n52069);
   clk_r_REG15243_S1 : DFF_X1 port map( D => n3174, CK => CLK, Q => n_3070, QN 
                           => n52068);
   clk_r_REG15478_S1 : DFF_X1 port map( D => n2938, CK => CLK, Q => n_3071, QN 
                           => n52067);
   clk_r_REG15241_S1 : DFF_X1 port map( D => n3175, CK => CLK, Q => n_3072, QN 
                           => n52066);
   clk_r_REG15191_S1 : DFF_X1 port map( D => n3200, CK => CLK, Q => n_3073, QN 
                           => n52065);
   clk_r_REG15239_S1 : DFF_X1 port map( D => n3176, CK => CLK, Q => n_3074, QN 
                           => n52064);
   clk_r_REG15189_S1 : DFF_X1 port map( D => n3201, CK => CLK, Q => n_3075, QN 
                           => n52063);
   clk_r_REG15187_S1 : DFF_X1 port map( D => n3202, CK => CLK, Q => n_3076, QN 
                           => n52062);
   clk_r_REG15576_S1 : DFF_X1 port map( D => n3006, CK => CLK, Q => n_3077, QN 
                           => n52061);
   clk_r_REG15128_S1 : DFF_X1 port map( D => n3166, CK => CLK, Q => n_3078, QN 
                           => n52060);
   clk_r_REG15126_S1 : DFF_X1 port map( D => n3167, CK => CLK, Q => n_3079, QN 
                           => n52059);
   clk_r_REG15176_S1 : DFF_X1 port map( D => n3142, CK => CLK, Q => n_3080, QN 
                           => n52058);
   clk_r_REG15174_S1 : DFF_X1 port map( D => n3143, CK => CLK, Q => n_3081, QN 
                           => n52057);
   clk_r_REG15514_S1 : DFF_X1 port map( D => n2973, CK => CLK, Q => n_3082, QN 
                           => n52056);
   clk_r_REG15124_S1 : DFF_X1 port map( D => n3168, CK => CLK, Q => n_3083, QN 
                           => n52055);
   clk_r_REG16518_S1 : DFF_X1 port map( D => n3110, CK => CLK, Q => n_3084, QN 
                           => n52054);
   clk_r_REG16516_S1 : DFF_X1 port map( D => n3111, CK => CLK, Q => n_3085, QN 
                           => n52053);
   clk_r_REG16466_S1 : DFF_X1 port map( D => n3136, CK => CLK, Q => n_3086, QN 
                           => n52052);
   clk_r_REG16514_S1 : DFF_X1 port map( D => n3112, CK => CLK, Q => n_3087, QN 
                           => n52051);
   clk_r_REG16464_S1 : DFF_X1 port map( D => n3137, CK => CLK, Q => n_3088, QN 
                           => n52050);
   clk_r_REG16453_S1 : DFF_X1 port map( D => n3078, CK => CLK, Q => n_3089, QN 
                           => n52049);
   clk_r_REG16451_S1 : DFF_X1 port map( D => n3079, CK => CLK, Q => n_3090, QN 
                           => n52048);
   clk_r_REG15060_S1 : DFF_X1 port map( D => n3070, CK => CLK, Q => n_3091, QN 
                           => n52047);
   clk_r_REG16401_S1 : DFF_X1 port map( D => n3104, CK => CLK, Q => n_3092, QN 
                           => n52046);
   clk_r_REG16449_S1 : DFF_X1 port map( D => n3080, CK => CLK, Q => n_3093, QN 
                           => n52045);
   clk_r_REG14967_S1 : DFF_X1 port map( D => n3270, CK => CLK, Q => n_3094, QN 
                           => n52044);
   clk_r_REG14965_S1 : DFF_X1 port map( D => n3271, CK => CLK, Q => n_3095, QN 
                           => n52043);
   clk_r_REG14915_S1 : DFF_X1 port map( D => n3296, CK => CLK, Q => n_3096, QN 
                           => n52042);
   clk_r_REG14963_S1 : DFF_X1 port map( D => n3272, CK => CLK, Q => n_3097, QN 
                           => n52041);
   clk_r_REG14913_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n_3098, QN 
                           => n52040);
   clk_r_REG14911_S1 : DFF_X1 port map( D => n3298, CK => CLK, Q => n_3099, QN 
                           => n52039);
   clk_r_REG15265_S1 : DFF_X1 port map( D => n3259, CK => CLK, Q => n_3100, QN 
                           => n52038);
   clk_r_REG15263_S1 : DFF_X1 port map( D => n3260, CK => CLK, Q => n_3101, QN 
                           => n52037);
   clk_r_REG15261_S1 : DFF_X1 port map( D => n3261, CK => CLK, Q => n_3102, QN 
                           => n52036);
   clk_r_REG15259_S1 : DFF_X1 port map( D => n3262, CK => CLK, Q => n_3103, QN 
                           => n52035);
   clk_r_REG15257_S1 : DFF_X1 port map( D => n3263, CK => CLK, Q => n_3104, QN 
                           => n52034);
   clk_r_REG15307_S1 : DFF_X1 port map( D => n3238, CK => CLK, Q => n_3105, QN 
                           => n52033);
   clk_r_REG14909_S1 : DFF_X1 port map( D => n3299, CK => CLK, Q => n_3106, QN 
                           => n52032);
   clk_r_REG15305_S1 : DFF_X1 port map( D => n3239, CK => CLK, Q => n_3107, QN 
                           => n52031);
   clk_r_REG15185_S1 : DFF_X1 port map( D => n3203, CK => CLK, Q => n_3108, QN 
                           => n52030);
   clk_r_REG16462_S1 : DFF_X1 port map( D => n3138, CK => CLK, Q => n_3109, QN 
                           => n52029);
   clk_r_REG16223_S1 : DFF_X1 port map( D => n2874, CK => CLK, Q => n_3110, QN 
                           => n52028);
   clk_r_REG15476_S1 : DFF_X1 port map( D => n2939, CK => CLK, Q => n_3111, QN 
                           => n52027);
   clk_r_REG15512_S1 : DFF_X1 port map( D => n2974, CK => CLK, Q => n_3112, QN 
                           => n52026);
   clk_r_REG15636_S1 : DFF_X1 port map( D => n3040, CK => CLK, Q => n_3113, QN 
                           => n52025);
   clk_r_REG15574_S1 : DFF_X1 port map( D => n3007, CK => CLK, Q => n_3114, QN 
                           => n52024);
   clk_r_REG15684_S1 : DFF_X1 port map( D => n3016, CK => CLK, Q => n_3115, QN 
                           => n52023);
   clk_r_REG15058_S1 : DFF_X1 port map( D => n3071, CK => CLK, Q => n_3116, QN 
                           => n52022);
   clk_r_REG16399_S1 : DFF_X1 port map( D => n3105, CK => CLK, Q => n_3117, QN 
                           => n52021);
   clk_r_REG16460_S1 : DFF_X1 port map( D => n3139, CK => CLK, Q => n_3118, QN 
                           => n52020);
   clk_r_REG15183_S1 : DFF_X1 port map( D => n3204, CK => CLK, Q => n_3119, QN 
                           => n52019);
   clk_r_REG15255_S1 : DFF_X1 port map( D => n3264, CK => CLK, Q => n_3120, QN 
                           => n52018);
   clk_r_REG14907_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n_3121, QN 
                           => n52017);
   clk_r_REG16221_S1 : DFF_X1 port map( D => n2875, CK => CLK, Q => n_3122, QN 
                           => n52016);
   clk_r_REG15474_S1 : DFF_X1 port map( D => n2940, CK => CLK, Q => n_3123, QN 
                           => n52015);
   clk_r_REG15510_S1 : DFF_X1 port map( D => n2975, CK => CLK, Q => n_3124, QN 
                           => n52014);
   clk_r_REG15624_S1 : DFF_X1 port map( D => n2982, CK => CLK, Q => n_3125, QN 
                           => n52013);
   clk_r_REG15108_S1 : DFF_X1 port map( D => n3046, CK => CLK, Q => n_3126, QN 
                           => n52012);
   clk_r_REG16089_S1 : DFF_X1 port map( D => n2813, CK => CLK, Q => n_3127, QN 
                           => n52011);
   clk_r_REG16199_S1 : DFF_X1 port map( D => n2822, CK => CLK, Q => n_3128, QN 
                           => n52010);
   clk_r_REG15386_S1 : DFF_X1 port map( D => n2909, CK => CLK, Q => n_3129, QN 
                           => n52009);
   clk_r_REG14777_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n_3130, QN 
                           => n52008);
   clk_r_REG16197_S1 : DFF_X1 port map( D => n2823, CK => CLK, Q => n_3131, QN 
                           => n52007);
   clk_r_REG15384_S1 : DFF_X1 port map( D => n2910, CK => CLK, Q => n_3132, QN 
                           => n52006);
   clk_r_REG15382_S1 : DFF_X1 port map( D => n2911, CK => CLK, Q => n_3133, QN 
                           => n52005);
   clk_r_REG14827_S1 : DFF_X1 port map( D => n3302, CK => CLK, Q => n_3134, QN 
                           => n52004);
   clk_r_REG14825_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n_3135, QN 
                           => n52003);
   clk_r_REG16147_S1 : DFF_X1 port map( D => n2848, CK => CLK, Q => n_3136, QN 
                           => n52002);
   clk_r_REG15432_S1 : DFF_X1 port map( D => n2886, CK => CLK, Q => n_3137, QN 
                           => n52001);
   clk_r_REG15430_S1 : DFF_X1 port map( D => n2887, CK => CLK, Q => n_3138, QN 
                           => n52000);
   clk_r_REG15380_S1 : DFF_X1 port map( D => n2912, CK => CLK, Q => n_3139, QN 
                           => n51999);
   clk_r_REG16548_S1 : DFF_X1 port map( D => n3223, CK => CLK, Q => n_3140, QN 
                           => n51998);
   clk_r_REG16546_S1 : DFF_X1 port map( D => n3224, CK => CLK, Q => n_3141, QN 
                           => n51997);
   clk_r_REG14775_S1 : DFF_X1 port map( D => n3328, CK => CLK, Q => n_3142, QN 
                           => n51996);
   clk_r_REG15370_S1 : DFF_X1 port map( D => n3334, CK => CLK, Q => n_3143, QN 
                           => n51995);
   clk_r_REG14823_S1 : DFF_X1 port map( D => n3304, CK => CLK, Q => n_3144, QN 
                           => n51994);
   clk_r_REG14683_S1 : DFF_X1 port map( D => n3366, CK => CLK, Q => n_3145, QN 
                           => n51993);
   clk_r_REG14429_S1 : DFF_X1 port map( D => n3398, CK => CLK, Q => n_3146, QN 
                           => n51992);
   clk_r_REG14759_S1 : DFF_X1 port map( D => n3430, CK => CLK, Q => n_3147, QN 
                           => n51991);
   clk_r_REG14899_S1 : DFF_X1 port map( D => n3462, CK => CLK, Q => n_3148, QN 
                           => n51990);
   clk_r_REG15041_S1 : DFF_X1 port map( D => n3494, CK => CLK, Q => n_3149, QN 
                           => n51989);
   clk_r_REG14897_S1 : DFF_X1 port map( D => n3463, CK => CLK, Q => n_3150, QN 
                           => n51988);
   clk_r_REG14757_S1 : DFF_X1 port map( D => n3431, CK => CLK, Q => n_3151, QN 
                           => n51987);
   clk_r_REG14427_S1 : DFF_X1 port map( D => n3399, CK => CLK, Q => n_3152, QN 
                           => n51986);
   clk_r_REG14681_S1 : DFF_X1 port map( D => n3367, CK => CLK, Q => n_3153, QN 
                           => n51985);
   clk_r_REG15039_S1 : DFF_X1 port map( D => n3495, CK => CLK, Q => n_3154, QN 
                           => n51984);
   clk_r_REG14773_S1 : DFF_X1 port map( D => n3329, CK => CLK, Q => n_3155, QN 
                           => n51983);
   clk_r_REG15368_S1 : DFF_X1 port map( D => n3335, CK => CLK, Q => n_3156, QN 
                           => n51982);
   clk_r_REG16544_S1 : DFF_X1 port map( D => n3225, CK => CLK, Q => n_3157, QN 
                           => n51981);
   clk_r_REG16628_S1 : DFF_X1 port map( D => n3551, CK => CLK, Q => n_3158, QN 
                           => n51980);
   clk_r_REG16678_S1 : DFF_X1 port map( D => n3526, CK => CLK, Q => n_3159, QN 
                           => n51979);
   clk_r_REG16542_S1 : DFF_X1 port map( D => n3226, CK => CLK, Q => n_3160, QN 
                           => n51978);
   clk_r_REG16676_S1 : DFF_X1 port map( D => n3527, CK => CLK, Q => n_3161, QN 
                           => n51977);
   clk_r_REG16540_S1 : DFF_X1 port map( D => n3227, CK => CLK, Q => n_3162, QN 
                           => n51976);
   clk_r_REG16626_S1 : DFF_X1 port map( D => n3552, CK => CLK, Q => n_3163, QN 
                           => n51975);
   clk_r_REG16538_S1 : DFF_X1 port map( D => n3228, CK => CLK, Q => n_3164, QN 
                           => n51974);
   clk_r_REG16674_S1 : DFF_X1 port map( D => n3528, CK => CLK, Q => n_3165, QN 
                           => n51973);
   clk_r_REG16536_S1 : DFF_X1 port map( D => n3229, CK => CLK, Q => n_3166, QN 
                           => n51972);
   clk_r_REG15622_S1 : DFF_X1 port map( D => n2983, CK => CLK, Q => n_3167, QN 
                           => n51971);
   clk_r_REG15572_S1 : DFF_X1 port map( D => n3008, CK => CLK, Q => n_3168, QN 
                           => n51970);
   clk_r_REG16534_S1 : DFF_X1 port map( D => n3230, CK => CLK, Q => n_3169, QN 
                           => n51969);
   clk_r_REG14771_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n_3170, QN 
                           => n51968);
   clk_r_REG14769_S1 : DFF_X1 port map( D => n3331, CK => CLK, Q => n_3171, QN 
                           => n51967);
   clk_r_REG14989_S1 : DFF_X1 port map( D => n3520, CK => CLK, Q => n_3172, QN 
                           => n51966);
   clk_r_REG15620_S1 : DFF_X1 port map( D => n2984, CK => CLK, Q => n_3173, QN 
                           => n51965);
   clk_r_REG15634_S1 : DFF_X1 port map( D => n3041, CK => CLK, Q => n_3174, QN 
                           => n51964);
   clk_r_REG14377_S1 : DFF_X1 port map( D => n3424, CK => CLK, Q => n_3175, QN 
                           => n51963);
   clk_r_REG15570_S1 : DFF_X1 port map( D => n3009, CK => CLK, Q => n_3176, QN 
                           => n51962);
   clk_r_REG15037_S1 : DFF_X1 port map( D => n3496, CK => CLK, Q => n_3177, QN 
                           => n51961);
   clk_r_REG15568_S1 : DFF_X1 port map( D => n3010, CK => CLK, Q => n_3178, QN 
                           => n51960);
   clk_r_REG14425_S1 : DFF_X1 port map( D => n3400, CK => CLK, Q => n_3179, QN 
                           => n51959);
   clk_r_REG16195_S1 : DFF_X1 port map( D => n2824, CK => CLK, Q => n_3180, QN 
                           => n51958);
   clk_r_REG14847_S1 : DFF_X1 port map( D => n3488, CK => CLK, Q => n_3181, QN 
                           => n51957);
   clk_r_REG16397_S1 : DFF_X1 port map( D => n3106, CK => CLK, Q => n_3182, QN 
                           => n51956);
   clk_r_REG14895_S1 : DFF_X1 port map( D => n3464, CK => CLK, Q => n_3183, QN 
                           => n51955);
   clk_r_REG14987_S1 : DFF_X1 port map( D => n3521, CK => CLK, Q => n_3184, QN 
                           => n51954);
   clk_r_REG14985_S1 : DFF_X1 port map( D => n3522, CK => CLK, Q => n_3185, QN 
                           => n51953);
   clk_r_REG14983_S1 : DFF_X1 port map( D => n3523, CK => CLK, Q => n_3186, QN 
                           => n51952);
   clk_r_REG14981_S1 : DFF_X1 port map( D => n3524, CK => CLK, Q => n_3187, QN 
                           => n51951);
   clk_r_REG15318_S1 : DFF_X1 port map( D => n3360, CK => CLK, Q => n_3188, QN 
                           => n51950);
   clk_r_REG14375_S1 : DFF_X1 port map( D => n3425, CK => CLK, Q => n_3189, QN 
                           => n51949);
   clk_r_REG14707_S1 : DFF_X1 port map( D => n3456, CK => CLK, Q => n_3190, QN 
                           => n51948);
   clk_r_REG14845_S1 : DFF_X1 port map( D => n3489, CK => CLK, Q => n_3191, QN 
                           => n51947);
   clk_r_REG14843_S1 : DFF_X1 port map( D => n3490, CK => CLK, Q => n_3192, QN 
                           => n51946);
   clk_r_REG14373_S1 : DFF_X1 port map( D => n3426, CK => CLK, Q => n_3193, QN 
                           => n51945);
   clk_r_REG14371_S1 : DFF_X1 port map( D => n3427, CK => CLK, Q => n_3194, QN 
                           => n51944);
   clk_r_REG14755_S1 : DFF_X1 port map( D => n3432, CK => CLK, Q => n_3195, QN 
                           => n51943);
   clk_r_REG14705_S1 : DFF_X1 port map( D => n3457, CK => CLK, Q => n_3196, QN 
                           => n51942);
   clk_r_REG14841_S1 : DFF_X1 port map( D => n3491, CK => CLK, Q => n_3197, QN 
                           => n51941);
   clk_r_REG16087_S1 : DFF_X1 port map( D => n2814, CK => CLK, Q => n_3198, QN 
                           => n51940);
   clk_r_REG14369_S1 : DFF_X1 port map( D => n3428, CK => CLK, Q => n_3199, QN 
                           => n51939);
   clk_r_REG15106_S1 : DFF_X1 port map( D => n3047, CK => CLK, Q => n_3200, QN 
                           => n51938);
   clk_r_REG14839_S1 : DFF_X1 port map( D => n3492, CK => CLK, Q => n_3201, QN 
                           => n51937);
   clk_r_REG14703_S1 : DFF_X1 port map( D => n3458, CK => CLK, Q => n_3202, QN 
                           => n51936);
   clk_r_REG15366_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n_3203, QN 
                           => n51935);
   clk_r_REG14631_S1 : DFF_X1 port map( D => n3392, CK => CLK, Q => n_3204, QN 
                           => n51934);
   clk_r_REG14701_S1 : DFF_X1 port map( D => n3459, CK => CLK, Q => n_3205, QN 
                           => n51933);
   clk_r_REG16624_S1 : DFF_X1 port map( D => n3553, CK => CLK, Q => n_3206, QN 
                           => n51932);
   clk_r_REG16622_S1 : DFF_X1 port map( D => n3554, CK => CLK, Q => n_3207, QN 
                           => n51931);
   clk_r_REG14699_S1 : DFF_X1 port map( D => n3460, CK => CLK, Q => n_3208, QN 
                           => n51930);
   clk_r_REG14679_S1 : DFF_X1 port map( D => n3368, CK => CLK, Q => n_3209, QN 
                           => n51929);
   clk_r_REG15056_S1 : DFF_X1 port map( D => n3072, CK => CLK, Q => n_3210, QN 
                           => n51928);
   clk_r_REG16219_S1 : DFF_X1 port map( D => n2876, CK => CLK, Q => n_3211, QN 
                           => n51927);
   clk_r_REG15472_S1 : DFF_X1 port map( D => n2941, CK => CLK, Q => n_3212, QN 
                           => n51926);
   clk_r_REG15560_S1 : DFF_X1 port map( D => n2950, CK => CLK, Q => n_3213, QN 
                           => n51925);
   clk_r_REG15558_S1 : DFF_X1 port map( D => n2951, CK => CLK, Q => n_3214, QN 
                           => n51924);
   clk_r_REG16085_S1 : DFF_X1 port map( D => n2815, CK => CLK, Q => n_3215, QN 
                           => n51923);
   clk_r_REG15508_S1 : DFF_X1 port map( D => n2976, CK => CLK, Q => n_3216, QN 
                           => n51922);
   clk_r_REG15428_S1 : DFF_X1 port map( D => n2888, CK => CLK, Q => n_3217, QN 
                           => n51921);
   clk_r_REG15378_S1 : DFF_X1 port map( D => n2913, CK => CLK, Q => n_3218, QN 
                           => n51920);
   clk_r_REG16217_S1 : DFF_X1 port map( D => n2877, CK => CLK, Q => n_3219, QN 
                           => n51919);
   clk_r_REG16215_S1 : DFF_X1 port map( D => n2878, CK => CLK, Q => n_3220, QN 
                           => n51918);
   clk_r_REG14629_S1 : DFF_X1 port map( D => n3393, CK => CLK, Q => n_3221, QN 
                           => n51917);
   clk_r_REG15470_S1 : DFF_X1 port map( D => n2942, CK => CLK, Q => n_3222, QN 
                           => n51916);
   clk_r_REG15104_S1 : DFF_X1 port map( D => n3048, CK => CLK, Q => n_3223, QN 
                           => n51915);
   clk_r_REG15054_S1 : DFF_X1 port map( D => n3073, CK => CLK, Q => n_3224, QN 
                           => n51914);
   clk_r_REG16213_S1 : DFF_X1 port map( D => n2879, CK => CLK, Q => n_3225, QN 
                           => n51913);
   clk_r_REG15316_S1 : DFF_X1 port map( D => n3361, CK => CLK, Q => n_3226, QN 
                           => n51912);
   clk_r_REG15314_S1 : DFF_X1 port map( D => n3362, CK => CLK, Q => n_3227, QN 
                           => n51911);
   clk_r_REG15312_S1 : DFF_X1 port map( D => n3363, CK => CLK, Q => n_3228, QN 
                           => n51910);
   clk_r_REG16263_S1 : DFF_X1 port map( D => n2854, CK => CLK, Q => n_3229, QN 
                           => n51909);
   clk_r_REG14627_S1 : DFF_X1 port map( D => n3394, CK => CLK, Q => n_3230, QN 
                           => n51908);
   clk_r_REG14625_S1 : DFF_X1 port map( D => n3395, CK => CLK, Q => n_3231, QN 
                           => n51907);
   clk_r_REG16135_S1 : DFF_X1 port map( D => n2790, CK => CLK, Q => n_3232, QN 
                           => n51906);
   clk_r_REG15556_S1 : DFF_X1 port map( D => n2952, CK => CLK, Q => n_3233, QN 
                           => n51905);
   clk_r_REG15506_S1 : DFF_X1 port map( D => n2977, CK => CLK, Q => n_3234, QN 
                           => n51904);
   clk_r_REG16145_S1 : DFF_X1 port map( D => n2849, CK => CLK, Q => n_3235, QN 
                           => n51903);
   clk_r_REG14623_S1 : DFF_X1 port map( D => n3396, CK => CLK, Q => n_3236, QN 
                           => n51902);
   clk_r_REG15310_S1 : DFF_X1 port map( D => n3364, CK => CLK, Q => n_3237, QN 
                           => n51901);
   clk_r_REG16133_S1 : DFF_X1 port map( D => n2791, CK => CLK, Q => n_3238, QN 
                           => n51900);
   clk_r_REG15052_S1 : DFF_X1 port map( D => n3074, CK => CLK, Q => n_3239, QN 
                           => n51899);
   clk_r_REG16458_S1 : DFF_X1 port map( D => n3140, CK => CLK, Q => n_3240, QN 
                           => n51898);
   clk_r_REG16395_S1 : DFF_X1 port map( D => n3107, CK => CLK, Q => n_3241, QN 
                           => n51897);
   clk_r_REG15050_S1 : DFF_X1 port map( D => n3075, CK => CLK, Q => n_3242, QN 
                           => n51896);
   clk_r_REG15504_S1 : DFF_X1 port map( D => n2978, CK => CLK, Q => n_3243, QN 
                           => n51895);
   clk_r_REG15468_S1 : DFF_X1 port map( D => n2943, CK => CLK, Q => n_3244, QN 
                           => n51894);
   clk_r_REG15376_S1 : DFF_X1 port map( D => n2914, CK => CLK, Q => n_3245, QN 
                           => n51893);
   clk_r_REG16143_S1 : DFF_X1 port map( D => n2850, CK => CLK, Q => n_3246, QN 
                           => n51892);
   clk_r_REG14767_S1 : DFF_X1 port map( D => n3332, CK => CLK, Q => n_3247, QN 
                           => n51891);
   clk_r_REG14078_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n_3248, QN 
                           => n51890);
   clk_r_REG13836_S1 : DFF_X1 port map( D => n3365, CK => CLK, Q => n_3249, QN 
                           => n51889);
   clk_r_REG14821_S1 : DFF_X1 port map( D => n3305, CK => CLK, Q => n_3250, QN 
                           => n51888);
   clk_r_REG14819_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n_3251, QN 
                           => n51887);
   clk_r_REG14159_S1 : DFF_X1 port map( D => n3429, CK => CLK, Q => n_3252, QN 
                           => n51886);
   clk_r_REG14119_S1 : DFF_X1 port map( D => n3461, CK => CLK, Q => n_3253, QN 
                           => n51885);
   clk_r_REG15364_S1 : DFF_X1 port map( D => n3337, CK => CLK, Q => n_3254, QN 
                           => n51884);
   clk_r_REG14065_S1 : DFF_X1 port map( D => n3493, CK => CLK, Q => n_3255, QN 
                           => n51883);
   clk_r_REG14893_S1 : DFF_X1 port map( D => n3465, CK => CLK, Q => n_3256, QN 
                           => n51882);
   clk_r_REG14817_S1 : DFF_X1 port map( D => n3307, CK => CLK, Q => n_3257, QN 
                           => n51881);
   clk_r_REG14891_S1 : DFF_X1 port map( D => n3466, CK => CLK, Q => n_3258, QN 
                           => n51880);
   clk_r_REG14889_S1 : DFF_X1 port map( D => n3467, CK => CLK, Q => n_3259, QN 
                           => n51879);
   clk_r_REG15362_S1 : DFF_X1 port map( D => n3338, CK => CLK, Q => n_3260, QN 
                           => n51878);
   clk_r_REG15360_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n_3261, QN 
                           => n51877);
   clk_r_REG14887_S1 : DFF_X1 port map( D => n3468, CK => CLK, Q => n_3262, QN 
                           => n51876);
   clk_r_REG14140_S1 : DFF_X1 port map( D => n3397, CK => CLK, Q => n_3263, QN 
                           => n51875);
   clk_r_REG14815_S1 : DFF_X1 port map( D => n3308, CK => CLK, Q => n_3264, QN 
                           => n51874);
   clk_r_REG15358_S1 : DFF_X1 port map( D => n3340, CK => CLK, Q => n_3265, QN 
                           => n51873);
   clk_r_REG15356_S1 : DFF_X1 port map( D => n3341, CK => CLK, Q => n_3266, QN 
                           => n51872);
   clk_r_REG16141_S1 : DFF_X1 port map( D => n2851, CK => CLK, Q => n_3267, QN 
                           => n51871);
   clk_r_REG14677_S1 : DFF_X1 port map( D => n3369, CK => CLK, Q => n_3268, QN 
                           => n51870);
   clk_r_REG14423_S1 : DFF_X1 port map( D => n3401, CK => CLK, Q => n_3269, QN 
                           => n51869);
   clk_r_REG15354_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n_3270, QN 
                           => n51868);
   clk_r_REG16083_S1 : DFF_X1 port map( D => n2816, CK => CLK, Q => n_3271, QN 
                           => n51867);
   clk_r_REG16139_S1 : DFF_X1 port map( D => n2852, CK => CLK, Q => n_3272, QN 
                           => n51866);
   clk_r_REG14675_S1 : DFF_X1 port map( D => n3370, CK => CLK, Q => n_3273, QN 
                           => n51865);
   clk_r_REG16081_S1 : DFF_X1 port map( D => n2817, CK => CLK, Q => n_3274, QN 
                           => n51864);
   clk_r_REG14813_S1 : DFF_X1 port map( D => n3309, CK => CLK, Q => n_3275, QN 
                           => n51863);
   clk_r_REG14753_S1 : DFF_X1 port map( D => n3433, CK => CLK, Q => n_3276, QN 
                           => n51862);
   clk_r_REG14673_S1 : DFF_X1 port map( D => n3371, CK => CLK, Q => n_3277, QN 
                           => n51861);
   clk_r_REG14671_S1 : DFF_X1 port map( D => n3372, CK => CLK, Q => n_3278, QN 
                           => n51860);
   clk_r_REG14010_S1 : DFF_X1 port map( D => n3525, CK => CLK, Q => n_3279, QN 
                           => n51859);
   clk_r_REG15035_S1 : DFF_X1 port map( D => n3497, CK => CLK, Q => n_3280, QN 
                           => n51858);
   clk_r_REG14669_S1 : DFF_X1 port map( D => n3373, CK => CLK, Q => n_3281, QN 
                           => n51857);
   clk_r_REG14421_S1 : DFF_X1 port map( D => n3402, CK => CLK, Q => n_3282, QN 
                           => n51856);
   clk_r_REG14751_S1 : DFF_X1 port map( D => n3434, CK => CLK, Q => n_3283, QN 
                           => n51855);
   clk_r_REG14885_S1 : DFF_X1 port map( D => n3469, CK => CLK, Q => n_3284, QN 
                           => n51854);
   clk_r_REG15033_S1 : DFF_X1 port map( D => n3498, CK => CLK, Q => n_3285, QN 
                           => n51853);
   clk_r_REG15374_S1 : DFF_X1 port map( D => n2915, CK => CLK, Q => n_3286, QN 
                           => n51852);
   clk_r_REG14811_S1 : DFF_X1 port map( D => n3310, CK => CLK, Q => n_3287, QN 
                           => n51851);
   clk_r_REG14667_S1 : DFF_X1 port map( D => n3374, CK => CLK, Q => n_3288, QN 
                           => n51850);
   clk_r_REG14419_S1 : DFF_X1 port map( D => n3403, CK => CLK, Q => n_3289, QN 
                           => n51849);
   clk_r_REG14417_S1 : DFF_X1 port map( D => n3404, CK => CLK, Q => n_3290, QN 
                           => n51848);
   clk_r_REG14415_S1 : DFF_X1 port map( D => n3405, CK => CLK, Q => n_3291, QN 
                           => n51847);
   clk_r_REG14413_S1 : DFF_X1 port map( D => n3406, CK => CLK, Q => n_3292, QN 
                           => n51846);
   clk_r_REG14749_S1 : DFF_X1 port map( D => n3435, CK => CLK, Q => n_3293, QN 
                           => n51845);
   clk_r_REG14747_S1 : DFF_X1 port map( D => n3436, CK => CLK, Q => n_3294, QN 
                           => n51844);
   clk_r_REG15031_S1 : DFF_X1 port map( D => n3499, CK => CLK, Q => n_3295, QN 
                           => n51843);
   clk_r_REG15029_S1 : DFF_X1 port map( D => n3500, CK => CLK, Q => n_3296, QN 
                           => n51842);
   clk_r_REG15027_S1 : DFF_X1 port map( D => n3501, CK => CLK, Q => n_3297, QN 
                           => n51841);
   clk_r_REG14745_S1 : DFF_X1 port map( D => n3437, CK => CLK, Q => n_3298, QN 
                           => n51840);
   clk_r_REG14743_S1 : DFF_X1 port map( D => n3438, CK => CLK, Q => n_3299, QN 
                           => n51839);
   clk_r_REG14883_S1 : DFF_X1 port map( D => n3470, CK => CLK, Q => n_3300, QN 
                           => n51838);
   clk_r_REG15025_S1 : DFF_X1 port map( D => n3502, CK => CLK, Q => n_3301, QN 
                           => n51837);
   clk_r_REG14741_S1 : DFF_X1 port map( D => n3439, CK => CLK, Q => n_3302, QN 
                           => n51836);
   clk_r_REG14881_S1 : DFF_X1 port map( D => n3471, CK => CLK, Q => n_3303, QN 
                           => n51835);
   clk_r_REG15023_S1 : DFF_X1 port map( D => n3503, CK => CLK, Q => n_3304, QN 
                           => n51834);
   clk_r_REG16532_S1 : DFF_X1 port map( D => n3231, CK => CLK, Q => n_3305, QN 
                           => n51833);
   clk_r_REG14665_S1 : DFF_X1 port map( D => n3375, CK => CLK, Q => n_3306, QN 
                           => n51832);
   clk_r_REG14411_S1 : DFF_X1 port map( D => n3407, CK => CLK, Q => n_3307, QN 
                           => n51831);
   clk_r_REG14809_S1 : DFF_X1 port map( D => n3311, CK => CLK, Q => n_3308, QN 
                           => n51830);
   clk_r_REG15172_S1 : DFF_X1 port map( D => n3144, CK => CLK, Q => n_3309, QN 
                           => n51829);
   clk_r_REG15352_S1 : DFF_X1 port map( D => n3343, CK => CLK, Q => n_3310, QN 
                           => n51828);
   clk_r_REG16620_S1 : DFF_X1 port map( D => n3555, CK => CLK, Q => n_3311, QN 
                           => n51827);
   clk_r_REG16393_S1 : DFF_X1 port map( D => n3108, CK => CLK, Q => n_3312, QN 
                           => n51826);
   clk_r_REG13673_S1 : DFF_X1 port map( D => n3141, CK => CLK, Q => n_3313, QN 
                           => n51825);
   clk_r_REG15632_S1 : DFF_X1 port map( D => n3042, CK => CLK, Q => n_3314, QN 
                           => n51824);
   clk_r_REG15048_S1 : DFF_X1 port map( D => n3076, CK => CLK, Q => n_3315, QN 
                           => n51823);
   clk_r_REG15502_S1 : DFF_X1 port map( D => n2979, CK => CLK, Q => n_3316, QN 
                           => n51822);
   clk_r_REG15466_S1 : DFF_X1 port map( D => n2928, CK => CLK, Q => n_3317, QN 
                           => n51821);
   clk_r_REG15372_S1 : DFF_X1 port map( D => n2916, CK => CLK, Q => n_3318, QN 
                           => n51820);
   clk_r_REG16261_S1 : DFF_X1 port map( D => n2855, CK => CLK, Q => n_3319, QN 
                           => n51819);
   clk_r_REG13727_S1 : DFF_X1 port map( D => n2853, CK => CLK, Q => n_3320, QN 
                           => n51818);
   clk_r_REG16131_S1 : DFF_X1 port map( D => n2792, CK => CLK, Q => n_3321, QN 
                           => n51817);
   clk_r_REG15630_S1 : DFF_X1 port map( D => n3043, CK => CLK, Q => n_3322, QN 
                           => n51816);
   clk_r_REG15628_S1 : DFF_X1 port map( D => n3044, CK => CLK, Q => n_3323, QN 
                           => n51815);
   clk_r_REG15566_S1 : DFF_X1 port map( D => n3011, CK => CLK, Q => n_3324, QN 
                           => n51814);
   clk_r_REG13794_S1 : DFF_X1 port map( D => n3045, CK => CLK, Q => n_3325, QN 
                           => n51813);
   clk_r_REG15682_S1 : DFF_X1 port map( D => n3017, CK => CLK, Q => n_3326, QN 
                           => n51812);
   clk_r_REG15680_S1 : DFF_X1 port map( D => n3018, CK => CLK, Q => n_3327, QN 
                           => n51811);
   clk_r_REG15678_S1 : DFF_X1 port map( D => n3019, CK => CLK, Q => n_3328, QN 
                           => n51810);
   clk_r_REG15676_S1 : DFF_X1 port map( D => n3020, CK => CLK, Q => n_3329, QN 
                           => n51809);
   clk_r_REG15564_S1 : DFF_X1 port map( D => n3012, CK => CLK, Q => n_3330, QN 
                           => n51808);
   clk_r_REG13803_S1 : DFF_X1 port map( D => n3013, CK => CLK, Q => n_3331, QN 
                           => n51807);
   clk_r_REG15618_S1 : DFF_X1 port map( D => n2985, CK => CLK, Q => n_3332, QN 
                           => n51806);
   clk_r_REG15616_S1 : DFF_X1 port map( D => n2986, CK => CLK, Q => n_3333, QN 
                           => n51805);
   clk_r_REG15614_S1 : DFF_X1 port map( D => n2987, CK => CLK, Q => n_3334, QN 
                           => n51804);
   clk_r_REG15612_S1 : DFF_X1 port map( D => n2988, CK => CLK, Q => n_3335, QN 
                           => n51803);
   clk_r_REG15610_S1 : DFF_X1 port map( D => n2989, CK => CLK, Q => n_3336, QN 
                           => n51802);
   clk_r_REG13868_S1 : DFF_X1 port map( D => n3205, CK => CLK, Q => n_3337, QN 
                           => n51801);
   clk_r_REG13824_S1 : DFF_X1 port map( D => n2917, CK => CLK, Q => n_3338, QN 
                           => n51800);
   clk_r_REG16211_S1 : DFF_X1 port map( D => n2880, CK => CLK, Q => n_3339, QN 
                           => n51799);
   clk_r_REG16259_S1 : DFF_X1 port map( D => n2856, CK => CLK, Q => n_3340, QN 
                           => n51798);
   clk_r_REG16209_S1 : DFF_X1 port map( D => n2881, CK => CLK, Q => n_3341, QN 
                           => n51797);
   clk_r_REG16207_S1 : DFF_X1 port map( D => n2882, CK => CLK, Q => n_3342, QN 
                           => n51796);
   clk_r_REG16205_S1 : DFF_X1 port map( D => n2883, CK => CLK, Q => n_3343, QN 
                           => n51795);
   clk_r_REG16203_S1 : DFF_X1 port map( D => n2884, CK => CLK, Q => n_3344, QN 
                           => n51794);
   clk_r_REG13720_S1 : DFF_X1 port map( D => n2885, CK => CLK, Q => n_3345, QN 
                           => n51793);
   clk_r_REG16582_S1 : DFF_X1 port map( D => n3206, CK => CLK, Q => n_3346, QN 
                           => n51792);
   clk_r_REG15303_S1 : DFF_X1 port map( D => n3240, CK => CLK, Q => n_3347, QN 
                           => n51791);
   clk_r_REG14031_S1 : DFF_X1 port map( D => n3301, CK => CLK, Q => n_3348, QN 
                           => n51790);
   clk_r_REG15237_S1 : DFF_X1 port map( D => n3177, CK => CLK, Q => n_3349, QN 
                           => n51789);
   clk_r_REG15122_S1 : DFF_X1 port map( D => n3169, CK => CLK, Q => n_3350, QN 
                           => n51788);
   clk_r_REG16512_S1 : DFF_X1 port map( D => n3113, CK => CLK, Q => n_3351, QN 
                           => n51787);
   clk_r_REG13687_S1 : DFF_X1 port map( D => n3109, CK => CLK, Q => n_3352, QN 
                           => n51786);
   clk_r_REG13917_S1 : DFF_X1 port map( D => n3077, CK => CLK, Q => n_3353, QN 
                           => n51785);
   clk_r_REG15500_S1 : DFF_X1 port map( D => n2980, CK => CLK, Q => n_3354, QN 
                           => n51784);
   clk_r_REG15464_S1 : DFF_X1 port map( D => n2927, CK => CLK, Q => n_3355, QN 
                           => n51783);
   clk_r_REG14961_S1 : DFF_X1 port map( D => n3273, CK => CLK, Q => n_3356, QN 
                           => n51782);
   clk_r_REG15253_S1 : DFF_X1 port map( D => n3265, CK => CLK, Q => n_3357, QN 
                           => n51781);
   clk_r_REG16580_S1 : DFF_X1 port map( D => n3207, CK => CLK, Q => n_3358, QN 
                           => n51780);
   clk_r_REG15235_S1 : DFF_X1 port map( D => n3178, CK => CLK, Q => n_3359, QN 
                           => n51779);
   clk_r_REG15120_S1 : DFF_X1 port map( D => n3170, CK => CLK, Q => n_3360, QN 
                           => n51778);
   clk_r_REG16079_S1 : DFF_X1 port map( D => n2818, CK => CLK, Q => n_3361, QN 
                           => n51777);
   clk_r_REG14959_S1 : DFF_X1 port map( D => n3274, CK => CLK, Q => n_3362, QN 
                           => n51776);
   clk_r_REG15251_S1 : DFF_X1 port map( D => n3266, CK => CLK, Q => n_3363, QN 
                           => n51775);
   clk_r_REG15233_S1 : DFF_X1 port map( D => n3179, CK => CLK, Q => n_3364, QN 
                           => n51774);
   clk_r_REG15231_S1 : DFF_X1 port map( D => n3180, CK => CLK, Q => n_3365, QN 
                           => n51773);
   clk_r_REG15229_S1 : DFF_X1 port map( D => n3181, CK => CLK, Q => n_3366, QN 
                           => n51772);
   clk_r_REG15227_S1 : DFF_X1 port map( D => n3182, CK => CLK, Q => n_3367, QN 
                           => n51771);
   clk_r_REG15118_S1 : DFF_X1 port map( D => n3171, CK => CLK, Q => n_3368, QN 
                           => n51770);
   clk_r_REG16510_S1 : DFF_X1 port map( D => n3114, CK => CLK, Q => n_3369, QN 
                           => n51769);
   clk_r_REG16447_S1 : DFF_X1 port map( D => n3081, CK => CLK, Q => n_3370, QN 
                           => n51768);
   clk_r_REG15102_S1 : DFF_X1 port map( D => n3049, CK => CLK, Q => n_3371, QN 
                           => n51767);
   clk_r_REG15608_S1 : DFF_X1 port map( D => n2990, CK => CLK, Q => n_3372, QN 
                           => n51766);
   clk_r_REG13810_S1 : DFF_X1 port map( D => n2981, CK => CLK, Q => n_3373, QN 
                           => n51765);
   clk_r_REG15444_S1 : DFF_X1 port map( D => n2944, CK => CLK, Q => n_3374, QN 
                           => n51764);
   clk_r_REG15426_S1 : DFF_X1 port map( D => n2889, CK => CLK, Q => n_3375, QN 
                           => n51763);
   clk_r_REG14879_S1 : DFF_X1 port map( D => n3472, CK => CLK, Q => n_3376, QN 
                           => n51762);
   clk_r_REG16530_S1 : DFF_X1 port map( D => n3232, CK => CLK, Q => n_3377, QN 
                           => n51761);
   clk_r_REG16193_S1 : DFF_X1 port map( D => n2825, CK => CLK, Q => n_3378, QN 
                           => n51760);
   clk_r_REG15116_S1 : DFF_X1 port map( D => n3172, CK => CLK, Q => n_3379, QN 
                           => n51759);
   clk_r_REG13904_S1 : DFF_X1 port map( D => n3173, CK => CLK, Q => n_3380, QN 
                           => n51758);
   clk_r_REG15170_S1 : DFF_X1 port map( D => n3145, CK => CLK, Q => n_3381, QN 
                           => n51757);
   clk_r_REG16077_S1 : DFF_X1 port map( D => n2819, CK => CLK, Q => n_3382, QN 
                           => n51756);
   clk_r_REG16508_S1 : DFF_X1 port map( D => n3115, CK => CLK, Q => n_3383, QN 
                           => n51755);
   clk_r_REG16578_S1 : DFF_X1 port map( D => n3208, CK => CLK, Q => n_3384, QN 
                           => n51754);
   clk_r_REG16506_S1 : DFF_X1 port map( D => n3116, CK => CLK, Q => n_3385, QN 
                           => n51753);
   clk_r_REG16528_S1 : DFF_X1 port map( D => n3233, CK => CLK, Q => n_3386, QN 
                           => n51752);
   clk_r_REG15249_S1 : DFF_X1 port map( D => n3267, CK => CLK, Q => n_3387, QN 
                           => n51751);
   clk_r_REG16504_S1 : DFF_X1 port map( D => n3117, CK => CLK, Q => n_3388, QN 
                           => n51750);
   clk_r_REG14957_S1 : DFF_X1 port map( D => n3275, CK => CLK, Q => n_3389, QN 
                           => n51749);
   clk_r_REG15247_S1 : DFF_X1 port map( D => n3268, CK => CLK, Q => n_3390, QN 
                           => n51748);
   clk_r_REG16445_S1 : DFF_X1 port map( D => n3082, CK => CLK, Q => n_3391, QN 
                           => n51747);
   clk_r_REG14955_S1 : DFF_X1 port map( D => n3276, CK => CLK, Q => n_3392, QN 
                           => n51746);
   clk_r_REG13849_S1 : DFF_X1 port map( D => n3269, CK => CLK, Q => n_3393, QN 
                           => n51745);
   clk_r_REG16526_S1 : DFF_X1 port map( D => n3234, CK => CLK, Q => n_3394, QN 
                           => n51744);
   clk_r_REG15021_S1 : DFF_X1 port map( D => n3504, CK => CLK, Q => n_3395, QN 
                           => n51743);
   clk_r_REG15225_S1 : DFF_X1 port map( D => n3183, CK => CLK, Q => n_3396, QN 
                           => n51742);
   clk_r_REG15168_S1 : DFF_X1 port map( D => n3146, CK => CLK, Q => n_3397, QN 
                           => n51741);
   clk_r_REG16502_S1 : DFF_X1 port map( D => n3118, CK => CLK, Q => n_3398, QN 
                           => n51740);
   clk_r_REG16443_S1 : DFF_X1 port map( D => n3083, CK => CLK, Q => n_3399, QN 
                           => n51739);
   clk_r_REG15100_S1 : DFF_X1 port map( D => n3050, CK => CLK, Q => n_3400, QN 
                           => n51738);
   clk_r_REG15098_S1 : DFF_X1 port map( D => n3051, CK => CLK, Q => n_3401, QN 
                           => n51737);
   clk_r_REG15096_S1 : DFF_X1 port map( D => n3052, CK => CLK, Q => n_3402, QN 
                           => n51736);
   clk_r_REG15554_S1 : DFF_X1 port map( D => n2953, CK => CLK, Q => n_3403, QN 
                           => n51735);
   clk_r_REG15094_S1 : DFF_X1 port map( D => n3053, CK => CLK, Q => n_3404, QN 
                           => n51734);
   clk_r_REG16524_S1 : DFF_X1 port map( D => n3235, CK => CLK, Q => n_3405, QN 
                           => n51733);
   clk_r_REG14409_S1 : DFF_X1 port map( D => n3408, CK => CLK, Q => n_3406, QN 
                           => n51732);
   clk_r_REG15301_S1 : DFF_X1 port map( D => n3241, CK => CLK, Q => n_3407, QN 
                           => n51731);
   clk_r_REG15299_S1 : DFF_X1 port map( D => n3242, CK => CLK, Q => n_3408, QN 
                           => n51730);
   clk_r_REG15297_S1 : DFF_X1 port map( D => n3243, CK => CLK, Q => n_3409, QN 
                           => n51729);
   clk_r_REG14953_S1 : DFF_X1 port map( D => n3277, CK => CLK, Q => n_3410, QN 
                           => n51728);
   clk_r_REG14951_S1 : DFF_X1 port map( D => n3278, CK => CLK, Q => n_3411, QN 
                           => n51727);
   clk_r_REG16522_S1 : DFF_X1 port map( D => n3236, CK => CLK, Q => n_3412, QN 
                           => n51726);
   clk_r_REG15092_S1 : DFF_X1 port map( D => n3054, CK => CLK, Q => n_3413, QN 
                           => n51725);
   clk_r_REG14949_S1 : DFF_X1 port map( D => n3279, CK => CLK, Q => n_3414, QN 
                           => n51724);
   clk_r_REG16075_S1 : DFF_X1 port map( D => n2820, CK => CLK, Q => n_3415, QN 
                           => n51723);
   clk_r_REG16191_S1 : DFF_X1 port map( D => n2826, CK => CLK, Q => n_3416, QN 
                           => n51722);
   clk_r_REG15350_S1 : DFF_X1 port map( D => n3344, CK => CLK, Q => n_3417, QN 
                           => n51721);
   clk_r_REG16441_S1 : DFF_X1 port map( D => n3084, CK => CLK, Q => n_3418, QN 
                           => n51720);
   clk_r_REG14947_S1 : DFF_X1 port map( D => n3280, CK => CLK, Q => n_3419, QN 
                           => n51719);
   clk_r_REG15462_S1 : DFF_X1 port map( D => n2926, CK => CLK, Q => n_3420, QN 
                           => n51718);
   clk_r_REG15552_S1 : DFF_X1 port map( D => n2954, CK => CLK, Q => n_3421, QN 
                           => n51717);
   clk_r_REG15424_S1 : DFF_X1 port map( D => n2890, CK => CLK, Q => n_3422, QN 
                           => n51716);
   clk_r_REG15422_S1 : DFF_X1 port map( D => n2891, CK => CLK, Q => n_3423, QN 
                           => n51715);
   clk_r_REG15420_S1 : DFF_X1 port map( D => n2892, CK => CLK, Q => n_3424, QN 
                           => n51714);
   clk_r_REG15442_S1 : DFF_X1 port map( D => n2945, CK => CLK, Q => n_3425, QN 
                           => n51713);
   clk_r_REG16500_S1 : DFF_X1 port map( D => n3119, CK => CLK, Q => n_3426, QN 
                           => n51712);
   clk_r_REG15440_S1 : DFF_X1 port map( D => n2946, CK => CLK, Q => n_3427, QN 
                           => n51711);
   clk_r_REG16439_S1 : DFF_X1 port map( D => n3085, CK => CLK, Q => n_3428, QN 
                           => n51710);
   clk_r_REG13734_S1 : DFF_X1 port map( D => n2821, CK => CLK, Q => n_3429, QN 
                           => n51709);
   clk_r_REG14663_S1 : DFF_X1 port map( D => n3376, CK => CLK, Q => n_3430, QN 
                           => n51708);
   clk_r_REG16189_S1 : DFF_X1 port map( D => n2827, CK => CLK, Q => n_3431, QN 
                           => n51707);
   clk_r_REG15418_S1 : DFF_X1 port map( D => n2893, CK => CLK, Q => n_3432, QN 
                           => n51706);
   clk_r_REG15166_S1 : DFF_X1 port map( D => n3147, CK => CLK, Q => n_3433, QN 
                           => n51705);
   clk_r_REG16187_S1 : DFF_X1 port map( D => n2828, CK => CLK, Q => n_3434, QN 
                           => n51704);
   clk_r_REG16437_S1 : DFF_X1 port map( D => n3086, CK => CLK, Q => n_3435, QN 
                           => n51703);
   clk_r_REG16257_S1 : DFF_X1 port map( D => n2857, CK => CLK, Q => n_3436, QN 
                           => n51702);
   clk_r_REG15550_S1 : DFF_X1 port map( D => n2955, CK => CLK, Q => n_3437, QN 
                           => n51701);
   clk_r_REG15438_S1 : DFF_X1 port map( D => n2947, CK => CLK, Q => n_3438, QN 
                           => n51700);
   clk_r_REG16129_S1 : DFF_X1 port map( D => n2793, CK => CLK, Q => n_3439, QN 
                           => n51699);
   clk_r_REG15548_S1 : DFF_X1 port map( D => n2956, CK => CLK, Q => n_3440, QN 
                           => n51698);
   clk_r_REG15546_S1 : DFF_X1 port map( D => n2957, CK => CLK, Q => n_3441, QN 
                           => n51697);
   clk_r_REG15674_S1 : DFF_X1 port map( D => n3021, CK => CLK, Q => n_3442, QN 
                           => n51696);
   clk_r_REG15223_S1 : DFF_X1 port map( D => n3184, CK => CLK, Q => n_3443, QN 
                           => n51695);
   clk_r_REG16185_S1 : DFF_X1 port map( D => n2829, CK => CLK, Q => n_3444, QN 
                           => n51694);
   clk_r_REG14739_S1 : DFF_X1 port map( D => n3440, CK => CLK, Q => n_3445, QN 
                           => n51693);
   clk_r_REG16127_S1 : DFF_X1 port map( D => n2794, CK => CLK, Q => n_3446, QN 
                           => n51692);
   clk_r_REG15436_S1 : DFF_X1 port map( D => n2948, CK => CLK, Q => n_3447, QN 
                           => n51691);
   clk_r_REG16618_S1 : DFF_X1 port map( D => n3556, CK => CLK, Q => n_3448, QN 
                           => n51690);
   clk_r_REG13648_S1 : DFF_X1 port map( D => n3557, CK => CLK, Q => n_3449, QN 
                           => n51689);
   clk_r_REG16672_S1 : DFF_X1 port map( D => n3529, CK => CLK, Q => n_3450, QN 
                           => n51688);
   clk_r_REG16670_S1 : DFF_X1 port map( D => n3530, CK => CLK, Q => n_3451, QN 
                           => n51687);
   clk_r_REG16668_S1 : DFF_X1 port map( D => n3531, CK => CLK, Q => n_3452, QN 
                           => n51686);
   clk_r_REG16666_S1 : DFF_X1 port map( D => n3532, CK => CLK, Q => n_3453, QN 
                           => n51685);
   clk_r_REG16664_S1 : DFF_X1 port map( D => n3533, CK => CLK, Q => n_3454, QN 
                           => n51684);
   clk_r_REG16662_S1 : DFF_X1 port map( D => n3534, CK => CLK, Q => n_3455, QN 
                           => n51683);
   clk_r_REG16660_S1 : DFF_X1 port map( D => n3535, CK => CLK, Q => n_3456, QN 
                           => n51682);
   clk_r_REG16658_S1 : DFF_X1 port map( D => n3536, CK => CLK, Q => n_3457, QN 
                           => n51681);
   clk_r_REG16369_S1 : DFF_X1 port map( D => n2576, CK => CLK, Q => n_3458, QN 
                           => n51680);
   clk_r_REG15858_S1 : DFF_X1 port map( D => n2672, CK => CLK, Q => n_3459, QN 
                           => n51679);
   clk_r_REG15986_S1 : DFF_X1 port map( D => n2736, CK => CLK, Q => n_3460, QN 
                           => n51678);
   clk_r_REG16367_S1 : DFF_X1 port map( D => n2577, CK => CLK, Q => n_3461, QN 
                           => n51677);
   clk_r_REG15856_S1 : DFF_X1 port map( D => n2673, CK => CLK, Q => n_3462, QN 
                           => n51676);
   clk_r_REG15794_S1 : DFF_X1 port map( D => n2640, CK => CLK, Q => n_3463, QN 
                           => n51675);
   clk_r_REG14807_S1 : DFF_X1 port map( D => n3312, CK => CLK, Q => n_3464, QN 
                           => n51674);
   clk_r_REG15792_S1 : DFF_X1 port map( D => n2641, CK => CLK, Q => n_3465, QN 
                           => n51673);
   clk_r_REG15790_S1 : DFF_X1 port map( D => n2642, CK => CLK, Q => n_3466, QN 
                           => n51672);
   clk_r_REG15788_S1 : DFF_X1 port map( D => n2643, CK => CLK, Q => n_3467, QN 
                           => n51671);
   clk_r_REG16255_S1 : DFF_X1 port map( D => n2858, CK => CLK, Q => n_3468, QN 
                           => n51670);
   clk_r_REG15164_S1 : DFF_X1 port map( D => n3148, CK => CLK, Q => n_3469, QN 
                           => n51669);
   clk_r_REG16305_S1 : DFF_X1 port map( D => n2544, CK => CLK, Q => n_3470, QN 
                           => n51668);
   clk_r_REG15416_S1 : DFF_X1 port map( D => n2894, CK => CLK, Q => n_3471, QN 
                           => n51667);
   clk_r_REG15984_S1 : DFF_X1 port map( D => n2737, CK => CLK, Q => n_3472, QN 
                           => n51666);
   clk_r_REG15982_S1 : DFF_X1 port map( D => n2738, CK => CLK, Q => n_3473, QN 
                           => n51665);
   clk_r_REG15980_S1 : DFF_X1 port map( D => n2739, CK => CLK, Q => n_3474, QN 
                           => n51664);
   clk_r_REG15854_S1 : DFF_X1 port map( D => n2674, CK => CLK, Q => n_3475, QN 
                           => n51663);
   clk_r_REG16050_S1 : DFF_X1 port map( D => n2768, CK => CLK, Q => n_3476, QN 
                           => n51662);
   clk_r_REG15852_S1 : DFF_X1 port map( D => n2675, CK => CLK, Q => n_3477, QN 
                           => n51661);
   clk_r_REG15942_S1 : DFF_X1 port map( D => n2704, CK => CLK, Q => n_3478, QN 
                           => n51660);
   clk_r_REG13817_S1 : DFF_X1 port map( D => n2949, CK => CLK, Q => n_3479, QN 
                           => n51659);
   clk_r_REG15730_S1 : DFF_X1 port map( D => n2608, CK => CLK, Q => n_3480, QN 
                           => n51658);
   clk_r_REG15728_S1 : DFF_X1 port map( D => n2609, CK => CLK, Q => n_3481, QN 
                           => n51657);
   clk_r_REG15414_S1 : DFF_X1 port map( D => n2895, CK => CLK, Q => n_3482, QN 
                           => n51656);
   clk_r_REG15940_S1 : DFF_X1 port map( D => n2705, CK => CLK, Q => n_3483, QN 
                           => n51655);
   clk_r_REG16048_S1 : DFF_X1 port map( D => n2769, CK => CLK, Q => n_3484, QN 
                           => n51654);
   clk_r_REG15850_S1 : DFF_X1 port map( D => n2676, CK => CLK, Q => n_3485, QN 
                           => n51653);
   clk_r_REG15978_S1 : DFF_X1 port map( D => n2740, CK => CLK, Q => n_3486, QN 
                           => n51652);
   clk_r_REG15786_S1 : DFF_X1 port map( D => n2644, CK => CLK, Q => n_3487, QN 
                           => n51651);
   clk_r_REG16365_S1 : DFF_X1 port map( D => n2578, CK => CLK, Q => n_3488, QN 
                           => n51650);
   clk_r_REG15938_S1 : DFF_X1 port map( D => n2706, CK => CLK, Q => n_3489, QN 
                           => n51649);
   clk_r_REG15726_S1 : DFF_X1 port map( D => n2610, CK => CLK, Q => n_3490, QN 
                           => n51648);
   clk_r_REG15784_S1 : DFF_X1 port map( D => n2645, CK => CLK, Q => n_3491, QN 
                           => n51647);
   clk_r_REG15976_S1 : DFF_X1 port map( D => n2741, CK => CLK, Q => n_3492, QN 
                           => n51646);
   clk_r_REG16303_S1 : DFF_X1 port map( D => n2545, CK => CLK, Q => n_3493, QN 
                           => n51645);
   clk_r_REG16363_S1 : DFF_X1 port map( D => n2579, CK => CLK, Q => n_3494, QN 
                           => n51644);
   clk_r_REG15782_S1 : DFF_X1 port map( D => n2646, CK => CLK, Q => n_3495, QN 
                           => n51643);
   clk_r_REG15848_S1 : DFF_X1 port map( D => n2677, CK => CLK, Q => n_3496, QN 
                           => n51642);
   clk_r_REG15846_S1 : DFF_X1 port map( D => n2678, CK => CLK, Q => n_3497, QN 
                           => n51641);
   clk_r_REG15780_S1 : DFF_X1 port map( D => n2647, CK => CLK, Q => n_3498, QN 
                           => n51640);
   clk_r_REG16361_S1 : DFF_X1 port map( D => n2580, CK => CLK, Q => n_3499, QN 
                           => n51639);
   clk_r_REG16125_S1 : DFF_X1 port map( D => n2795, CK => CLK, Q => n_3500, QN 
                           => n51638);
   clk_r_REG15974_S1 : DFF_X1 port map( D => n2742, CK => CLK, Q => n_3501, QN 
                           => n51637);
   clk_r_REG15972_S1 : DFF_X1 port map( D => n2743, CK => CLK, Q => n_3502, QN 
                           => n51636);
   clk_r_REG15844_S1 : DFF_X1 port map( D => n2679, CK => CLK, Q => n_3503, QN 
                           => n51635);
   clk_r_REG15778_S1 : DFF_X1 port map( D => n2648, CK => CLK, Q => n_3504, QN 
                           => n51634);
   clk_r_REG16359_S1 : DFF_X1 port map( D => n2581, CK => CLK, Q => n_3505, QN 
                           => n51633);
   clk_r_REG15162_S1 : DFF_X1 port map( D => n3149, CK => CLK, Q => n_3506, QN 
                           => n51632);
   clk_r_REG15970_S1 : DFF_X1 port map( D => n2744, CK => CLK, Q => n_3507, QN 
                           => n51631);
   clk_r_REG15842_S1 : DFF_X1 port map( D => n2680, CK => CLK, Q => n_3508, QN 
                           => n51630);
   clk_r_REG16357_S1 : DFF_X1 port map( D => n2582, CK => CLK, Q => n_3509, QN 
                           => n51629);
   clk_r_REG15776_S1 : DFF_X1 port map( D => n2649, CK => CLK, Q => n_3510, QN 
                           => n51628);
   clk_r_REG16301_S1 : DFF_X1 port map( D => n2546, CK => CLK, Q => n_3511, QN 
                           => n51627);
   clk_r_REG13659_S1 : DFF_X1 port map( D => n3237, CK => CLK, Q => n_3512, QN 
                           => n51626);
   clk_r_REG16046_S1 : DFF_X1 port map( D => n2770, CK => CLK, Q => n_3513, QN 
                           => n51625);
   clk_r_REG16355_S1 : DFF_X1 port map( D => n2583, CK => CLK, Q => n_3514, QN 
                           => n51624);
   clk_r_REG16123_S1 : DFF_X1 port map( D => n2796, CK => CLK, Q => n_3515, QN 
                           => n51623);
   clk_r_REG16044_S1 : DFF_X1 port map( D => n2771, CK => CLK, Q => n_3516, QN 
                           => n51622);
   clk_r_REG16253_S1 : DFF_X1 port map( D => n2859, CK => CLK, Q => n_3517, QN 
                           => n51621);
   clk_r_REG16042_S1 : DFF_X1 port map( D => n2772, CK => CLK, Q => n_3518, QN 
                           => n51620);
   clk_r_REG15672_S1 : DFF_X1 port map( D => n3022, CK => CLK, Q => n_3519, QN 
                           => n51619);
   clk_r_REG15968_S1 : DFF_X1 port map( D => n2745, CK => CLK, Q => n_3520, QN 
                           => n51618);
   clk_r_REG16299_S1 : DFF_X1 port map( D => n2547, CK => CLK, Q => n_3521, QN 
                           => n51617);
   clk_r_REG16576_S1 : DFF_X1 port map( D => n3209, CK => CLK, Q => n_3522, QN 
                           => n51616);
   clk_r_REG15412_S1 : DFF_X1 port map( D => n2896, CK => CLK, Q => n_3523, QN 
                           => n51615);
   clk_r_REG16353_S1 : DFF_X1 port map( D => n2584, CK => CLK, Q => n_3524, QN 
                           => n51614);
   clk_r_REG15840_S1 : DFF_X1 port map( D => n2681, CK => CLK, Q => n_3525, QN 
                           => n51613);
   clk_r_REG15936_S1 : DFF_X1 port map( D => n2707, CK => CLK, Q => n_3526, QN 
                           => n51612);
   clk_r_REG15460_S1 : DFF_X1 port map( D => n2925, CK => CLK, Q => n_3527, QN 
                           => n51611);
   clk_r_REG15934_S1 : DFF_X1 port map( D => n2708, CK => CLK, Q => n_3528, QN 
                           => n51610);
   clk_r_REG16040_S1 : DFF_X1 port map( D => n2773, CK => CLK, Q => n_3529, QN 
                           => n51609);
   clk_r_REG16574_S1 : DFF_X1 port map( D => n3210, CK => CLK, Q => n_3530, QN 
                           => n51608);
   clk_r_REG16251_S1 : DFF_X1 port map( D => n2860, CK => CLK, Q => n_3531, QN 
                           => n51607);
   clk_r_REG15724_S1 : DFF_X1 port map( D => n2611, CK => CLK, Q => n_3532, QN 
                           => n51606);
   clk_r_REG15966_S1 : DFF_X1 port map( D => n2746, CK => CLK, Q => n_3533, QN 
                           => n51605);
   clk_r_REG16297_S1 : DFF_X1 port map( D => n2548, CK => CLK, Q => n_3534, QN 
                           => n51604);
   clk_r_REG16038_S1 : DFF_X1 port map( D => n2774, CK => CLK, Q => n_3535, QN 
                           => n51603);
   clk_r_REG16249_S1 : DFF_X1 port map( D => n2861, CK => CLK, Q => n_3536, QN 
                           => n51602);
   clk_r_REG16572_S1 : DFF_X1 port map( D => n3211, CK => CLK, Q => n_3537, QN 
                           => n51601);
   clk_r_REG16036_S1 : DFF_X1 port map( D => n2775, CK => CLK, Q => n_3538, QN 
                           => n51600);
   clk_r_REG15670_S1 : DFF_X1 port map( D => n3023, CK => CLK, Q => n_3539, QN 
                           => n51599);
   clk_r_REG15932_S1 : DFF_X1 port map( D => n2709, CK => CLK, Q => n_3540, QN 
                           => n51598);
   clk_r_REG15774_S1 : DFF_X1 port map( D => n2650, CK => CLK, Q => n_3541, QN 
                           => n51597);
   clk_r_REG16295_S1 : DFF_X1 port map( D => n2549, CK => CLK, Q => n_3542, QN 
                           => n51596);
   clk_r_REG16034_S1 : DFF_X1 port map( D => n2776, CK => CLK, Q => n_3543, QN 
                           => n51595);
   clk_r_REG15722_S1 : DFF_X1 port map( D => n2612, CK => CLK, Q => n_3544, QN 
                           => n51594);
   clk_r_REG16032_S1 : DFF_X1 port map( D => n2777, CK => CLK, Q => n_3545, QN 
                           => n51593);
   clk_r_REG15295_S1 : DFF_X1 port map( D => n3244, CK => CLK, Q => n_3546, QN 
                           => n51592);
   clk_r_REG15930_S1 : DFF_X1 port map( D => n2710, CK => CLK, Q => n_3547, QN 
                           => n51591);
   clk_r_REG15606_S1 : DFF_X1 port map( D => n2991, CK => CLK, Q => n_3548, QN 
                           => n51590);
   clk_r_REG15928_S1 : DFF_X1 port map( D => n2711, CK => CLK, Q => n_3549, QN 
                           => n51589);
   clk_r_REG15720_S1 : DFF_X1 port map( D => n2613, CK => CLK, Q => n_3550, QN 
                           => n51588);
   clk_r_REG15718_S1 : DFF_X1 port map( D => n2614, CK => CLK, Q => n_3551, QN 
                           => n51587);
   clk_r_REG15544_S1 : DFF_X1 port map( D => n2958, CK => CLK, Q => n_3552, QN 
                           => n51586);
   clk_r_REG15604_S1 : DFF_X1 port map( D => n2992, CK => CLK, Q => n_3553, QN 
                           => n51585);
   clk_r_REG16030_S1 : DFF_X1 port map( D => n2778, CK => CLK, Q => n_3554, QN 
                           => n51584);
   clk_r_REG16293_S1 : DFF_X1 port map( D => n2550, CK => CLK, Q => n_3555, QN 
                           => n51583);
   clk_r_REG16570_S1 : DFF_X1 port map( D => n3212, CK => CLK, Q => n_3556, QN 
                           => n51582);
   clk_r_REG16568_S1 : DFF_X1 port map( D => n3213, CK => CLK, Q => n_3557, QN 
                           => n51581);
   clk_r_REG16291_S1 : DFF_X1 port map( D => n2551, CK => CLK, Q => n_3558, QN 
                           => n51580);
   clk_r_REG16566_S1 : DFF_X1 port map( D => n3214, CK => CLK, Q => n_3559, QN 
                           => n51579);
   clk_r_REG16564_S1 : DFF_X1 port map( D => n3215, CK => CLK, Q => n_3560, QN 
                           => n51578);
   clk_r_REG15716_S1 : DFF_X1 port map( D => n2615, CK => CLK, Q => n_3561, QN 
                           => n51577);
   clk_r_REG15964_S1 : DFF_X1 port map( D => n2747, CK => CLK, Q => n_3562, QN 
                           => n51576);
   clk_r_REG16247_S1 : DFF_X1 port map( D => n2862, CK => CLK, Q => n_3563, QN 
                           => n51575);
   clk_r_REG15962_S1 : DFF_X1 port map( D => n2748, CK => CLK, Q => n_3564, QN 
                           => n51574);
   clk_r_REG15960_S1 : DFF_X1 port map( D => n2749, CK => CLK, Q => n_3565, QN 
                           => n51573);
   clk_r_REG15926_S1 : DFF_X1 port map( D => n2712, CK => CLK, Q => n_3566, QN 
                           => n51572);
   clk_r_REG15772_S1 : DFF_X1 port map( D => n2651, CK => CLK, Q => n_3567, QN 
                           => n51571);
   clk_r_REG16289_S1 : DFF_X1 port map( D => n2552, CK => CLK, Q => n_3568, QN 
                           => n51570);
   clk_r_REG15958_S1 : DFF_X1 port map( D => n2750, CK => CLK, Q => n_3569, QN 
                           => n51569);
   clk_r_REG15714_S1 : DFF_X1 port map( D => n2616, CK => CLK, Q => n_3570, QN 
                           => n51568);
   clk_r_REG15924_S1 : DFF_X1 port map( D => n2713, CK => CLK, Q => n_3571, QN 
                           => n51567);
   clk_r_REG16287_S1 : DFF_X1 port map( D => n2553, CK => CLK, Q => n_3572, QN 
                           => n51566);
   clk_r_REG16285_S1 : DFF_X1 port map( D => n2554, CK => CLK, Q => n_3573, QN 
                           => n51565);
   clk_r_REG16351_S1 : DFF_X1 port map( D => n2585, CK => CLK, Q => n_3574, QN 
                           => n51564);
   clk_r_REG15712_S1 : DFF_X1 port map( D => n2617, CK => CLK, Q => n_3575, QN 
                           => n51563);
   clk_r_REG16562_S1 : DFF_X1 port map( D => n3216, CK => CLK, Q => n_3576, QN 
                           => n51562);
   clk_r_REG15770_S1 : DFF_X1 port map( D => n2652, CK => CLK, Q => n_3577, QN 
                           => n51561);
   clk_r_REG15458_S1 : DFF_X1 port map( D => n2924, CK => CLK, Q => n_3578, QN 
                           => n51560);
   clk_r_REG15838_S1 : DFF_X1 port map( D => n2682, CK => CLK, Q => n_3579, QN 
                           => n51559);
   clk_r_REG16028_S1 : DFF_X1 port map( D => n2779, CK => CLK, Q => n_3580, QN 
                           => n51558);
   clk_r_REG16283_S1 : DFF_X1 port map( D => n2555, CK => CLK, Q => n_3581, QN 
                           => n51557);
   clk_r_REG16281_S1 : DFF_X1 port map( D => n2556, CK => CLK, Q => n_3582, QN 
                           => n51556);
   clk_r_REG16279_S1 : DFF_X1 port map( D => n2557, CK => CLK, Q => n_3583, QN 
                           => n51555);
   clk_r_REG16026_S1 : DFF_X1 port map( D => n2780, CK => CLK, Q => n_3584, QN 
                           => n51554);
   clk_r_REG15456_S1 : DFF_X1 port map( D => n2923, CK => CLK, Q => n_3585, QN 
                           => n51553);
   clk_r_REG15293_S1 : DFF_X1 port map( D => n3245, CK => CLK, Q => n_3586, QN 
                           => n51552);
   clk_r_REG15922_S1 : DFF_X1 port map( D => n2714, CK => CLK, Q => n_3587, QN 
                           => n51551);
   clk_r_REG15768_S1 : DFF_X1 port map( D => n2653, CK => CLK, Q => n_3588, QN 
                           => n51550);
   clk_r_REG15766_S1 : DFF_X1 port map( D => n2654, CK => CLK, Q => n_3589, QN 
                           => n51549);
   clk_r_REG16277_S1 : DFF_X1 port map( D => n2558, CK => CLK, Q => n_3590, QN 
                           => n51548);
   clk_r_REG15920_S1 : DFF_X1 port map( D => n2715, CK => CLK, Q => n_3591, QN 
                           => n51547);
   clk_r_REG15918_S1 : DFF_X1 port map( D => n2716, CK => CLK, Q => n_3592, QN 
                           => n51546);
   clk_r_REG15291_S1 : DFF_X1 port map( D => n3246, CK => CLK, Q => n_3593, QN 
                           => n51545);
   clk_r_REG15542_S1 : DFF_X1 port map( D => n2959, CK => CLK, Q => n_3594, QN 
                           => n51544);
   clk_r_REG16024_S1 : DFF_X1 port map( D => n2781, CK => CLK, Q => n_3595, QN 
                           => n51543);
   clk_r_REG15916_S1 : DFF_X1 port map( D => n2717, CK => CLK, Q => n_3596, QN 
                           => n51542);
   clk_r_REG15090_S1 : DFF_X1 port map( D => n3055, CK => CLK, Q => n_3597, QN 
                           => n51541);
   clk_r_REG16349_S1 : DFF_X1 port map( D => n2586, CK => CLK, Q => n_3598, QN 
                           => n51540);
   clk_r_REG15289_S1 : DFF_X1 port map( D => n3247, CK => CLK, Q => n_3599, QN 
                           => n51539);
   clk_r_REG16347_S1 : DFF_X1 port map( D => n2587, CK => CLK, Q => n_3600, QN 
                           => n51538);
   clk_r_REG15454_S1 : DFF_X1 port map( D => n2922, CK => CLK, Q => n_3601, QN 
                           => n51537);
   clk_r_REG15836_S1 : DFF_X1 port map( D => n2683, CK => CLK, Q => n_3602, QN 
                           => n51536);
   clk_r_REG16345_S1 : DFF_X1 port map( D => n2588, CK => CLK, Q => n_3603, QN 
                           => n51535);
   clk_r_REG15710_S1 : DFF_X1 port map( D => n2618, CK => CLK, Q => n_3604, QN 
                           => n51534);
   clk_r_REG15287_S1 : DFF_X1 port map( D => n3248, CK => CLK, Q => n_3605, QN 
                           => n51533);
   clk_r_REG15088_S1 : DFF_X1 port map( D => n3056, CK => CLK, Q => n_3606, QN 
                           => n51532);
   clk_r_REG15914_S1 : DFF_X1 port map( D => n2718, CK => CLK, Q => n_3607, QN 
                           => n51531);
   clk_r_REG16022_S1 : DFF_X1 port map( D => n2782, CK => CLK, Q => n_3608, QN 
                           => n51530);
   clk_r_REG15834_S1 : DFF_X1 port map( D => n2684, CK => CLK, Q => n_3609, QN 
                           => n51529);
   clk_r_REG15832_S1 : DFF_X1 port map( D => n2685, CK => CLK, Q => n_3610, QN 
                           => n51528);
   clk_r_REG15668_S1 : DFF_X1 port map( D => n3024, CK => CLK, Q => n_3611, QN 
                           => n51527);
   clk_r_REG16245_S1 : DFF_X1 port map( D => n2863, CK => CLK, Q => n_3612, QN 
                           => n51526);
   clk_r_REG15830_S1 : DFF_X1 port map( D => n2686, CK => CLK, Q => n_3613, QN 
                           => n51525);
   clk_r_REG15708_S1 : DFF_X1 port map( D => n2619, CK => CLK, Q => n_3614, QN 
                           => n51524);
   clk_r_REG15706_S1 : DFF_X1 port map( D => n2620, CK => CLK, Q => n_3615, QN 
                           => n51523);
   clk_r_REG16343_S1 : DFF_X1 port map( D => n2589, CK => CLK, Q => n_3616, QN 
                           => n51522);
   clk_r_REG16121_S1 : DFF_X1 port map( D => n2797, CK => CLK, Q => n_3617, QN 
                           => n51521);
   clk_r_REG15540_S1 : DFF_X1 port map( D => n2960, CK => CLK, Q => n_3618, QN 
                           => n51520);
   clk_r_REG16341_S1 : DFF_X1 port map( D => n2590, CK => CLK, Q => n_3619, QN 
                           => n51519);
   clk_r_REG15704_S1 : DFF_X1 port map( D => n2621, CK => CLK, Q => n_3620, QN 
                           => n51518);
   clk_r_REG15702_S1 : DFF_X1 port map( D => n2622, CK => CLK, Q => n_3621, QN 
                           => n51517);
   clk_r_REG15452_S1 : DFF_X1 port map( D => n2921, CK => CLK, Q => n_3622, QN 
                           => n51516);
   clk_r_REG16020_S1 : DFF_X1 port map( D => n2783, CK => CLK, Q => n_3623, QN 
                           => n51515);
   clk_r_REG15450_S1 : DFF_X1 port map( D => n2920, CK => CLK, Q => n_3624, QN 
                           => n51514);
   clk_r_REG15160_S1 : DFF_X1 port map( D => n3150, CK => CLK, Q => n_3625, QN 
                           => n51513);
   clk_r_REG15448_S1 : DFF_X1 port map( D => n2919, CK => CLK, Q => n_3626, QN 
                           => n51512);
   clk_r_REG16275_S1 : DFF_X1 port map( D => n2559, CK => CLK, Q => n_3627, QN 
                           => n51511);
   clk_r_REG16498_S1 : DFF_X1 port map( D => n3120, CK => CLK, Q => n_3628, QN 
                           => n51510);
   clk_r_REG16243_S1 : DFF_X1 port map( D => n2864, CK => CLK, Q => n_3629, QN 
                           => n51509);
   clk_r_REG15446_S1 : DFF_X1 port map( D => n2918, CK => CLK, Q => n_3630, QN 
                           => n51508);
   clk_r_REG16070_S1 : DFF_X1 port map( D => n2758, CK => CLK, Q => n_3631, QN 
                           => n51507);
   clk_r_REG15814_S1 : DFF_X1 port map( D => n2630, CK => CLK, Q => n_3632, QN 
                           => n51506);
   clk_r_REG15764_S1 : DFF_X1 port map( D => n2655, CK => CLK, Q => n_3633, QN 
                           => n51505);
   clk_r_REG16068_S1 : DFF_X1 port map( D => n2759, CK => CLK, Q => n_3634, QN 
                           => n51504);
   clk_r_REG15762_S1 : DFF_X1 port map( D => n2656, CK => CLK, Q => n_3635, QN 
                           => n51503);
   clk_r_REG15956_S1 : DFF_X1 port map( D => n2751, CK => CLK, Q => n_3636, QN 
                           => n51502);
   clk_r_REG16018_S1 : DFF_X1 port map( D => n2784, CK => CLK, Q => n_3637, QN 
                           => n51501);
   clk_r_REG16183_S1 : DFF_X1 port map( D => n2830, CK => CLK, Q => n_3638, QN 
                           => n51500);
   clk_r_REG16016_S1 : DFF_X1 port map( D => n2785, CK => CLK, Q => n_3639, QN 
                           => n51499);
   clk_r_REG16119_S1 : DFF_X1 port map( D => n2798, CK => CLK, Q => n_3640, QN 
                           => n51498);
   clk_r_REG15700_S1 : DFF_X1 port map( D => n2623, CK => CLK, Q => n_3641, QN 
                           => n51497);
   clk_r_REG16339_S1 : DFF_X1 port map( D => n2591, CK => CLK, Q => n_3642, QN 
                           => n51496);
   clk_r_REG16181_S1 : DFF_X1 port map( D => n2831, CK => CLK, Q => n_3643, QN 
                           => n51495);
   clk_r_REG15828_S1 : DFF_X1 port map( D => n2687, CK => CLK, Q => n_3644, QN 
                           => n51494);
   clk_r_REG16273_S1 : DFF_X1 port map( D => n2560, CK => CLK, Q => n_3645, QN 
                           => n51493);
   clk_r_REG15750_S1 : DFF_X1 port map( D => n2598, CK => CLK, Q => n_3646, QN 
                           => n51492);
   clk_r_REG15912_S1 : DFF_X1 port map( D => n2719, CK => CLK, Q => n_3647, QN 
                           => n51491);
   clk_r_REG15748_S1 : DFF_X1 port map( D => n2599, CK => CLK, Q => n_3648, QN 
                           => n51490);
   clk_r_REG15698_S1 : DFF_X1 port map( D => n2624, CK => CLK, Q => n_3649, QN 
                           => n51489);
   clk_r_REG15910_S1 : DFF_X1 port map( D => n2720, CK => CLK, Q => n_3650, QN 
                           => n51488);
   clk_r_REG15954_S1 : DFF_X1 port map( D => n2752, CK => CLK, Q => n_3651, QN 
                           => n51487);
   clk_r_REG15696_S1 : DFF_X1 port map( D => n2625, CK => CLK, Q => n_3652, QN 
                           => n51486);
   clk_r_REG15908_S1 : DFF_X1 port map( D => n2703, CK => CLK, Q => n_3653, QN 
                           => n51485);
   clk_r_REG16014_S1 : DFF_X1 port map( D => n2786, CK => CLK, Q => n_3654, QN 
                           => n51484);
   clk_r_REG16435_S1 : DFF_X1 port map( D => n3087, CK => CLK, Q => n_3655, QN 
                           => n51483);
   clk_r_REG16433_S1 : DFF_X1 port map( D => n3088, CK => CLK, Q => n_3656, QN 
                           => n51482);
   clk_r_REG16117_S1 : DFF_X1 port map( D => n2799, CK => CLK, Q => n_3657, QN 
                           => n51481);
   clk_r_REG16115_S1 : DFF_X1 port map( D => n2800, CK => CLK, Q => n_3658, QN 
                           => n51480);
   clk_r_REG15826_S1 : DFF_X1 port map( D => n2688, CK => CLK, Q => n_3659, QN 
                           => n51479);
   clk_r_REG16325_S1 : DFF_X1 port map( D => n2534, CK => CLK, Q => n_3660, QN 
                           => n51478);
   clk_r_REG16006_S1 : DFF_X1 port map( D => n2726, CK => CLK, Q => n_3661, QN 
                           => n51477);
   clk_r_REG15158_S1 : DFF_X1 port map( D => n3151, CK => CLK, Q => n_3662, QN 
                           => n51476);
   clk_r_REG15906_S1 : DFF_X1 port map( D => n2702, CK => CLK, Q => n_3663, QN 
                           => n51475);
   clk_r_REG15878_S1 : DFF_X1 port map( D => n2662, CK => CLK, Q => n_3664, QN 
                           => n51474);
   clk_r_REG16012_S1 : DFF_X1 port map( D => n2787, CK => CLK, Q => n_3665, QN 
                           => n51473);
   clk_r_REG15694_S1 : DFF_X1 port map( D => n2626, CK => CLK, Q => n_3666, QN 
                           => n51472);
   clk_r_REG16004_S1 : DFF_X1 port map( D => n2727, CK => CLK, Q => n_3667, QN 
                           => n51471);
   clk_r_REG16323_S1 : DFF_X1 port map( D => n2535, CK => CLK, Q => n_3668, QN 
                           => n51470);
   clk_r_REG15876_S1 : DFF_X1 port map( D => n2663, CK => CLK, Q => n_3669, QN 
                           => n51469);
   clk_r_REG15952_S1 : DFF_X1 port map( D => n2753, CK => CLK, Q => n_3670, QN 
                           => n51468);
   clk_r_REG15888_S1 : DFF_X1 port map( D => n2721, CK => CLK, Q => n_3671, QN 
                           => n51467);
   clk_r_REG15886_S1 : DFF_X1 port map( D => n2722, CK => CLK, Q => n_3672, QN 
                           => n51466);
   clk_r_REG16271_S1 : DFF_X1 port map( D => n2561, CK => CLK, Q => n_3673, QN 
                           => n51465);
   clk_r_REG16269_S1 : DFF_X1 port map( D => n2562, CK => CLK, Q => n_3674, QN 
                           => n51464);
   clk_r_REG16337_S1 : DFF_X1 port map( D => n2592, CK => CLK, Q => n_3675, QN 
                           => n51463);
   clk_r_REG16389_S1 : DFF_X1 port map( D => n2566, CK => CLK, Q => n_3676, QN 
                           => n51462);
   clk_r_REG16387_S1 : DFF_X1 port map( D => n2567, CK => CLK, Q => n_3677, QN 
                           => n51461);
   clk_r_REG15692_S1 : DFF_X1 port map( D => n2627, CK => CLK, Q => n_3678, QN 
                           => n51460);
   clk_r_REG15690_S1 : DFF_X1 port map( D => n2628, CK => CLK, Q => n_3679, QN 
                           => n51459);
   clk_r_REG15884_S1 : DFF_X1 port map( D => n2723, CK => CLK, Q => n_3680, QN 
                           => n51458);
   clk_r_REG15882_S1 : DFF_X1 port map( D => n2724, CK => CLK, Q => n_3681, QN 
                           => n51457);
   clk_r_REG15950_S1 : DFF_X1 port map( D => n2754, CK => CLK, Q => n_3682, QN 
                           => n51456);
   clk_r_REG16267_S1 : DFF_X1 port map( D => n2563, CK => CLK, Q => n_3683, QN 
                           => n51455);
   clk_r_REG15812_S1 : DFF_X1 port map( D => n2631, CK => CLK, Q => n_3684, QN 
                           => n51454);
   clk_r_REG15824_S1 : DFF_X1 port map( D => n2689, CK => CLK, Q => n_3685, QN 
                           => n51453);
   clk_r_REG16265_S1 : DFF_X1 port map( D => n2564, CK => CLK, Q => n_3686, QN 
                           => n51452);
   clk_r_REG15822_S1 : DFF_X1 port map( D => n2690, CK => CLK, Q => n_3687, QN 
                           => n51451);
   clk_r_REG15760_S1 : DFF_X1 port map( D => n2657, CK => CLK, Q => n_3688, QN 
                           => n51450);
   clk_r_REG15156_S1 : DFF_X1 port map( D => n3152, CK => CLK, Q => n_3689, QN 
                           => n51449);
   clk_r_REG15758_S1 : DFF_X1 port map( D => n2658, CK => CLK, Q => n_3690, QN 
                           => n51448);
   clk_r_REG15756_S1 : DFF_X1 port map( D => n2659, CK => CLK, Q => n_3691, QN 
                           => n51447);
   clk_r_REG16335_S1 : DFF_X1 port map( D => n2593, CK => CLK, Q => n_3692, QN 
                           => n51446);
   clk_r_REG16179_S1 : DFF_X1 port map( D => n2832, CK => CLK, Q => n_3693, QN 
                           => n51445);
   clk_r_REG16333_S1 : DFF_X1 port map( D => n2594, CK => CLK, Q => n_3694, QN 
                           => n51444);
   clk_r_REG16010_S1 : DFF_X1 port map( D => n2788, CK => CLK, Q => n_3695, QN 
                           => n51443);
   clk_r_REG15754_S1 : DFF_X1 port map( D => n2660, CK => CLK, Q => n_3696, QN 
                           => n51442);
   clk_r_REG16331_S1 : DFF_X1 port map( D => n2595, CK => CLK, Q => n_3697, QN 
                           => n51441);
   clk_r_REG15948_S1 : DFF_X1 port map( D => n2755, CK => CLK, Q => n_3698, QN 
                           => n51440);
   clk_r_REG15820_S1 : DFF_X1 port map( D => n2691, CK => CLK, Q => n_3699, QN 
                           => n51439);
   clk_r_REG15818_S1 : DFF_X1 port map( D => n2692, CK => CLK, Q => n_3700, QN 
                           => n51438);
   clk_r_REG15946_S1 : DFF_X1 port map( D => n2756, CK => CLK, Q => n_3701, QN 
                           => n51437);
   clk_r_REG16329_S1 : DFF_X1 port map( D => n2596, CK => CLK, Q => n_3702, QN 
                           => n51436);
   clk_r_REG13741_S1 : DFF_X1 port map( D => n2789, CK => CLK, Q => n_3703, QN 
                           => n51435);
   clk_r_REG13778_S1 : DFF_X1 port map( D => n2629, CK => CLK, Q => n_3704, QN 
                           => n51434);
   clk_r_REG15746_S1 : DFF_X1 port map( D => n2600, CK => CLK, Q => n_3705, QN 
                           => n51433);
   clk_r_REG15744_S1 : DFF_X1 port map( D => n2601, CK => CLK, Q => n_3706, QN 
                           => n51432);
   clk_r_REG15742_S1 : DFF_X1 port map( D => n2602, CK => CLK, Q => n_3707, QN 
                           => n51431);
   clk_r_REG13757_S1 : DFF_X1 port map( D => n2725, CK => CLK, Q => n_3708, QN 
                           => n51430);
   clk_r_REG15904_S1 : DFF_X1 port map( D => n2701, CK => CLK, Q => n_3709, QN 
                           => n51429);
   clk_r_REG13771_S1 : DFF_X1 port map( D => n2661, CK => CLK, Q => n_3710, QN 
                           => n51428);
   clk_r_REG15902_S1 : DFF_X1 port map( D => n2700, CK => CLK, Q => n_3711, QN 
                           => n51427);
   clk_r_REG15810_S1 : DFF_X1 port map( D => n2632, CK => CLK, Q => n_3712, QN 
                           => n51426);
   clk_r_REG15900_S1 : DFF_X1 port map( D => n2699, CK => CLK, Q => n_3713, QN 
                           => n51425);
   clk_r_REG15740_S1 : DFF_X1 port map( D => n2603, CK => CLK, Q => n_3714, QN 
                           => n51424);
   clk_r_REG13764_S1 : DFF_X1 port map( D => n2693, CK => CLK, Q => n_3715, QN 
                           => n51423);
   clk_r_REG15874_S1 : DFF_X1 port map( D => n2664, CK => CLK, Q => n_3716, QN 
                           => n51422);
   clk_r_REG13701_S1 : DFF_X1 port map( D => n2597, CK => CLK, Q => n_3717, QN 
                           => n51421);
   clk_r_REG16385_S1 : DFF_X1 port map( D => n2568, CK => CLK, Q => n_3718, QN 
                           => n51420);
   clk_r_REG15808_S1 : DFF_X1 port map( D => n2633, CK => CLK, Q => n_3719, QN 
                           => n51419);
   clk_r_REG15806_S1 : DFF_X1 port map( D => n2634, CK => CLK, Q => n_3720, QN 
                           => n51418);
   clk_r_REG15872_S1 : DFF_X1 port map( D => n2665, CK => CLK, Q => n_3721, QN 
                           => n51417);
   clk_r_REG15870_S1 : DFF_X1 port map( D => n2666, CK => CLK, Q => n_3722, QN 
                           => n51416);
   clk_r_REG15804_S1 : DFF_X1 port map( D => n2635, CK => CLK, Q => n_3723, QN 
                           => n51415);
   clk_r_REG16383_S1 : DFF_X1 port map( D => n2569, CK => CLK, Q => n_3724, QN 
                           => n51414);
   clk_r_REG16381_S1 : DFF_X1 port map( D => n2570, CK => CLK, Q => n_3725, QN 
                           => n51413);
   clk_r_REG13750_S1 : DFF_X1 port map( D => n2757, CK => CLK, Q => n_3726, QN 
                           => n51412);
   clk_r_REG16379_S1 : DFF_X1 port map( D => n2571, CK => CLK, Q => n_3727, QN 
                           => n51411);
   clk_r_REG15868_S1 : DFF_X1 port map( D => n2667, CK => CLK, Q => n_3728, QN 
                           => n51410);
   clk_r_REG13708_S1 : DFF_X1 port map( D => n2565, CK => CLK, Q => n_3729, QN 
                           => n51409);
   clk_r_REG16066_S1 : DFF_X1 port map( D => n2760, CK => CLK, Q => n_3730, QN 
                           => n51408);
   clk_r_REG16377_S1 : DFF_X1 port map( D => n2572, CK => CLK, Q => n_3731, QN 
                           => n51407);
   clk_r_REG15738_S1 : DFF_X1 port map( D => n2604, CK => CLK, Q => n_3732, QN 
                           => n51406);
   clk_r_REG16321_S1 : DFF_X1 port map( D => n2536, CK => CLK, Q => n_3733, QN 
                           => n51405);
   clk_r_REG15802_S1 : DFF_X1 port map( D => n2636, CK => CLK, Q => n_3734, QN 
                           => n51404);
   clk_r_REG15898_S1 : DFF_X1 port map( D => n2698, CK => CLK, Q => n_3735, QN 
                           => n51403);
   clk_r_REG15866_S1 : DFF_X1 port map( D => n2668, CK => CLK, Q => n_3736, QN 
                           => n51402);
   clk_r_REG15896_S1 : DFF_X1 port map( D => n2697, CK => CLK, Q => n_3737, QN 
                           => n51401);
   clk_r_REG15736_S1 : DFF_X1 port map( D => n2605, CK => CLK, Q => n_3738, QN 
                           => n51400);
   clk_r_REG15894_S1 : DFF_X1 port map( D => n2696, CK => CLK, Q => n_3739, QN 
                           => n51399);
   clk_r_REG16002_S1 : DFF_X1 port map( D => n2728, CK => CLK, Q => n_3740, QN 
                           => n51398);
   clk_r_REG16000_S1 : DFF_X1 port map( D => n2729, CK => CLK, Q => n_3741, QN 
                           => n51397);
   clk_r_REG16064_S1 : DFF_X1 port map( D => n2761, CK => CLK, Q => n_3742, QN 
                           => n51396);
   clk_r_REG16319_S1 : DFF_X1 port map( D => n2537, CK => CLK, Q => n_3743, QN 
                           => n51395);
   clk_r_REG16317_S1 : DFF_X1 port map( D => n2538, CK => CLK, Q => n_3744, QN 
                           => n51394);
   clk_r_REG15998_S1 : DFF_X1 port map( D => n2730, CK => CLK, Q => n_3745, QN 
                           => n51393);
   clk_r_REG15734_S1 : DFF_X1 port map( D => n2606, CK => CLK, Q => n_3746, QN 
                           => n51392);
   clk_r_REG16062_S1 : DFF_X1 port map( D => n2762, CK => CLK, Q => n_3747, QN 
                           => n51391);
   clk_r_REG16315_S1 : DFF_X1 port map( D => n2539, CK => CLK, Q => n_3748, QN 
                           => n51390);
   clk_r_REG16313_S1 : DFF_X1 port map( D => n2540, CK => CLK, Q => n_3749, QN 
                           => n51389);
   clk_r_REG15892_S1 : DFF_X1 port map( D => n2695, CK => CLK, Q => n_3750, QN 
                           => n51388);
   clk_r_REG16311_S1 : DFF_X1 port map( D => n2541, CK => CLK, Q => n_3751, QN 
                           => n51387);
   clk_r_REG15996_S1 : DFF_X1 port map( D => n2731, CK => CLK, Q => n_3752, QN 
                           => n51386);
   clk_r_REG15864_S1 : DFF_X1 port map( D => n2669, CK => CLK, Q => n_3753, QN 
                           => n51385);
   clk_r_REG16060_S1 : DFF_X1 port map( D => n2763, CK => CLK, Q => n_3754, QN 
                           => n51384);
   clk_r_REG15890_S1 : DFF_X1 port map( D => n2694, CK => CLK, Q => n_3755, QN 
                           => n51383);
   clk_r_REG16375_S1 : DFF_X1 port map( D => n2573, CK => CLK, Q => n_3756, QN 
                           => n51382);
   clk_r_REG16373_S1 : DFF_X1 port map( D => n2574, CK => CLK, Q => n_3757, QN 
                           => n51381);
   clk_r_REG16058_S1 : DFF_X1 port map( D => n2764, CK => CLK, Q => n_3758, QN 
                           => n51380);
   clk_r_REG15800_S1 : DFF_X1 port map( D => n2637, CK => CLK, Q => n_3759, QN 
                           => n51379);
   clk_r_REG16056_S1 : DFF_X1 port map( D => n2765, CK => CLK, Q => n_3760, QN 
                           => n51378);
   clk_r_REG15862_S1 : DFF_X1 port map( D => n2670, CK => CLK, Q => n_3761, QN 
                           => n51377);
   clk_r_REG15994_S1 : DFF_X1 port map( D => n2732, CK => CLK, Q => n_3762, QN 
                           => n51376);
   clk_r_REG15992_S1 : DFF_X1 port map( D => n2733, CK => CLK, Q => n_3763, QN 
                           => n51375);
   clk_r_REG15990_S1 : DFF_X1 port map( D => n2734, CK => CLK, Q => n_3764, QN 
                           => n51374);
   clk_r_REG15798_S1 : DFF_X1 port map( D => n2638, CK => CLK, Q => n_3765, QN 
                           => n51373);
   clk_r_REG16371_S1 : DFF_X1 port map( D => n2575, CK => CLK, Q => n_3766, QN 
                           => n51372);
   clk_r_REG16309_S1 : DFF_X1 port map( D => n2542, CK => CLK, Q => n_3767, QN 
                           => n51371);
   clk_r_REG16307_S1 : DFF_X1 port map( D => n2543, CK => CLK, Q => n_3768, QN 
                           => n51370);
   clk_r_REG16054_S1 : DFF_X1 port map( D => n2766, CK => CLK, Q => n_3769, QN 
                           => n51369);
   clk_r_REG15796_S1 : DFF_X1 port map( D => n2639, CK => CLK, Q => n_3770, QN 
                           => n51368);
   clk_r_REG16052_S1 : DFF_X1 port map( D => n2767, CK => CLK, Q => n_3771, QN 
                           => n51367);
   clk_r_REG15732_S1 : DFF_X1 port map( D => n2607, CK => CLK, Q => n_3772, QN 
                           => n51366);
   clk_r_REG15860_S1 : DFF_X1 port map( D => n2671, CK => CLK, Q => n_3773, QN 
                           => n51365);
   clk_r_REG15988_S1 : DFF_X1 port map( D => n2735, CK => CLK, Q => n_3774, QN 
                           => n51364);
   clk_r_REG16942_S7 : DFFR_X1 port map( D => n3570, CK => CLK, RN => RESET_BAR
                           , Q => n53566, QN => n_3775);
   clk_r_REG16939_S7 : DFFR_X1 port map( D => n3569, CK => CLK, RN => RESET_BAR
                           , Q => n53579, QN => n_3776);
   clk_r_REG16843_S7 : DFFR_X1 port map( D => n3566, CK => CLK, RN => RESET_BAR
                           , Q => n53547, QN => n_3777);
   clk_r_REG16923_S7 : DFFR_X1 port map( D => n49090, CK => CLK, RN => 
                           RESET_BAR, Q => n52427, QN => n_3778);
   clk_r_REG16901_S7 : DFFR_X1 port map( D => n49088, CK => CLK, RN => 
                           RESET_BAR, Q => n52425, QN => n_3779);
   clk_r_REG16851_S7 : DFFS_X1 port map( D => n3564, CK => CLK, SN => RESET_BAR
                           , Q => n_3780, QN => n52401);
   clk_r_REG16879_S7 : DFFS_X1 port map( D => n3563, CK => CLK, SN => RESET_BAR
                           , Q => n_3781, QN => n52482);
   clk_r_REG16872_S7 : DFFS_X1 port map( D => n3561, CK => CLK, SN => RESET_BAR
                           , Q => n_3782, QN => n52481);
   clk_r_REG16844_S7 : DFFS_X1 port map( D => n3565, CK => CLK, SN => RESET_BAR
                           , Q => n_3783, QN => n52479);
   clk_r_REG16886_S7 : DFFR_X1 port map( D => n3562, CK => CLK, RN => RESET_BAR
                           , Q => n_3784, QN => n52402);
   clk_r_REG16952_S7 : DFFS_X1 port map( D => n3572, CK => CLK, SN => RESET_BAR
                           , Q => n_3785, QN => n52400);
   clk_r_REG16858_S7 : DFFS_X1 port map( D => n3559, CK => CLK, SN => RESET_BAR
                           , Q => n_3786, QN => n52480);
   clk_r_REG16703_S5 : DFFS_X2 port map( D => n40605, CK => CLK, SN => 
                           RESET_BAR, Q => n52436, QN => n_3787);
   clk_r_REG16708_S5 : DFFS_X2 port map( D => n40610, CK => CLK, SN => 
                           RESET_BAR, Q => n52441, QN => n_3788);
   clk_r_REG16709_S5 : DFFS_X2 port map( D => n40611, CK => CLK, SN => 
                           RESET_BAR, Q => n52442, QN => n_3789);
   clk_r_REG16718_S5 : DFFS_X2 port map( D => n40612, CK => CLK, SN => 
                           RESET_BAR, Q => n52443, QN => n_3790);
   clk_r_REG16719_S5 : DFFS_X2 port map( D => n40613, CK => CLK, SN => 
                           RESET_BAR, Q => n52444, QN => n_3791);
   clk_r_REG16720_S5 : DFFS_X2 port map( D => n40614, CK => CLK, SN => 
                           RESET_BAR, Q => n52445, QN => n_3792);
   clk_r_REG16721_S5 : DFFS_X2 port map( D => n40615, CK => CLK, SN => 
                           RESET_BAR, Q => n52446, QN => n_3793);
   clk_r_REG16722_S5 : DFFS_X2 port map( D => n40616, CK => CLK, SN => 
                           RESET_BAR, Q => n52447, QN => n_3794);
   clk_r_REG16723_S5 : DFFS_X2 port map( D => n40617, CK => CLK, SN => 
                           RESET_BAR, Q => n52448, QN => n_3795);
   clk_r_REG16724_S5 : DFFS_X2 port map( D => n40618, CK => CLK, SN => 
                           RESET_BAR, Q => n52449, QN => n_3796);
   clk_r_REG16725_S5 : DFFS_X2 port map( D => n40619, CK => CLK, SN => 
                           RESET_BAR, Q => n52450, QN => n_3797);
   clk_r_REG16710_S5 : DFFS_X2 port map( D => n40620, CK => CLK, SN => 
                           RESET_BAR, Q => n52451, QN => n_3798);
   clk_r_REG16711_S5 : DFFS_X2 port map( D => n40621, CK => CLK, SN => 
                           RESET_BAR, Q => n52452, QN => n_3799);
   clk_r_REG16712_S5 : DFFS_X2 port map( D => n40622, CK => CLK, SN => 
                           RESET_BAR, Q => n52453, QN => n_3800);
   clk_r_REG16713_S5 : DFFS_X2 port map( D => n40623, CK => CLK, SN => 
                           RESET_BAR, Q => n52454, QN => n_3801);
   clk_r_REG16714_S5 : DFFS_X2 port map( D => n40624, CK => CLK, SN => 
                           RESET_BAR, Q => n52455, QN => n_3802);
   clk_r_REG16715_S5 : DFFS_X2 port map( D => n40625, CK => CLK, SN => 
                           RESET_BAR, Q => n52456, QN => n_3803);
   clk_r_REG16716_S5 : DFFS_X2 port map( D => n40626, CK => CLK, SN => 
                           RESET_BAR, Q => n52457, QN => n_3804);
   clk_r_REG16717_S5 : DFFS_X2 port map( D => n40627, CK => CLK, SN => 
                           RESET_BAR, Q => n52458, QN => n_3805);
   clk_r_REG16726_S5 : DFFS_X2 port map( D => n40628, CK => CLK, SN => 
                           RESET_BAR, Q => n52459, QN => n_3806);
   clk_r_REG16727_S5 : DFFS_X2 port map( D => n40632, CK => CLK, SN => 
                           RESET_BAR, Q => n52463, QN => n_3807);
   clk_r_REG16728_S5 : DFFS_X2 port map( D => n40636, CK => CLK, SN => 
                           RESET_BAR, Q => n52467, QN => n_3808);
   clk_r_REG16729_S5 : DFFS_X2 port map( D => n40637, CK => CLK, SN => 
                           RESET_BAR, Q => n52468, QN => n_3809);
   clk_r_REG16730_S5 : DFFS_X2 port map( D => n40638, CK => CLK, SN => 
                           RESET_BAR, Q => n52469, QN => n_3810);
   clk_r_REG16731_S5 : DFFS_X2 port map( D => n40642, CK => CLK, SN => 
                           RESET_BAR, Q => n52473, QN => n_3811);
   clk_r_REG16732_S5 : DFFS_X2 port map( D => n40646, CK => CLK, SN => 
                           RESET_BAR, Q => n52477, QN => n_3812);
   clk_r_REG16733_S5 : DFFS_X2 port map( D => n40647, CK => CLK, SN => 
                           RESET_BAR, Q => n52478, QN => n_3813);
   clk_r_REG16706_S5 : DFFS_X2 port map( D => n40608, CK => CLK, SN => 
                           RESET_BAR, Q => n52439, QN => n_3814);
   clk_r_REG16707_S5 : DFFS_X2 port map( D => n40609, CK => CLK, SN => 
                           RESET_BAR, Q => n52440, QN => n_3815);
   clk_r_REG16704_S5 : DFFS_X2 port map( D => n40606, CK => CLK, SN => 
                           RESET_BAR, Q => n52437, QN => n_3816);
   clk_r_REG16705_S5 : DFFS_X2 port map( D => n40607, CK => CLK, SN => 
                           RESET_BAR, Q => n52438, QN => n_3817);
   clk_r_REG16702_S5 : DFFS_X2 port map( D => n40604, CK => CLK, SN => 
                           RESET_BAR, Q => n52435, QN => n_3818);
   U3 : CLKBUF_X1 port map( A => n60059, Z => n59857);
   U4 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n53629, A3 => n53627, ZN => 
                           n60774);
   U5 : CLKBUF_X1 port map( A => n60774, Z => n60727);
   U6 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => ADD_RD1(2),
                           ZN => n41690);
   U7 : INV_X1 port map( A => n41690, ZN => n3562);
   U8 : INV_X1 port map( A => ADD_RD1(1), ZN => n58175);
   U9 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), ZN => n58170);
   U10 : NOR2_X1 port map( A1 => n58175, A2 => n58170, ZN => n41688);
   U11 : INV_X1 port map( A => n41688, ZN => n3561);
   U12 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n58170, ZN => n41692);
   U13 : INV_X1 port map( A => n41692, ZN => n3559);
   U14 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => ADD_RD2(0)
                           , ZN => n3568);
   U15 : NAND2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), ZN => n58171);
   U16 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => n58171, ZN => n3575);
   U17 : INV_X1 port map( A => ADD_RD2(1), ZN => n58176);
   U18 : NOR2_X1 port map( A1 => n58176, A2 => n58171, ZN => n3574);
   U19 : INV_X1 port map( A => ADD_RD2(2), ZN => n58177);
   U20 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n58177, ZN => n58172);
   U21 : NOR2_X1 port map( A1 => n58176, A2 => n58172, ZN => n3570);
   U22 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => n58172, ZN => n3569);
   U23 : INV_X1 port map( A => ADD_RD1(2), ZN => n58173);
   U24 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => n58173, ZN
                           => n3566);
   U25 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n58175, ZN
                           => n41686);
   U26 : INV_X1 port map( A => n41686, ZN => n3564);
   U27 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => n58175, A3 => n58173, ZN => 
                           n3560);
   U28 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n58173, ZN => n58174);
   U29 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n58174, ZN => n41687);
   U30 : INV_X1 port map( A => n41687, ZN => n3565);
   U31 : INV_X1 port map( A => ADD_RD1(3), ZN => n3558);
   U32 : NOR2_X1 port map( A1 => n58175, A2 => n58174, ZN => n41689);
   U33 : INV_X1 port map( A => n41689, ZN => n3563);
   U34 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => n58177, ZN
                           => n3573);
   U35 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => n58176, ZN
                           => n41691);
   U36 : INV_X1 port map( A => n41691, ZN => n3572);
   U37 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => n58177, A3 => n58176, ZN => 
                           n3571);
   U38 : INV_X1 port map( A => ADD_RD2(3), ZN => n3567);
   U39 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53599, ZN => n58783);
   U40 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52458, ZN => n59006);
   U41 : OAI22_X1 port map( A1 => n52458, A2 => n58783, B1 => n52512, B2 => 
                           n59006, ZN => n58178);
   U42 : INV_X1 port map( A => n58178, ZN => n3249);
   U43 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53600, ZN => n59173);
   U44 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52456, ZN => n58982);
   U45 : OAI22_X1 port map( A1 => n52456, A2 => n59173, B1 => n52513, B2 => 
                           n58982, ZN => n58179);
   U46 : INV_X1 port map( A => n58179, ZN => n3218);
   U47 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53603, ZN => n58717);
   U48 : OAI22_X1 port map( A1 => n52456, A2 => n58717, B1 => n52514, B2 => 
                           n58982, ZN => n58180);
   U49 : INV_X1 port map( A => n58180, ZN => n3121);
   U50 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53598, ZN => n58915);
   U51 : OAI22_X1 port map( A1 => n52456, A2 => n58915, B1 => n52515, B2 => 
                           n58982, ZN => n58181);
   U52 : INV_X1 port map( A => n58181, ZN => n3281);
   U53 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53601, ZN => n59213);
   U54 : OAI22_X1 port map( A1 => n52456, A2 => n59213, B1 => n52519, B2 => 
                           n58982, ZN => n58182);
   U55 : INV_X1 port map( A => n58182, ZN => n3187);
   U56 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53602, ZN => n58761);
   U57 : OAI22_X1 port map( A1 => n52456, A2 => n58761, B1 => n52520, B2 => 
                           n58982, ZN => n58183);
   U58 : INV_X1 port map( A => n58183, ZN => n3153);
   U59 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53611, ZN => n58721);
   U60 : OAI22_X1 port map( A1 => n52458, A2 => n58721, B1 => n52521, B2 => 
                           n59006, ZN => n58184);
   U61 : INV_X1 port map( A => n58184, ZN => n2865);
   U62 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53604, ZN => n58789);
   U63 : OAI22_X1 port map( A1 => n52456, A2 => n58789, B1 => n52523, B2 => 
                           n58982, ZN => n58185);
   U64 : INV_X1 port map( A => n58185, ZN => n3090);
   U65 : OAI22_X1 port map( A1 => n52458, A2 => n58717, B1 => n52525, B2 => 
                           n59006, ZN => n58186);
   U66 : INV_X1 port map( A => n58186, ZN => n3124);
   U67 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53609, ZN => n58793);
   U68 : OAI22_X1 port map( A1 => n52458, A2 => n58793, B1 => n52526, B2 => 
                           n59006, ZN => n58187);
   U69 : INV_X1 port map( A => n58187, ZN => n2930);
   U70 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53608, ZN => n58913);
   U71 : OAI22_X1 port map( A1 => n52456, A2 => n58913, B1 => n52527, B2 => 
                           n58982, ZN => n58188);
   U72 : INV_X1 port map( A => n58188, ZN => n2962);
   U73 : OAI22_X1 port map( A1 => n52458, A2 => n59213, B1 => n52532, B2 => 
                           n59006, ZN => n58189);
   U74 : INV_X1 port map( A => n58189, ZN => n3188);
   U75 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52451, ZN => n58999);
   U76 : OAI22_X1 port map( A1 => n52451, A2 => n58915, B1 => n52591, B2 => 
                           n58999, ZN => n58190);
   U77 : INV_X1 port map( A => n58190, ZN => n3287);
   U78 : CLKBUF_X1 port map( A => n59213, Z => n58736);
   U79 : OAI22_X1 port map( A1 => n52451, A2 => n58736, B1 => n52596, B2 => 
                           n58999, ZN => n58191);
   U80 : INV_X1 port map( A => n58191, ZN => n3194);
   U81 : OAI22_X1 port map( A1 => n52451, A2 => n58761, B1 => n52597, B2 => 
                           n58999, ZN => n58192);
   U82 : INV_X1 port map( A => n58192, ZN => n3158);
   U83 : CLKBUF_X1 port map( A => n58717, Z => n58745);
   U84 : OAI22_X1 port map( A1 => n52451, A2 => n58745, B1 => n52598, B2 => 
                           n58999, ZN => n58193);
   U85 : INV_X1 port map( A => n58193, ZN => n3130);
   U86 : OAI22_X1 port map( A1 => n52451, A2 => n58789, B1 => n52599, B2 => 
                           n58999, ZN => n58194);
   U87 : INV_X1 port map( A => n58194, ZN => n3096);
   U88 : OAI22_X1 port map( A1 => n52451, A2 => n58913, B1 => n52600, B2 => 
                           n58999, ZN => n58195);
   U89 : INV_X1 port map( A => n58195, ZN => n2967);
   U90 : OAI22_X1 port map( A1 => n52451, A2 => n58793, B1 => n52601, B2 => 
                           n58999, ZN => n58196);
   U91 : INV_X1 port map( A => n58196, ZN => n2936);
   U92 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53610, ZN => n58800);
   U93 : OAI22_X1 port map( A1 => n52451, A2 => n58800, B1 => n52602, B2 => 
                           n58999, ZN => n58197);
   U94 : INV_X1 port map( A => n58197, ZN => n2897);
   U95 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53612, ZN => n58759);
   U96 : OAI22_X1 port map( A1 => n52451, A2 => n58759, B1 => n52603, B2 => 
                           n58999, ZN => n58198);
   U97 : INV_X1 port map( A => n58198, ZN => n2833);
   U98 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53613, ZN => n58741);
   U99 : OAI22_X1 port map( A1 => n52451, A2 => n58741, B1 => n52604, B2 => 
                           n58999, ZN => n58199);
   U100 : INV_X1 port map( A => n58199, ZN => n2801);
   U101 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52449, ZN => n58976);
   U102 : OAI22_X1 port map( A1 => n52449, A2 => n58741, B1 => n52606, B2 => 
                           n58976, ZN => n58200);
   U103 : INV_X1 port map( A => n58200, ZN => n2802);
   U104 : OAI22_X1 port map( A1 => n52449, A2 => n58759, B1 => n52607, B2 => 
                           n58976, ZN => n58201);
   U105 : INV_X1 port map( A => n58201, ZN => n2834);
   U106 : OAI22_X1 port map( A1 => n52449, A2 => n58800, B1 => n52608, B2 => 
                           n58976, ZN => n58202);
   U107 : INV_X1 port map( A => n58202, ZN => n2898);
   U108 : OAI22_X1 port map( A1 => n52449, A2 => n58793, B1 => n52609, B2 => 
                           n58976, ZN => n58203);
   U109 : INV_X1 port map( A => n58203, ZN => n2937);
   U110 : OAI22_X1 port map( A1 => n52451, A2 => n58721, B1 => n52611, B2 => 
                           n58999, ZN => n58204);
   U111 : INV_X1 port map( A => n58204, ZN => n2871);
   U112 : OAI22_X1 port map( A1 => n52449, A2 => n58721, B1 => n52612, B2 => 
                           n58976, ZN => n58205);
   U113 : INV_X1 port map( A => n58205, ZN => n2872);
   U114 : OAI22_X1 port map( A1 => n52449, A2 => n58913, B1 => n52614, B2 => 
                           n58976, ZN => n58206);
   U115 : INV_X1 port map( A => n58206, ZN => n2968);
   U116 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53591, ZN => n58813);
   U117 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52446, ZN => n58978);
   U118 : OAI22_X1 port map( A1 => n52446, A2 => n58813, B1 => n52757, B2 => 
                           n58978, ZN => n58207);
   U119 : INV_X1 port map( A => n58207, ZN => n3517);
   U120 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53594, ZN => n58811);
   U121 : OAI22_X1 port map( A1 => n52446, A2 => n58811, B1 => n52756, B2 => 
                           n58978, ZN => n58208);
   U122 : INV_X1 port map( A => n58208, ZN => n3420);
   U123 : OAI22_X1 port map( A1 => n52449, A2 => n58813, B1 => n52752, B2 => 
                           n58976, ZN => n58209);
   U124 : INV_X1 port map( A => n58209, ZN => n3515);
   U125 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53590, ZN => n59209);
   U126 : OAI22_X1 port map( A1 => n52449, A2 => n59209, B1 => n52750, B2 => 
                           n58976, ZN => n58210);
   U127 : INV_X1 port map( A => n58210, ZN => n3548);
   U128 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53605, ZN => n58781);
   U129 : OAI22_X1 port map( A1 => n52446, A2 => n58781, B1 => n52749, B2 => 
                           n58978, ZN => n58211);
   U130 : INV_X1 port map( A => n58211, ZN => n3068);
   U131 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53597, ZN => n59166);
   U132 : OAI22_X1 port map( A1 => n52446, A2 => n59166, B1 => n52747, B2 => 
                           n58978, ZN => n58212);
   U133 : INV_X1 port map( A => n58212, ZN => n3323);
   U134 : OAI22_X1 port map( A1 => n52446, A2 => n58915, B1 => n52736, B2 => 
                           n58978, ZN => n58213);
   U135 : INV_X1 port map( A => n58213, ZN => n3293);
   U136 : OAI22_X1 port map( A1 => n52446, A2 => n58913, B1 => n52735, B2 => 
                           n58978, ZN => n58214);
   U137 : INV_X1 port map( A => n58214, ZN => n2971);
   U138 : OAI22_X1 port map( A1 => n52446, A2 => n58759, B1 => n52731, B2 => 
                           n58978, ZN => n58215);
   U139 : INV_X1 port map( A => n58215, ZN => n2843);
   U140 : OAI22_X1 port map( A1 => n52446, A2 => n58741, B1 => n52728, B2 => 
                           n58978, ZN => n58216);
   U141 : INV_X1 port map( A => n58216, ZN => n2809);
   U142 : OAI22_X1 port map( A1 => n52446, A2 => n58800, B1 => n52725, B2 => 
                           n58978, ZN => n58217);
   U143 : INV_X1 port map( A => n58217, ZN => n2905);
   U144 : OAI22_X1 port map( A1 => n52446, A2 => n58789, B1 => n52724, B2 => 
                           n58978, ZN => n58218);
   U145 : INV_X1 port map( A => n58218, ZN => n3101);
   U146 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52455, ZN => n58985);
   U147 : OAI22_X1 port map( A1 => n52455, A2 => n58789, B1 => n52723, B2 => 
                           n58985, ZN => n58219);
   U148 : INV_X1 port map( A => n58219, ZN => n3100);
   U149 : OAI22_X1 port map( A1 => n52455, A2 => n58783, B1 => n52722, B2 => 
                           n58985, ZN => n58220);
   U150 : INV_X1 port map( A => n58220, ZN => n3257);
   U151 : OAI22_X1 port map( A1 => n52455, A2 => n58741, B1 => n52721, B2 => 
                           n58985, ZN => n58221);
   U152 : INV_X1 port map( A => n58221, ZN => n2808);
   U153 : OAI22_X1 port map( A1 => n52455, A2 => n58915, B1 => n52720, B2 => 
                           n58985, ZN => n58222);
   U154 : INV_X1 port map( A => n58222, ZN => n3292);
   U155 : OAI22_X1 port map( A1 => n52455, A2 => n58717, B1 => n52717, B2 => 
                           n58985, ZN => n58223);
   U156 : INV_X1 port map( A => n58223, ZN => n3132);
   U157 : OAI22_X1 port map( A1 => n52455, A2 => n59213, B1 => n52713, B2 => 
                           n58985, ZN => n58224);
   U158 : INV_X1 port map( A => n58224, ZN => n3196);
   U159 : OAI22_X1 port map( A1 => n52455, A2 => n59209, B1 => n52712, B2 => 
                           n58985, ZN => n58225);
   U160 : INV_X1 port map( A => n58225, ZN => n3547);
   U161 : OAI22_X1 port map( A1 => n52446, A2 => n59173, B1 => n52710, B2 => 
                           n58978, ZN => n58226);
   U162 : INV_X1 port map( A => n58226, ZN => n3221);
   U163 : OAI22_X1 port map( A1 => n52451, A2 => n59173, B1 => n52707, B2 => 
                           n58999, ZN => n58227);
   U164 : INV_X1 port map( A => n58227, ZN => n3219);
   U165 : OAI22_X1 port map( A1 => n52458, A2 => n59209, B1 => n52705, B2 => 
                           n59006, ZN => n58228);
   U166 : INV_X1 port map( A => n58228, ZN => n3546);
   U167 : OAI22_X1 port map( A1 => n52456, A2 => n59209, B1 => n52704, B2 => 
                           n58982, ZN => n58229);
   U168 : INV_X1 port map( A => n58229, ZN => n3545);
   U169 : OAI22_X1 port map( A1 => n52456, A2 => n58759, B1 => n52695, B2 => 
                           n58982, ZN => n58230);
   U170 : INV_X1 port map( A => n58230, ZN => n2838);
   U171 : OAI22_X1 port map( A1 => n52456, A2 => n58741, B1 => n52694, B2 => 
                           n58982, ZN => n58231);
   U172 : INV_X1 port map( A => n58231, ZN => n2806);
   U173 : OAI22_X1 port map( A1 => n52458, A2 => n58759, B1 => n52691, B2 => 
                           n59006, ZN => n58232);
   U174 : INV_X1 port map( A => n58232, ZN => n2836);
   U175 : OAI22_X1 port map( A1 => n52458, A2 => n58741, B1 => n52690, B2 => 
                           n59006, ZN => n58233);
   U176 : INV_X1 port map( A => n58233, ZN => n2804);
   U177 : OAI22_X1 port map( A1 => n52458, A2 => n58761, B1 => n52681, B2 => 
                           n59006, ZN => n58234);
   U178 : INV_X1 port map( A => n58234, ZN => n3160);
   U179 : OAI22_X1 port map( A1 => n52458, A2 => n58789, B1 => n52678, B2 => 
                           n59006, ZN => n58235);
   U180 : INV_X1 port map( A => n58235, ZN => n3098);
   U181 : OAI22_X1 port map( A1 => n52456, A2 => n58800, B1 => n52664, B2 => 
                           n58982, ZN => n58236);
   U182 : INV_X1 port map( A => n58236, ZN => n2900);
   U183 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53607, ZN => n58730);
   U184 : OAI22_X1 port map( A1 => n52456, A2 => n58730, B1 => n52661, B2 => 
                           n58982, ZN => n58237);
   U185 : INV_X1 port map( A => n58237, ZN => n3004);
   U186 : OAI22_X1 port map( A1 => n52455, A2 => n58813, B1 => n52659, B2 => 
                           n58985, ZN => n58238);
   U187 : INV_X1 port map( A => n58238, ZN => n3513);
   U188 : OAI22_X1 port map( A1 => n52455, A2 => n58811, B1 => n52658, B2 => 
                           n58985, ZN => n58239);
   U189 : INV_X1 port map( A => n58239, ZN => n3417);
   U190 : OAI22_X1 port map( A1 => n52455, A2 => n58730, B1 => n52657, B2 => 
                           n58985, ZN => n58240);
   U191 : INV_X1 port map( A => n58240, ZN => n3003);
   U192 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53596, ZN => n58819);
   U193 : OAI22_X1 port map( A1 => n52455, A2 => n58819, B1 => n52655, B2 => 
                           n58985, ZN => n58241);
   U194 : INV_X1 port map( A => n58241, ZN => n3353);
   U195 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53595, ZN => n58910);
   U196 : OAI22_X1 port map( A1 => n52455, A2 => n58910, B1 => n52654, B2 => 
                           n58985, ZN => n58242);
   U197 : INV_X1 port map( A => n58242, ZN => n3385);
   U198 : OAI22_X1 port map( A1 => n52455, A2 => n58781, B1 => n52653, B2 => 
                           n58985, ZN => n58243);
   U199 : INV_X1 port map( A => n58243, ZN => n3065);
   U200 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53592, ZN => n59169);
   U201 : OAI22_X1 port map( A1 => n52455, A2 => n59169, B1 => n52652, B2 => 
                           n58985, ZN => n58244);
   U202 : INV_X1 port map( A => n58244, ZN => n3479);
   U203 : OAI22_X1 port map( A1 => n52455, A2 => n59166, B1 => n52651, B2 => 
                           n58985, ZN => n58245);
   U204 : INV_X1 port map( A => n58245, ZN => n3316);
   U205 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53593, ZN => n58826);
   U206 : OAI22_X1 port map( A1 => n52455, A2 => n58826, B1 => n52650, B2 => 
                           n58985, ZN => n58246);
   U207 : INV_X1 port map( A => n58246, ZN => n3449);
   U208 : OAI22_X1 port map( A1 => n52449, A2 => n58915, B1 => n52648, B2 => 
                           n58976, ZN => n58247);
   U209 : INV_X1 port map( A => n58247, ZN => n3289);
   U210 : OAI22_X1 port map( A1 => n52449, A2 => n58783, B1 => n52647, B2 => 
                           n58976, ZN => n58248);
   U211 : INV_X1 port map( A => n58248, ZN => n3255);
   U212 : OAI22_X1 port map( A1 => n52446, A2 => n58730, B1 => n52645, B2 => 
                           n58978, ZN => n58249);
   U213 : INV_X1 port map( A => n58249, ZN => n3000);
   U214 : OAI22_X1 port map( A1 => n52458, A2 => n59169, B1 => n52642, B2 => 
                           n59006, ZN => n58250);
   U215 : INV_X1 port map( A => n58250, ZN => n3478);
   U216 : OAI22_X1 port map( A1 => n52456, A2 => n58910, B1 => n52641, B2 => 
                           n58982, ZN => n58251);
   U217 : INV_X1 port map( A => n58251, ZN => n3384);
   U218 : OAI22_X1 port map( A1 => n52458, A2 => n58819, B1 => n52639, B2 => 
                           n59006, ZN => n58252);
   U219 : INV_X1 port map( A => n58252, ZN => n3352);
   U220 : OAI22_X1 port map( A1 => n52458, A2 => n58910, B1 => n52638, B2 => 
                           n59006, ZN => n58253);
   U221 : INV_X1 port map( A => n58253, ZN => n3383);
   U222 : OAI22_X1 port map( A1 => n52456, A2 => n58813, B1 => n52637, B2 => 
                           n58982, ZN => n58254);
   U223 : INV_X1 port map( A => n58254, ZN => n3512);
   U224 : OAI22_X1 port map( A1 => n52456, A2 => n58819, B1 => n52636, B2 => 
                           n58982, ZN => n58255);
   U225 : INV_X1 port map( A => n58255, ZN => n3351);
   U226 : OAI22_X1 port map( A1 => n52458, A2 => n58811, B1 => n52634, B2 => 
                           n59006, ZN => n58256);
   U227 : INV_X1 port map( A => n58256, ZN => n3416);
   U228 : OAI22_X1 port map( A1 => n52456, A2 => n58811, B1 => n52632, B2 => 
                           n58982, ZN => n58257);
   U229 : INV_X1 port map( A => n58257, ZN => n3415);
   U230 : OAI22_X1 port map( A1 => n52458, A2 => n58730, B1 => n52631, B2 => 
                           n59006, ZN => n58258);
   U231 : INV_X1 port map( A => n58258, ZN => n2999);
   U232 : OAI22_X1 port map( A1 => n52456, A2 => n58781, B1 => n52630, B2 => 
                           n58982, ZN => n58259);
   U233 : INV_X1 port map( A => n58259, ZN => n3064);
   U234 : OAI22_X1 port map( A1 => n52456, A2 => n58826, B1 => n52629, B2 => 
                           n58982, ZN => n58260);
   U235 : INV_X1 port map( A => n58260, ZN => n3447);
   U236 : OAI22_X1 port map( A1 => n52458, A2 => n58781, B1 => n52628, B2 => 
                           n59006, ZN => n58261);
   U237 : INV_X1 port map( A => n58261, ZN => n3063);
   U238 : OAI22_X1 port map( A1 => n52458, A2 => n59166, B1 => n52624, B2 => 
                           n59006, ZN => n58262);
   U239 : INV_X1 port map( A => n58262, ZN => n3314);
   U240 : OAI22_X1 port map( A1 => n52449, A2 => n59213, B1 => n52619, B2 => 
                           n58976, ZN => n58263);
   U241 : INV_X1 port map( A => n58263, ZN => n3195);
   U242 : OAI22_X1 port map( A1 => n52449, A2 => n58761, B1 => n52618, B2 => 
                           n58976, ZN => n58264);
   U243 : INV_X1 port map( A => n58264, ZN => n3159);
   U244 : OAI22_X1 port map( A1 => n52449, A2 => n58717, B1 => n52617, B2 => 
                           n58976, ZN => n58265);
   U245 : INV_X1 port map( A => n58265, ZN => n3131);
   U246 : OAI22_X1 port map( A1 => n52449, A2 => n58789, B1 => n52616, B2 => 
                           n58976, ZN => n58266);
   U247 : INV_X1 port map( A => n58266, ZN => n3097);
   U248 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52459, ZN => n58993);
   U249 : OAI22_X1 port map( A1 => n52459, A2 => n58793, B1 => n52954, B2 => 
                           n58993, ZN => n58267);
   U250 : INV_X1 port map( A => n58267, ZN => n2942);
   U251 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52436, ZN => n59124);
   U252 : OAI22_X1 port map( A1 => n52436, A2 => n58761, B1 => n53421, B2 => 
                           n59124, ZN => n58268);
   U253 : INV_X1 port map( A => n58268, ZN => n3152);
   U254 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52445, ZN => n58967);
   U255 : OAI22_X1 port map( A1 => n52445, A2 => n58783, B1 => n53122, B2 => 
                           n58967, ZN => n58269);
   U256 : INV_X1 port map( A => n58269, ZN => n3268);
   U257 : CLKBUF_X1 port map( A => n58730, Z => n58616);
   U258 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52454, ZN => n59120);
   U259 : OAI22_X1 port map( A1 => n52454, A2 => n58616, B1 => n53064, B2 => 
                           n59120, ZN => n58270);
   U260 : INV_X1 port map( A => n58270, ZN => n2985);
   U261 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52478, ZN => n58980);
   U262 : OAI22_X1 port map( A1 => n52478, A2 => n58789, B1 => n52914, B2 => 
                           n58980, ZN => n58271);
   U263 : INV_X1 port map( A => n58271, ZN => n3106);
   U264 : OAI22_X1 port map( A1 => n52445, A2 => n58745, B1 => n53120, B2 => 
                           n58967, ZN => n58272);
   U265 : INV_X1 port map( A => n58272, ZN => n3117);
   U266 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52469, ZN => n58996);
   U267 : OAI22_X1 port map( A1 => n52469, A2 => n58813, B1 => n52918, B2 => 
                           n58996, ZN => n58273);
   U268 : INV_X1 port map( A => n58273, ZN => n3523);
   U269 : OAI22_X1 port map( A1 => n52478, A2 => n58819, B1 => n52920, B2 => 
                           n58980, ZN => n58274);
   U270 : INV_X1 port map( A => n58274, ZN => n3360);
   U271 : OAI22_X1 port map( A1 => n52478, A2 => n58741, B1 => n53389, B2 => 
                           n58980, ZN => n58275);
   U272 : INV_X1 port map( A => n58275, ZN => n2799);
   U273 : OAI22_X1 port map( A1 => n52436, A2 => n58759, B1 => n53425, B2 => 
                           n59124, ZN => n58276);
   U274 : INV_X1 port map( A => n58276, ZN => n2832);
   U275 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52444, ZN => n59128);
   U276 : OAI22_X1 port map( A1 => n52444, A2 => n58616, B1 => n53067, B2 => 
                           n59128, ZN => n58277);
   U277 : INV_X1 port map( A => n58277, ZN => n2988);
   U278 : OAI22_X1 port map( A1 => n52469, A2 => n58730, B1 => n52910, B2 => 
                           n58996, ZN => n58278);
   U279 : INV_X1 port map( A => n58278, ZN => n3010);
   U280 : OAI22_X1 port map( A1 => n52459, A2 => n58789, B1 => n53387, B2 => 
                           n58993, ZN => n58279);
   U281 : INV_X1 port map( A => n58279, ZN => n3087);
   U282 : OAI22_X1 port map( A1 => n52459, A2 => n58783, B1 => n52832, B2 => 
                           n58993, ZN => n58280);
   U283 : INV_X1 port map( A => n58280, ZN => n3259);
   U284 : OAI22_X1 port map( A1 => n52459, A2 => n58915, B1 => n52831, B2 => 
                           n58993, ZN => n58281);
   U285 : INV_X1 port map( A => n58281, ZN => n3298);
   U286 : OAI22_X1 port map( A1 => n52445, A2 => n58616, B1 => n53068, B2 => 
                           n58967, ZN => n58282);
   U287 : INV_X1 port map( A => n58282, ZN => n2989);
   U288 : OAI22_X1 port map( A1 => n52478, A2 => n58915, B1 => n52828, B2 => 
                           n58980, ZN => n58283);
   U289 : INV_X1 port map( A => n58283, ZN => n3296);
   U290 : OAI22_X1 port map( A1 => n52444, A2 => n58741, B1 => n53114, B2 => 
                           n59128, ZN => n58284);
   U291 : INV_X1 port map( A => n58284, ZN => n2819);
   U292 : OAI22_X1 port map( A1 => n52459, A2 => n58741, B1 => n53372, B2 => 
                           n58993, ZN => n58285);
   U293 : INV_X1 port map( A => n58285, ZN => n2798);
   U294 : OAI22_X1 port map( A1 => n52469, A2 => n58811, B1 => n52907, B2 => 
                           n58996, ZN => n58286);
   U295 : INV_X1 port map( A => n58286, ZN => n3424);
   U296 : OAI22_X1 port map( A1 => n52478, A2 => n58781, B1 => n52823, B2 => 
                           n58980, ZN => n58287);
   U297 : INV_X1 port map( A => n58287, ZN => n3070);
   U298 : OAI22_X1 port map( A1 => n52478, A2 => n58826, B1 => n52922, B2 => 
                           n58980, ZN => n58288);
   U299 : INV_X1 port map( A => n58288, ZN => n3456);
   U300 : OAI22_X1 port map( A1 => n52478, A2 => n58721, B1 => n53361, B2 => 
                           n58980, ZN => n58289);
   U301 : INV_X1 port map( A => n58289, ZN => n2864);
   U302 : OAI22_X1 port map( A1 => n52459, A2 => n58717, B1 => n52820, B2 => 
                           n58993, ZN => n58290);
   U303 : INV_X1 port map( A => n58290, ZN => n3137);
   U304 : OAI22_X1 port map( A1 => n52469, A2 => n58717, B1 => n53360, B2 => 
                           n58996, ZN => n58291);
   U305 : INV_X1 port map( A => n58291, ZN => n3120);
   U306 : OAI22_X1 port map( A1 => n52478, A2 => n58745, B1 => n52819, B2 => 
                           n58980, ZN => n58292);
   U307 : INV_X1 port map( A => n58292, ZN => n3112);
   U308 : OAI22_X1 port map( A1 => n52444, A2 => n59173, B1 => n53109, B2 => 
                           n59128, ZN => n58293);
   U309 : INV_X1 port map( A => n58293, ZN => n3232);
   U310 : OAI22_X1 port map( A1 => n52459, A2 => n58616, B1 => n52905, B2 => 
                           n58993, ZN => n58294);
   U311 : INV_X1 port map( A => n58294, ZN => n2984);
   U312 : OAI22_X1 port map( A1 => n52444, A2 => n58793, B1 => n53106, B2 => 
                           n59128, ZN => n58295);
   U313 : INV_X1 port map( A => n58295, ZN => n2944);
   U314 : OAI22_X1 port map( A1 => n52478, A2 => n59169, B1 => n52923, B2 => 
                           n58980, ZN => n58296);
   U315 : INV_X1 port map( A => n58296, ZN => n3489);
   U316 : OAI22_X1 port map( A1 => n52444, A2 => n58913, B1 => n53105, B2 => 
                           n59128, ZN => n58297);
   U317 : INV_X1 port map( A => n58297, ZN => n2981);
   U318 : OAI22_X1 port map( A1 => n52478, A2 => n58913, B1 => n52814, B2 => 
                           n58980, ZN => n58298);
   U319 : INV_X1 port map( A => n58298, ZN => n2973);
   U320 : OAI22_X1 port map( A1 => n52478, A2 => n58813, B1 => n52904, B2 => 
                           n58980, ZN => n58299);
   U321 : INV_X1 port map( A => n58299, ZN => n3520);
   U322 : OAI22_X1 port map( A1 => n52436, A2 => n59166, B1 => n52902, B2 => 
                           n59124, ZN => n58300);
   U323 : INV_X1 port map( A => n58300, ZN => n3330);
   U324 : OAI22_X1 port map( A1 => n52444, A2 => n59209, B1 => n53043, B2 => 
                           n59128, ZN => n58301);
   U325 : INV_X1 port map( A => n58301, ZN => n3555);
   U326 : OAI22_X1 port map( A1 => n52469, A2 => n58783, B1 => n52836, B2 => 
                           n58996, ZN => n58302);
   U327 : INV_X1 port map( A => n58302, ZN => n3263);
   U328 : OAI22_X1 port map( A1 => n52451, A2 => n58781, B1 => n53338, B2 => 
                           n58999, ZN => n58303);
   U329 : INV_X1 port map( A => n58303, ZN => n3056);
   U330 : OAI22_X1 port map( A1 => n52444, A2 => n58745, B1 => n53101, B2 => 
                           n59128, ZN => n58304);
   U331 : INV_X1 port map( A => n58304, ZN => n3114);
   U332 : OAI22_X1 port map( A1 => n52469, A2 => n58761, B1 => n52811, B2 => 
                           n58996, ZN => n58305);
   U333 : INV_X1 port map( A => n58305, ZN => n3167);
   U334 : OAI22_X1 port map( A1 => n52459, A2 => n59173, B1 => n52901, B2 => 
                           n58993, ZN => n58306);
   U335 : INV_X1 port map( A => n58306, ZN => n3230);
   U336 : OAI22_X1 port map( A1 => n52478, A2 => n58730, B1 => n52809, B2 => 
                           n58980, ZN => n58307);
   U337 : INV_X1 port map( A => n58307, ZN => n3006);
   U338 : OAI22_X1 port map( A1 => n52459, A2 => n59213, B1 => n52808, B2 => 
                           n58993, ZN => n58308);
   U339 : INV_X1 port map( A => n58308, ZN => n3202);
   U340 : OAI22_X1 port map( A1 => n52478, A2 => n59213, B1 => n52807, B2 => 
                           n58980, ZN => n58309);
   U341 : INV_X1 port map( A => n58309, ZN => n3201);
   U342 : OAI22_X1 port map( A1 => n52446, A2 => n58783, B1 => n53337, B2 => 
                           n58978, ZN => n58310);
   U343 : INV_X1 port map( A => n58310, ZN => n3248);
   U344 : OAI22_X1 port map( A1 => n52444, A2 => n58761, B1 => n53100, B2 => 
                           n59128, ZN => n58311);
   U345 : INV_X1 port map( A => n58311, ZN => n3171);
   U346 : OAI22_X1 port map( A1 => n52469, A2 => n58736, B1 => n52804, B2 => 
                           n58996, ZN => n58312);
   U347 : INV_X1 port map( A => n58312, ZN => n3175);
   U348 : OAI22_X1 port map( A1 => n52478, A2 => n58793, B1 => n52803, B2 => 
                           n58980, ZN => n58313);
   U349 : INV_X1 port map( A => n58313, ZN => n2938);
   U350 : OAI22_X1 port map( A1 => n52469, A2 => n59173, B1 => n52898, B2 => 
                           n58996, ZN => n58314);
   U351 : INV_X1 port map( A => n58314, ZN => n3229);
   U352 : CLKBUF_X1 port map( A => n58721, Z => n58725);
   U353 : OAI22_X1 port map( A1 => n52436, A2 => n58725, B1 => n52842, B2 => 
                           n59124, ZN => n58315);
   U354 : INV_X1 port map( A => n58315, ZN => n2874);
   U355 : OAI22_X1 port map( A1 => n52436, A2 => n58793, B1 => n52843, B2 => 
                           n59124, ZN => n58316);
   U356 : INV_X1 port map( A => n58316, ZN => n2939);
   U357 : OAI22_X1 port map( A1 => n52436, A2 => n58913, B1 => n52844, B2 => 
                           n59124, ZN => n58317);
   U358 : INV_X1 port map( A => n58317, ZN => n2974);
   U359 : OAI22_X1 port map( A1 => n52478, A2 => n59209, B1 => n52895, B2 => 
                           n58980, ZN => n58318);
   U360 : INV_X1 port map( A => n58318, ZN => n3552);
   U361 : OAI22_X1 port map( A1 => n52449, A2 => n58819, B1 => n52796, B2 => 
                           n58976, ZN => n58319);
   U362 : INV_X1 port map( A => n58319, ZN => n3359);
   U363 : OAI22_X1 port map( A1 => n52459, A2 => n59209, B1 => n52890, B2 => 
                           n58993, ZN => n58320);
   U364 : INV_X1 port map( A => n58320, ZN => n3551);
   U365 : OAI22_X1 port map( A1 => n52446, A2 => n58717, B1 => n52794, B2 => 
                           n58978, ZN => n58321);
   U366 : INV_X1 port map( A => n58321, ZN => n3135);
   U367 : OAI22_X1 port map( A1 => n52449, A2 => n58811, B1 => n52793, B2 => 
                           n58976, ZN => n58322);
   U368 : INV_X1 port map( A => n58322, ZN => n3423);
   U369 : OAI22_X1 port map( A1 => n52451, A2 => n58819, B1 => n52792, B2 => 
                           n58999, ZN => n58323);
   U370 : INV_X1 port map( A => n58323, ZN => n3358);
   U371 : OAI22_X1 port map( A1 => n52446, A2 => n58721, B1 => n53295, B2 => 
                           n58978, ZN => n58324);
   U372 : INV_X1 port map( A => n58324, ZN => n2862);
   U373 : OAI22_X1 port map( A1 => n52449, A2 => n59173, B1 => n53292, B2 => 
                           n58976, ZN => n58325);
   U374 : INV_X1 port map( A => n58325, ZN => n3215);
   U375 : OAI22_X1 port map( A1 => n52446, A2 => n59169, B1 => n52788, B2 => 
                           n58978, ZN => n58326);
   U376 : INV_X1 port map( A => n58326, ZN => n3486);
   U377 : OAI22_X1 port map( A1 => n52451, A2 => n58730, B1 => n53285, B2 => 
                           n58999, ZN => n58327);
   U378 : INV_X1 port map( A => n58327, ZN => n2992);
   U379 : OAI22_X1 port map( A1 => n52449, A2 => n59166, B1 => n52787, B2 => 
                           n58976, ZN => n58328);
   U380 : INV_X1 port map( A => n58328, ZN => n3326);
   U381 : OAI22_X1 port map( A1 => n52458, A2 => n58913, B1 => n53284, B2 => 
                           n59006, ZN => n58329);
   U382 : INV_X1 port map( A => n58329, ZN => n2958);
   U383 : OAI22_X1 port map( A1 => n52449, A2 => n58730, B1 => n53280, B2 => 
                           n58976, ZN => n58330);
   U384 : INV_X1 port map( A => n58330, ZN => n2991);
   U385 : OAI22_X1 port map( A1 => n52455, A2 => n58725, B1 => n53268, B2 => 
                           n58985, ZN => n58331);
   U386 : INV_X1 port map( A => n58331, ZN => n2861);
   U387 : OAI22_X1 port map( A1 => n52456, A2 => n58725, B1 => n53263, B2 => 
                           n58982, ZN => n58332);
   U388 : INV_X1 port map( A => n58332, ZN => n2860);
   U389 : OAI22_X1 port map( A1 => n52454, A2 => n58761, B1 => n53092, B2 => 
                           n59120, ZN => n58333);
   U390 : INV_X1 port map( A => n58333, ZN => n3170);
   U391 : OAI22_X1 port map( A1 => n52445, A2 => n59213, B1 => n53099, B2 => 
                           n58967, ZN => n58334);
   U392 : INV_X1 port map( A => n58334, ZN => n3182);
   U393 : OAI22_X1 port map( A1 => n52454, A2 => n58721, B1 => n53073, B2 => 
                           n59120, ZN => n58335);
   U394 : INV_X1 port map( A => n58335, ZN => n2881);
   U395 : OAI22_X1 port map( A1 => n52444, A2 => n58910, B1 => n53020, B2 => 
                           n59128, ZN => n58336);
   U396 : INV_X1 port map( A => n58336, ZN => n3374);
   U397 : OAI22_X1 port map( A1 => n52444, A2 => n58819, B1 => n53002, B2 => 
                           n59128, ZN => n58337);
   U398 : INV_X1 port map( A => n58337, ZN => n3342);
   U399 : OAI22_X1 port map( A1 => n52444, A2 => n58721, B1 => n53076, B2 => 
                           n59128, ZN => n58338);
   U400 : INV_X1 port map( A => n58338, ZN => n2884);
   U401 : OAI22_X1 port map( A1 => n52459, A2 => n58826, B1 => n52928, B2 => 
                           n58993, ZN => n58339);
   U402 : INV_X1 port map( A => n58339, ZN => n3457);
   U403 : OAI22_X1 port map( A1 => n52445, A2 => n58721, B1 => n53077, B2 => 
                           n58967, ZN => n58340);
   U404 : INV_X1 port map( A => n58340, ZN => n2885);
   U405 : OAI22_X1 port map( A1 => n52478, A2 => n58811, B1 => n52931, B2 => 
                           n58980, ZN => n58341);
   U406 : INV_X1 port map( A => n58341, ZN => n3428);
   U407 : OAI22_X1 port map( A1 => n52459, A2 => n59169, B1 => n52933, B2 => 
                           n58993, ZN => n58342);
   U408 : INV_X1 port map( A => n58342, ZN => n3492);
   U409 : OAI22_X1 port map( A1 => n52444, A2 => n58736, B1 => n53098, B2 => 
                           n59128, ZN => n58343);
   U410 : INV_X1 port map( A => n58343, ZN => n3181);
   U411 : OAI22_X1 port map( A1 => n52459, A2 => n58761, B1 => n52815, B2 => 
                           n58993, ZN => n58344);
   U412 : INV_X1 port map( A => n58344, ZN => n3168);
   U413 : OAI22_X1 port map( A1 => n52445, A2 => n59173, B1 => n53144, B2 => 
                           n58967, ZN => n58345);
   U414 : INV_X1 port map( A => n58345, ZN => n3236);
   U415 : OAI22_X1 port map( A1 => n52454, A2 => n58800, B1 => n52977, B2 => 
                           n59120, ZN => n58346);
   U416 : INV_X1 port map( A => n58346, ZN => n2914);
   U417 : OAI22_X1 port map( A1 => n52454, A2 => n58913, B1 => n52975, B2 => 
                           n59120, ZN => n58347);
   U418 : INV_X1 port map( A => n58347, ZN => n2978);
   U419 : OAI22_X1 port map( A1 => n52454, A2 => n58781, B1 => n52974, B2 => 
                           n59120, ZN => n58348);
   U420 : INV_X1 port map( A => n58348, ZN => n3075);
   U421 : OAI22_X1 port map( A1 => n52454, A2 => n58789, B1 => n52973, B2 => 
                           n59120, ZN => n58349);
   U422 : INV_X1 port map( A => n58349, ZN => n3107);
   U423 : OAI22_X1 port map( A1 => n52449, A2 => n58910, B1 => n52760, B2 => 
                           n58976, ZN => n58350);
   U424 : INV_X1 port map( A => n58350, ZN => n3387);
   U425 : OAI22_X1 port map( A1 => n52454, A2 => n58717, B1 => n52972, B2 => 
                           n59120, ZN => n58351);
   U426 : INV_X1 port map( A => n58351, ZN => n3140);
   U427 : OAI22_X1 port map( A1 => n52469, A2 => n58781, B1 => n52971, B2 => 
                           n58996, ZN => n58352);
   U428 : INV_X1 port map( A => n58352, ZN => n3074);
   U429 : OAI22_X1 port map( A1 => n52449, A2 => n58826, B1 => n52762, B2 => 
                           n58976, ZN => n58353);
   U430 : INV_X1 port map( A => n58353, ZN => n3451);
   U431 : CLKBUF_X1 port map( A => n58741, Z => n58655);
   U432 : OAI22_X1 port map( A1 => n52469, A2 => n58655, B1 => n52970, B2 => 
                           n58996, ZN => n58354);
   U433 : INV_X1 port map( A => n58354, ZN => n2791);
   U434 : OAI22_X1 port map( A1 => n52459, A2 => n58819, B1 => n52969, B2 => 
                           n58993, ZN => n58355);
   U435 : INV_X1 port map( A => n58355, ZN => n3364);
   U436 : OAI22_X1 port map( A1 => n52454, A2 => n58759, B1 => n52978, B2 => 
                           n59120, ZN => n58356);
   U437 : INV_X1 port map( A => n58356, ZN => n2850);
   U438 : OAI22_X1 port map( A1 => n52459, A2 => n58913, B1 => n52966, B2 => 
                           n58993, ZN => n58357);
   U439 : INV_X1 port map( A => n58357, ZN => n2977);
   U440 : OAI22_X1 port map( A1 => n52445, A2 => n59166, B1 => n52979, B2 => 
                           n58967, ZN => n58358);
   U441 : INV_X1 port map( A => n58358, ZN => n3332);
   U442 : OAI22_X1 port map( A1 => n52436, A2 => n58655, B1 => n52964, B2 => 
                           n59124, ZN => n58359);
   U443 : INV_X1 port map( A => n58359, ZN => n2790);
   U444 : OAI22_X1 port map( A1 => n52454, A2 => n58736, B1 => n53091, B2 => 
                           n59120, ZN => n58360);
   U445 : INV_X1 port map( A => n58360, ZN => n3178);
   U446 : OAI22_X1 port map( A1 => n52459, A2 => n58910, B1 => n52962, B2 => 
                           n58993, ZN => n58361);
   U447 : INV_X1 port map( A => n58361, ZN => n3394);
   U448 : OAI22_X1 port map( A1 => n52454, A2 => n59166, B1 => n52980, B2 => 
                           n59120, ZN => n58362);
   U449 : INV_X1 port map( A => n58362, ZN => n3333);
   U450 : OAI22_X1 port map( A1 => n52446, A2 => n58826, B1 => n52764, B2 => 
                           n58978, ZN => n58363);
   U451 : INV_X1 port map( A => n58363, ZN => n3453);
   U452 : OAI22_X1 port map( A1 => n52444, A2 => n58783, B1 => n53095, B2 => 
                           n59128, ZN => n58364);
   U453 : INV_X1 port map( A => n58364, ZN => n3266);
   U454 : OAI22_X1 port map( A1 => n52445, A2 => n58655, B1 => n53171, B2 => 
                           n58967, ZN => n58365);
   U455 : INV_X1 port map( A => n58365, ZN => n2793);
   U456 : OAI22_X1 port map( A1 => n52454, A2 => n58655, B1 => n53178, B2 => 
                           n59120, ZN => n58366);
   U457 : INV_X1 port map( A => n58366, ZN => n2794);
   U458 : OAI22_X1 port map( A1 => n52445, A2 => n58793, B1 => n53179, B2 => 
                           n58967, ZN => n58367);
   U459 : INV_X1 port map( A => n58367, ZN => n2948);
   U460 : OAI22_X1 port map( A1 => n52454, A2 => n59209, B1 => n53180, B2 => 
                           n59120, ZN => n58368);
   U461 : INV_X1 port map( A => n58368, ZN => n3556);
   U462 : OAI22_X1 port map( A1 => n52445, A2 => n59209, B1 => n53181, B2 => 
                           n58967, ZN => n58369);
   U463 : INV_X1 port map( A => n58369, ZN => n3557);
   U464 : OAI22_X1 port map( A1 => n52469, A2 => n58819, B1 => n52959, B2 => 
                           n58996, ZN => n58370);
   U465 : INV_X1 port map( A => n58370, ZN => n3362);
   U466 : OAI22_X1 port map( A1 => n52436, A2 => n58915, B1 => n52853, B2 => 
                           n59124, ZN => n58371);
   U467 : INV_X1 port map( A => n58371, ZN => n3300);
   U468 : OAI22_X1 port map( A1 => n52449, A2 => n59169, B1 => n52767, B2 => 
                           n58976, ZN => n58372);
   U469 : INV_X1 port map( A => n58372, ZN => n3484);
   U470 : OAI22_X1 port map( A1 => n52451, A2 => n58811, B1 => n52768, B2 => 
                           n58999, ZN => n58373);
   U471 : INV_X1 port map( A => n58373, ZN => n3421);
   U472 : OAI22_X1 port map( A1 => n52446, A2 => n59209, B1 => n52769, B2 => 
                           n58978, ZN => n58374);
   U473 : INV_X1 port map( A => n58374, ZN => n3549);
   U474 : OAI22_X1 port map( A1 => n52451, A2 => n58826, B1 => n52770, B2 => 
                           n58999, ZN => n58375);
   U475 : INV_X1 port map( A => n58375, ZN => n3454);
   U476 : OAI22_X1 port map( A1 => n52451, A2 => n59169, B1 => n52771, B2 => 
                           n58999, ZN => n58376);
   U477 : INV_X1 port map( A => n58376, ZN => n3485);
   U478 : OAI22_X1 port map( A1 => n52446, A2 => n59213, B1 => n52772, B2 => 
                           n58978, ZN => n58377);
   U479 : INV_X1 port map( A => n58377, ZN => n3198);
   U480 : OAI22_X1 port map( A1 => n52451, A2 => n59166, B1 => n53196, B2 => 
                           n58999, ZN => n58378);
   U481 : INV_X1 port map( A => n58378, ZN => n3312);
   U482 : OAI22_X1 port map( A1 => n52469, A2 => n58721, B1 => n52957, B2 => 
                           n58996, ZN => n58379);
   U483 : INV_X1 port map( A => n58379, ZN => n2879);
   U484 : OAI22_X1 port map( A1 => n52451, A2 => n59209, B1 => n52773, B2 => 
                           n58999, ZN => n58380);
   U485 : INV_X1 port map( A => n58380, ZN => n3550);
   U486 : OAI22_X1 port map( A1 => n52436, A2 => n58783, B1 => n52852, B2 => 
                           n59124, ZN => n58381);
   U487 : INV_X1 port map( A => n58381, ZN => n3264);
   U488 : OAI22_X1 port map( A1 => n52436, A2 => n59213, B1 => n52851, B2 => 
                           n59124, ZN => n58382);
   U489 : INV_X1 port map( A => n58382, ZN => n3204);
   U490 : OAI22_X1 port map( A1 => n52454, A2 => n58783, B1 => n53089, B2 => 
                           n59120, ZN => n58383);
   U491 : INV_X1 port map( A => n58383, ZN => n3265);
   U492 : OAI22_X1 port map( A1 => n52478, A2 => n58910, B1 => n52953, B2 => 
                           n58980, ZN => n58384);
   U493 : INV_X1 port map( A => n58384, ZN => n3393);
   U494 : OAI22_X1 port map( A1 => n52436, A2 => n58717, B1 => n52850, B2 => 
                           n59124, ZN => n58385);
   U495 : INV_X1 port map( A => n58385, ZN => n3139);
   U496 : OAI22_X1 port map( A1 => n52436, A2 => n58789, B1 => n52849, B2 => 
                           n59124, ZN => n58386);
   U497 : INV_X1 port map( A => n58386, ZN => n3105);
   U498 : OAI22_X1 port map( A1 => n52451, A2 => n58813, B1 => n52776, B2 => 
                           n58999, ZN => n58387);
   U499 : INV_X1 port map( A => n58387, ZN => n3519);
   U500 : OAI22_X1 port map( A1 => n52454, A2 => n58793, B1 => n52976, B2 => 
                           n59120, ZN => n58388);
   U501 : INV_X1 port map( A => n58388, ZN => n2943);
   U502 : OAI22_X1 port map( A1 => n52446, A2 => n58761, B1 => n52780, B2 => 
                           n58978, ZN => n58389);
   U503 : INV_X1 port map( A => n58389, ZN => n3164);
   U504 : OAI22_X1 port map( A1 => n52446, A2 => n58819, B1 => n52783, B2 => 
                           n58978, ZN => n58390);
   U505 : INV_X1 port map( A => n58390, ZN => n3356);
   U506 : OAI22_X1 port map( A1 => n52458, A2 => n58800, B1 => n53214, B2 => 
                           n59006, ZN => n58391);
   U507 : INV_X1 port map( A => n58391, ZN => n2895);
   U508 : OAI22_X1 port map( A1 => n52478, A2 => n59166, B1 => n52862, B2 => 
                           n58980, ZN => n58392);
   U509 : INV_X1 port map( A => n58392, ZN => n3327);
   U510 : OAI22_X1 port map( A1 => n52436, A2 => n59173, B1 => n52873, B2 => 
                           n59124, ZN => n58393);
   U511 : INV_X1 port map( A => n58393, ZN => n3224);
   U512 : OAI22_X1 port map( A1 => n52446, A2 => n58910, B1 => n52777, B2 => 
                           n58978, ZN => n58394);
   U513 : INV_X1 port map( A => n58394, ZN => n3389);
   U514 : OAI22_X1 port map( A1 => n52469, A2 => n59209, B1 => n52938, B2 => 
                           n58996, ZN => n58395);
   U515 : INV_X1 port map( A => n58395, ZN => n3553);
   U516 : OAI22_X1 port map( A1 => n52451, A2 => n58910, B1 => n52784, B2 => 
                           n58999, ZN => n58396);
   U517 : INV_X1 port map( A => n58396, ZN => n3391);
   U518 : OAI22_X1 port map( A1 => n52459, A2 => n58781, B1 => n52942, B2 => 
                           n58993, ZN => n58397);
   U519 : INV_X1 port map( A => n58397, ZN => n3072);
   U520 : OAI22_X1 port map( A1 => n52469, A2 => n58826, B1 => n52940, B2 => 
                           n58996, ZN => n58398);
   U521 : INV_X1 port map( A => n58398, ZN => n3460);
   U522 : OAI22_X1 port map( A1 => n52436, A2 => n58781, B1 => n52848, B2 => 
                           n59124, ZN => n58399);
   U523 : INV_X1 port map( A => n58399, ZN => n3071);
   U524 : OAI22_X1 port map( A1 => n52436, A2 => n58730, B1 => n52846, B2 => 
                           n59124, ZN => n58400);
   U525 : INV_X1 port map( A => n58400, ZN => n3007);
   U526 : OAI22_X1 port map( A1 => n52436, A2 => n58800, B1 => n52950, B2 => 
                           n59124, ZN => n58401);
   U527 : INV_X1 port map( A => n58401, ZN => n2913);
   U528 : OAI22_X1 port map( A1 => n52436, A2 => n59209, B1 => n52939, B2 => 
                           n59124, ZN => n58402);
   U529 : INV_X1 port map( A => n58402, ZN => n3554);
   U530 : OAI22_X1 port map( A1 => n52478, A2 => n58800, B1 => n52864, B2 => 
                           n58980, ZN => n58403);
   U531 : INV_X1 port map( A => n58403, ZN => n2910);
   U532 : OAI22_X1 port map( A1 => n52469, A2 => n58800, B1 => n52865, B2 => 
                           n58996, ZN => n58404);
   U533 : INV_X1 port map( A => n58404, ZN => n2911);
   U534 : OAI22_X1 port map( A1 => n52459, A2 => n58721, B1 => n52943, B2 => 
                           n58993, ZN => n58405);
   U535 : INV_X1 port map( A => n58405, ZN => n2876);
   U536 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52468, ZN => n59082);
   U537 : OAI22_X1 port map( A1 => n52468, A2 => n58910, B1 => n52968, B2 => 
                           n59082, ZN => n58406);
   U538 : INV_X1 port map( A => n58406, ZN => n3396);
   U539 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52473, ZN => n59130);
   U540 : OAI22_X1 port map( A1 => n52473, A2 => n59173, B1 => n52894, B2 => 
                           n59130, ZN => n58407);
   U541 : INV_X1 port map( A => n58407, ZN => n3227);
   U542 : OAI22_X1 port map( A1 => n52468, A2 => n59169, B1 => n52913, B2 => 
                           n59082, ZN => n58408);
   U543 : INV_X1 port map( A => n58408, ZN => n3488);
   U544 : OAI22_X1 port map( A1 => n52468, A2 => n58730, B1 => n52908, B2 => 
                           n59082, ZN => n58409);
   U545 : INV_X1 port map( A => n58409, ZN => n3009);
   U546 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52477, ZN => n59126);
   U547 : OAI22_X1 port map( A1 => n52477, A2 => n58730, B1 => n52900, B2 => 
                           n59126, ZN => n58410);
   U548 : INV_X1 port map( A => n58410, ZN => n3008);
   U549 : OAI22_X1 port map( A1 => n52473, A2 => n58616, B1 => n52899, B2 => 
                           n59130, ZN => n58411);
   U550 : INV_X1 port map( A => n58411, ZN => n2983);
   U551 : OAI22_X1 port map( A1 => n52468, A2 => n59173, B1 => n52896, B2 => 
                           n59082, ZN => n58412);
   U552 : INV_X1 port map( A => n58412, ZN => n3228);
   U553 : OAI22_X1 port map( A1 => n52468, A2 => n58725, B1 => n52961, B2 => 
                           n59082, ZN => n58413);
   U554 : INV_X1 port map( A => n58413, ZN => n2854);
   U555 : OAI22_X1 port map( A1 => n52473, A2 => n58819, B1 => n52960, B2 => 
                           n59130, ZN => n58414);
   U556 : INV_X1 port map( A => n58414, ZN => n3363);
   U557 : OAI22_X1 port map( A1 => n52468, A2 => n58819, B1 => n52958, B2 => 
                           n59082, ZN => n58415);
   U558 : INV_X1 port map( A => n58415, ZN => n3361);
   U559 : OAI22_X1 port map( A1 => n52468, A2 => n58781, B1 => n52956, B2 => 
                           n59082, ZN => n58416);
   U560 : INV_X1 port map( A => n58416, ZN => n3073);
   U561 : OAI22_X1 port map( A1 => n52473, A2 => n58721, B1 => n52952, B2 => 
                           n59130, ZN => n58417);
   U562 : INV_X1 port map( A => n58417, ZN => n2878);
   U563 : OAI22_X1 port map( A1 => n52477, A2 => n58721, B1 => n52951, B2 => 
                           n59126, ZN => n58418);
   U564 : INV_X1 port map( A => n58418, ZN => n2877);
   U565 : OAI22_X1 port map( A1 => n52468, A2 => n58913, B1 => n52948, B2 => 
                           n59082, ZN => n58419);
   U566 : INV_X1 port map( A => n58419, ZN => n2976);
   U567 : OAI22_X1 port map( A1 => n52477, A2 => n58793, B1 => n52944, B2 => 
                           n59126, ZN => n58420);
   U568 : INV_X1 port map( A => n58420, ZN => n2941);
   U569 : OAI22_X1 port map( A1 => n52473, A2 => n58826, B1 => n52937, B2 => 
                           n59130, ZN => n58421);
   U570 : INV_X1 port map( A => n58421, ZN => n3459);
   U571 : OAI22_X1 port map( A1 => n52477, A2 => n58910, B1 => n52936, B2 => 
                           n59126, ZN => n58422);
   U572 : INV_X1 port map( A => n58422, ZN => n3392);
   U573 : OAI22_X1 port map( A1 => n52477, A2 => n58826, B1 => n52934, B2 => 
                           n59126, ZN => n58423);
   U574 : INV_X1 port map( A => n58423, ZN => n3458);
   U575 : OAI22_X1 port map( A1 => n52473, A2 => n58741, B1 => n52930, B2 => 
                           n59130, ZN => n58424);
   U576 : INV_X1 port map( A => n58424, ZN => n2814);
   U577 : OAI22_X1 port map( A1 => n52477, A2 => n59169, B1 => n52929, B2 => 
                           n59126, ZN => n58425);
   U578 : INV_X1 port map( A => n58425, ZN => n3491);
   U579 : OAI22_X1 port map( A1 => n52468, A2 => n58736, B1 => n52802, B2 => 
                           n59082, ZN => n58426);
   U580 : INV_X1 port map( A => n58426, ZN => n3174);
   U581 : OAI22_X1 port map( A1 => n52473, A2 => n59213, B1 => n52805, B2 => 
                           n59130, ZN => n58427);
   U582 : INV_X1 port map( A => n58427, ZN => n3200);
   U583 : OAI22_X1 port map( A1 => n52477, A2 => n58736, B1 => n52806, B2 => 
                           n59126, ZN => n58428);
   U584 : INV_X1 port map( A => n58428, ZN => n3176);
   U585 : OAI22_X1 port map( A1 => n52468, A2 => n58761, B1 => n52810, B2 => 
                           n59082, ZN => n58429);
   U586 : INV_X1 port map( A => n58429, ZN => n3166);
   U587 : OAI22_X1 port map( A1 => n52468, A2 => n58783, B1 => n52834, B2 => 
                           n59082, ZN => n58430);
   U588 : INV_X1 port map( A => n58430, ZN => n3261);
   U589 : OAI22_X1 port map( A1 => n52473, A2 => n58783, B1 => n52835, B2 => 
                           n59130, ZN => n58431);
   U590 : INV_X1 port map( A => n58431, ZN => n3262);
   U591 : OAI22_X1 port map( A1 => n52473, A2 => n58811, B1 => n52926, B2 => 
                           n59130, ZN => n58432);
   U592 : INV_X1 port map( A => n58432, ZN => n3427);
   U593 : OAI22_X1 port map( A1 => n52477, A2 => n58811, B1 => n52925, B2 => 
                           n59126, ZN => n58433);
   U594 : INV_X1 port map( A => n58433, ZN => n3426);
   U595 : OAI22_X1 port map( A1 => n52473, A2 => n59169, B1 => n52924, B2 => 
                           n59130, ZN => n58434);
   U596 : INV_X1 port map( A => n58434, ZN => n3490);
   U597 : OAI22_X1 port map( A1 => n52468, A2 => n58745, B1 => n52816, B2 => 
                           n59082, ZN => n58435);
   U598 : INV_X1 port map( A => n58435, ZN => n3110);
   U599 : OAI22_X1 port map( A1 => n52473, A2 => n58910, B1 => n52963, B2 => 
                           n59130, ZN => n58436);
   U600 : INV_X1 port map( A => n58436, ZN => n3395);
   U601 : OAI22_X1 port map( A1 => n52473, A2 => n58745, B1 => n52817, B2 => 
                           n59130, ZN => n58437);
   U602 : INV_X1 port map( A => n58437, ZN => n3111);
   U603 : OAI22_X1 port map( A1 => n52477, A2 => n58761, B1 => n53357, B2 => 
                           n59126, ZN => n58438);
   U604 : INV_X1 port map( A => n58438, ZN => n3150);
   U605 : OAI22_X1 port map( A1 => n52473, A2 => n58759, B1 => n53375, B2 => 
                           n59130, ZN => n58439);
   U606 : INV_X1 port map( A => n58439, ZN => n2831);
   U607 : OAI22_X1 port map( A1 => n52477, A2 => n58717, B1 => n52818, B2 => 
                           n59126, ZN => n58440);
   U608 : INV_X1 port map( A => n58440, ZN => n3136);
   U609 : OAI22_X1 port map( A1 => n52468, A2 => n59166, B1 => n52887, B2 => 
                           n59082, ZN => n58441);
   U610 : INV_X1 port map( A => n58441, ZN => n3329);
   U611 : OAI22_X1 port map( A1 => n52468, A2 => n58741, B1 => n52859, B2 => 
                           n59082, ZN => n58442);
   U612 : INV_X1 port map( A => n58442, ZN => n2813);
   U613 : OAI22_X1 port map( A1 => n52477, A2 => n59166, B1 => n52874, B2 => 
                           n59126, ZN => n58443);
   U614 : INV_X1 port map( A => n58443, ZN => n3328);
   U615 : OAI22_X1 port map( A1 => n52468, A2 => n58759, B1 => n53370, B2 => 
                           n59082, ZN => n58444);
   U616 : INV_X1 port map( A => n58444, ZN => n2830);
   U617 : OAI22_X1 port map( A1 => n52477, A2 => n58741, B1 => n53390, B2 => 
                           n59126, ZN => n58445);
   U618 : INV_X1 port map( A => n58445, ZN => n2800);
   U619 : OAI22_X1 port map( A1 => n52468, A2 => n58813, B1 => n52919, B2 => 
                           n59082, ZN => n58446);
   U620 : INV_X1 port map( A => n58446, ZN => n3524);
   U621 : OAI22_X1 port map( A1 => n52477, A2 => n58783, B1 => n52833, B2 => 
                           n59126, ZN => n58447);
   U622 : INV_X1 port map( A => n58447, ZN => n3260);
   U623 : OAI22_X1 port map( A1 => n52468, A2 => n58811, B1 => n52921, B2 => 
                           n59082, ZN => n58448);
   U624 : INV_X1 port map( A => n58448, ZN => n3425);
   U625 : OAI22_X1 port map( A1 => n52477, A2 => n58789, B1 => n52824, B2 => 
                           n59126, ZN => n58449);
   U626 : INV_X1 port map( A => n58449, ZN => n3104);
   U627 : OAI22_X1 port map( A1 => n52477, A2 => n59173, B1 => n52889, B2 => 
                           n59126, ZN => n58450);
   U628 : INV_X1 port map( A => n58450, ZN => n3225);
   U629 : OAI22_X1 port map( A1 => n52477, A2 => n58813, B1 => n52916, B2 => 
                           n59126, ZN => n58451);
   U630 : INV_X1 port map( A => n58451, ZN => n3521);
   U631 : OAI22_X1 port map( A1 => n52473, A2 => n58813, B1 => n52917, B2 => 
                           n59130, ZN => n58452);
   U632 : INV_X1 port map( A => n58452, ZN => n3522);
   U633 : OAI22_X1 port map( A1 => n52473, A2 => n58800, B1 => n52861, B2 => 
                           n59130, ZN => n58453);
   U634 : INV_X1 port map( A => n58453, ZN => n2909);
   U635 : OAI22_X1 port map( A1 => n52468, A2 => n58915, B1 => n52830, B2 => 
                           n59082, ZN => n58454);
   U636 : INV_X1 port map( A => n58454, ZN => n3297);
   U637 : OAI22_X1 port map( A1 => n52477, A2 => n58759, B1 => n52868, B2 => 
                           n59126, ZN => n58455);
   U638 : INV_X1 port map( A => n58455, ZN => n2848);
   U639 : OAI22_X1 port map( A1 => n52468, A2 => n58800, B1 => n52871, B2 => 
                           n59082, ZN => n58456);
   U640 : INV_X1 port map( A => n58456, ZN => n2912);
   U641 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53606, ZN => n59112);
   U642 : OAI22_X1 port map( A1 => n52456, A2 => n59112, B1 => n53271, B2 => 
                           n58982, ZN => n58457);
   U643 : INV_X1 port map( A => n58457, ZN => n3023);
   U644 : OAI22_X1 port map( A1 => n52449, A2 => n59112, B1 => n53251, B2 => 
                           n58976, ZN => n58458);
   U645 : INV_X1 port map( A => n58458, ZN => n3022);
   U646 : OAI22_X1 port map( A1 => n52458, A2 => n59112, B1 => n52522, B2 => 
                           n59006, ZN => n58459);
   U647 : INV_X1 port map( A => n58459, ZN => n3025);
   U648 : OAI22_X1 port map( A1 => n52478, A2 => n59112, B1 => n52906, B2 => 
                           n58980, ZN => n58460);
   U649 : INV_X1 port map( A => n58460, ZN => n3041);
   U650 : OAI22_X1 port map( A1 => n52455, A2 => n59112, B1 => n52716, B2 => 
                           n58985, ZN => n58461);
   U651 : INV_X1 port map( A => n58461, ZN => n3035);
   U652 : OAI22_X1 port map( A1 => n52451, A2 => n59112, B1 => n52675, B2 => 
                           n58999, ZN => n58462);
   U653 : INV_X1 port map( A => n58462, ZN => n3031);
   U654 : OAI22_X1 port map( A1 => n52459, A2 => n59112, B1 => n52797, B2 => 
                           n58993, ZN => n58463);
   U655 : INV_X1 port map( A => n58463, ZN => n3037);
   U656 : OAI22_X1 port map( A1 => n52446, A2 => n59112, B1 => n52700, B2 => 
                           n58978, ZN => n58464);
   U657 : INV_X1 port map( A => n58464, ZN => n3033);
   U658 : OAI22_X1 port map( A1 => n52469, A2 => n59112, B1 => n52799, B2 => 
                           n58996, ZN => n58465);
   U659 : INV_X1 port map( A => n58465, ZN => n3039);
   U660 : OAI22_X1 port map( A1 => n52468, A2 => n59112, B1 => n52798, B2 => 
                           n59082, ZN => n58466);
   U661 : INV_X1 port map( A => n58466, ZN => n3038);
   U662 : OAI22_X1 port map( A1 => n52445, A2 => n59112, B1 => n53057, B2 => 
                           n58967, ZN => n58467);
   U663 : INV_X1 port map( A => n58467, ZN => n3045);
   U664 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52440, ZN => n59152);
   U665 : OAI22_X1 port map( A1 => n52440, A2 => n59173, B1 => n53291, B2 => 
                           n59152, ZN => n58468);
   U666 : INV_X1 port map( A => n58468, ZN => n3214);
   U667 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52443, ZN => n59158);
   U668 : OAI22_X1 port map( A1 => n52443, A2 => n59173, B1 => n53308, B2 => 
                           n59158, ZN => n58469);
   U669 : INV_X1 port map( A => n58469, ZN => n3216);
   U670 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52437, ZN => n59150);
   U671 : OAI22_X1 port map( A1 => n52437, A2 => n58783, B1 => n53325, B2 => 
                           n59150, ZN => n58470);
   U672 : INV_X1 port map( A => n58470, ZN => n3246);
   U673 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52447, ZN => n59144);
   U674 : OAI22_X1 port map( A1 => n52447, A2 => n59173, B1 => n52758, B2 => 
                           n59144, ZN => n58471);
   U675 : INV_X1 port map( A => n58471, ZN => n3222);
   U676 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52448, ZN => n59171);
   U677 : OAI22_X1 port map( A1 => n52448, A2 => n58819, B1 => n52981, B2 => 
                           n59171, ZN => n58472);
   U678 : INV_X1 port map( A => n58472, ZN => n3365);
   U679 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52450, ZN => n59175);
   U680 : OAI22_X1 port map( A1 => n52450, A2 => n58811, B1 => n52984, B2 => 
                           n59175, ZN => n58473);
   U681 : INV_X1 port map( A => n58473, ZN => n3429);
   U682 : OAI22_X1 port map( A1 => n52450, A2 => n58826, B1 => n52985, B2 => 
                           n59175, ZN => n58474);
   U683 : INV_X1 port map( A => n58474, ZN => n3461);
   U684 : OAI22_X1 port map( A1 => n52450, A2 => n58910, B1 => n52995, B2 => 
                           n59175, ZN => n58475);
   U685 : INV_X1 port map( A => n58475, ZN => n3397);
   U686 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52467, ZN => n59212);
   U687 : OAI22_X1 port map( A1 => n52467, A2 => n58759, B1 => n53004, B2 => 
                           n59212, ZN => n58476);
   U688 : INV_X1 port map( A => n58476, ZN => n2852);
   U689 : OAI22_X1 port map( A1 => n52467, A2 => n58741, B1 => n53006, B2 => 
                           n59212, ZN => n58477);
   U690 : INV_X1 port map( A => n58477, ZN => n2817);
   U691 : OAI22_X1 port map( A1 => n52448, A2 => n58813, B1 => n53011, B2 => 
                           n59171, ZN => n58478);
   U692 : INV_X1 port map( A => n58478, ZN => n3525);
   U693 : OAI22_X1 port map( A1 => n52467, A2 => n58800, B1 => n53018, B2 => 
                           n59212, ZN => n58479);
   U694 : INV_X1 port map( A => n58479, ZN => n2915);
   U695 : OAI22_X1 port map( A1 => n52467, A2 => n59166, B1 => n53019, B2 => 
                           n59212, ZN => n58480);
   U696 : INV_X1 port map( A => n58480, ZN => n3310);
   U697 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52442, ZN => n59168);
   U698 : OAI22_X1 port map( A1 => n52442, A2 => n58811, B1 => n53024, B2 => 
                           n59168, ZN => n58481);
   U699 : INV_X1 port map( A => n58481, ZN => n3406);
   U700 : OAI22_X1 port map( A1 => n52448, A2 => n58826, B1 => n53031, B2 => 
                           n59171, ZN => n58482);
   U701 : INV_X1 port map( A => n58482, ZN => n3438);
   U702 : OAI22_X1 port map( A1 => n52450, A2 => n59169, B1 => n53032, B2 => 
                           n59175, ZN => n58483);
   U703 : INV_X1 port map( A => n58483, ZN => n3470);
   U704 : OAI22_X1 port map( A1 => n52450, A2 => n58813, B1 => n53033, B2 => 
                           n59175, ZN => n58484);
   U705 : INV_X1 port map( A => n58484, ZN => n3502);
   U706 : OAI22_X1 port map( A1 => n52450, A2 => n58721, B1 => n53071, B2 => 
                           n59175, ZN => n58485);
   U707 : INV_X1 port map( A => n58485, ZN => n2880);
   U708 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52441, ZN => n59161);
   U709 : OAI22_X1 port map( A1 => n52441, A2 => n58721, B1 => n53074, B2 => 
                           n59161, ZN => n58486);
   U710 : INV_X1 port map( A => n58486, ZN => n2882);
   U711 : OAI22_X1 port map( A1 => n52442, A2 => n58721, B1 => n53075, B2 => 
                           n59168, ZN => n58487);
   U712 : INV_X1 port map( A => n58487, ZN => n2883);
   U713 : OAI22_X1 port map( A1 => n52450, A2 => n58741, B1 => n53093, B2 => 
                           n59175, ZN => n58488);
   U714 : INV_X1 port map( A => n58488, ZN => n2818);
   U715 : OAI22_X1 port map( A1 => n52442, A2 => n58736, B1 => n53097, B2 => 
                           n59168, ZN => n58489);
   U716 : INV_X1 port map( A => n58489, ZN => n3180);
   U717 : OAI22_X1 port map( A1 => n52467, A2 => n58730, B1 => n53104, B2 => 
                           n59212, ZN => n58490);
   U718 : INV_X1 port map( A => n58490, ZN => n2990);
   U719 : OAI22_X1 port map( A1 => n52467, A2 => n59169, B1 => n53108, B2 => 
                           n59212, ZN => n58491);
   U720 : INV_X1 port map( A => n58491, ZN => n3472);
   U721 : OAI22_X1 port map( A1 => n52441, A2 => n58761, B1 => n53111, B2 => 
                           n59161, ZN => n58492);
   U722 : INV_X1 port map( A => n58492, ZN => n3172);
   U723 : OAI22_X1 port map( A1 => n52442, A2 => n58761, B1 => n53112, B2 => 
                           n59168, ZN => n58493);
   U724 : INV_X1 port map( A => n58493, ZN => n3173);
   U725 : OAI22_X1 port map( A1 => n52441, A2 => n58745, B1 => n53115, B2 => 
                           n59161, ZN => n58494);
   U726 : INV_X1 port map( A => n58494, ZN => n3115);
   U727 : OAI22_X1 port map( A1 => n52442, A2 => n58745, B1 => n53117, B2 => 
                           n59168, ZN => n58495);
   U728 : INV_X1 port map( A => n58495, ZN => n3116);
   U729 : OAI22_X1 port map( A1 => n52442, A2 => n58616, B1 => n53066, B2 => 
                           n59168, ZN => n58496);
   U730 : INV_X1 port map( A => n58496, ZN => n2987);
   U731 : OAI22_X1 port map( A1 => n52441, A2 => n58616, B1 => n53065, B2 => 
                           n59161, ZN => n58497);
   U732 : INV_X1 port map( A => n58497, ZN => n2986);
   U733 : OAI22_X1 port map( A1 => n52450, A2 => n58717, B1 => n53130, B2 => 
                           n59175, ZN => n58498);
   U734 : INV_X1 port map( A => n58498, ZN => n3118);
   U735 : OAI22_X1 port map( A1 => n52448, A2 => n59173, B1 => n53137, B2 => 
                           n59171, ZN => n58499);
   U736 : INV_X1 port map( A => n58499, ZN => n3235);
   U737 : OAI22_X1 port map( A1 => n52467, A2 => n58811, B1 => n53138, B2 => 
                           n59212, ZN => n58500);
   U738 : INV_X1 port map( A => n58500, ZN => n3408);
   U739 : OAI22_X1 port map( A1 => n52441, A2 => n58736, B1 => n53096, B2 => 
                           n59161, ZN => n58501);
   U740 : INV_X1 port map( A => n58501, ZN => n3179);
   U741 : OAI22_X1 port map( A1 => n52441, A2 => n58915, B1 => n53143, B2 => 
                           n59161, ZN => n58502);
   U742 : INV_X1 port map( A => n58502, ZN => n3278);
   U743 : OAI22_X1 port map( A1 => n52467, A2 => n58781, B1 => n53145, B2 => 
                           n59212, ZN => n58503);
   U744 : INV_X1 port map( A => n58503, ZN => n3054);
   U745 : OAI22_X1 port map( A1 => n52467, A2 => n58915, B1 => n53146, B2 => 
                           n59212, ZN => n58504);
   U746 : INV_X1 port map( A => n58504, ZN => n3279);
   U747 : OAI22_X1 port map( A1 => n52442, A2 => n58741, B1 => n53147, B2 => 
                           n59168, ZN => n58505);
   U748 : INV_X1 port map( A => n58505, ZN => n2820);
   U749 : OAI22_X1 port map( A1 => n52450, A2 => n58730, B1 => n53062, B2 => 
                           n59175, ZN => n58506);
   U750 : INV_X1 port map( A => n58506, ZN => n3012);
   U751 : OAI22_X1 port map( A1 => n52467, A2 => n58819, B1 => n53149, B2 => 
                           n59212, ZN => n58507);
   U752 : INV_X1 port map( A => n58507, ZN => n3344);
   U753 : OAI22_X1 port map( A1 => n52448, A2 => n58915, B1 => n53151, B2 => 
                           n59171, ZN => n58508);
   U754 : INV_X1 port map( A => n58508, ZN => n3280);
   U755 : OAI22_X1 port map( A1 => n52450, A2 => n58793, B1 => n53152, B2 => 
                           n59175, ZN => n58509);
   U756 : INV_X1 port map( A => n58509, ZN => n2926);
   U757 : OAI22_X1 port map( A1 => n52442, A2 => n58793, B1 => n53157, B2 => 
                           n59168, ZN => n58510);
   U758 : INV_X1 port map( A => n58510, ZN => n2945);
   U759 : OAI22_X1 port map( A1 => n52467, A2 => n58717, B1 => n53158, B2 => 
                           n59212, ZN => n58511);
   U760 : INV_X1 port map( A => n58511, ZN => n3119);
   U761 : OAI22_X1 port map( A1 => n52448, A2 => n58730, B1 => n53056, B2 => 
                           n59171, ZN => n58512);
   U762 : INV_X1 port map( A => n58512, ZN => n3011);
   U763 : OAI22_X1 port map( A1 => n52441, A2 => n58793, B1 => n53159, B2 => 
                           n59161, ZN => n58513);
   U764 : INV_X1 port map( A => n58513, ZN => n2946);
   U765 : OAI22_X1 port map( A1 => n52442, A2 => n59112, B1 => n53055, B2 => 
                           n59168, ZN => n58514);
   U766 : INV_X1 port map( A => n58514, ZN => n3044);
   U767 : OAI22_X1 port map( A1 => n52441, A2 => n58741, B1 => n53161, B2 => 
                           n59161, ZN => n58515);
   U768 : INV_X1 port map( A => n58515, ZN => n2821);
   U769 : OAI22_X1 port map( A1 => n52467, A2 => n58910, B1 => n53162, B2 => 
                           n59212, ZN => n58516);
   U770 : INV_X1 port map( A => n58516, ZN => n3376);
   U771 : OAI22_X1 port map( A1 => n52441, A2 => n58789, B1 => n53167, B2 => 
                           n59161, ZN => n58517);
   U772 : INV_X1 port map( A => n58517, ZN => n3086);
   U773 : OAI22_X1 port map( A1 => n52441, A2 => n59112, B1 => n53054, B2 => 
                           n59161, ZN => n58518);
   U774 : INV_X1 port map( A => n58518, ZN => n3043);
   U775 : OAI22_X1 port map( A1 => n52467, A2 => n58725, B1 => n53168, B2 => 
                           n59212, ZN => n58519);
   U776 : INV_X1 port map( A => n58519, ZN => n2857);
   U777 : OAI22_X1 port map( A1 => n52467, A2 => n58793, B1 => n53170, B2 => 
                           n59212, ZN => n58520);
   U778 : INV_X1 port map( A => n58520, ZN => n2947);
   U779 : OAI22_X1 port map( A1 => n52467, A2 => n58826, B1 => n53177, B2 => 
                           n59212, ZN => n58521);
   U780 : INV_X1 port map( A => n58521, ZN => n3440);
   U781 : OAI22_X1 port map( A1 => n52448, A2 => n58655, B1 => n53053, B2 => 
                           n59171, ZN => n58522);
   U782 : INV_X1 port map( A => n58522, ZN => n2792);
   U783 : OAI22_X1 port map( A1 => n52448, A2 => n58759, B1 => n53052, B2 => 
                           n59171, ZN => n58523);
   U784 : INV_X1 port map( A => n58523, ZN => n2853);
   U785 : OAI22_X1 port map( A1 => n52448, A2 => n58725, B1 => n53051, B2 => 
                           n59171, ZN => n58524);
   U786 : INV_X1 port map( A => n58524, ZN => n2855);
   U787 : OAI22_X1 port map( A1 => n52450, A2 => n58783, B1 => n53125, B2 => 
                           n59175, ZN => n58525);
   U788 : INV_X1 port map( A => n58525, ZN => n3269);
   U789 : OAI22_X1 port map( A1 => n52467, A2 => n59209, B1 => n53187, B2 => 
                           n59212, ZN => n58526);
   U790 : INV_X1 port map( A => n58526, ZN => n3534);
   U791 : OAI22_X1 port map( A1 => n52442, A2 => n59209, B1 => n53188, B2 => 
                           n59168, ZN => n58527);
   U792 : INV_X1 port map( A => n58527, ZN => n3535);
   U793 : OAI22_X1 port map( A1 => n52450, A2 => n59173, B1 => n53126, B2 => 
                           n59175, ZN => n58528);
   U794 : INV_X1 port map( A => n58528, ZN => n3234);
   U795 : OAI22_X1 port map( A1 => n52440, A2 => n58725, B1 => n53200, B2 => 
                           n59152, ZN => n58529);
   U796 : INV_X1 port map( A => n58529, ZN => n2858);
   U797 : OAI22_X1 port map( A1 => n52448, A2 => n58800, B1 => n53050, B2 => 
                           n59171, ZN => n58530);
   U798 : INV_X1 port map( A => n58530, ZN => n2916);
   U799 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52457, ZN => n59156);
   U800 : OAI22_X1 port map( A1 => n52457, A2 => n58800, B1 => n53203, B2 => 
                           n59156, ZN => n58531);
   U801 : INV_X1 port map( A => n58531, ZN => n2894);
   U802 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52435, ZN => n59164);
   U803 : OAI22_X1 port map( A1 => n52435, A2 => n58761, B1 => n53394, B2 => 
                           n59164, ZN => n58532);
   U804 : INV_X1 port map( A => n58532, ZN => n3151);
   U805 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52439, ZN => n59154);
   U806 : OAI22_X1 port map( A1 => n52439, A2 => n58793, B1 => n53211, B2 => 
                           n59154, ZN => n58533);
   U807 : INV_X1 port map( A => n58533, ZN => n2949);
   U808 : OAI22_X1 port map( A1 => n52435, A2 => n58789, B1 => n53388, B2 => 
                           n59164, ZN => n58534);
   U809 : INV_X1 port map( A => n58534, ZN => n3088);
   U810 : OAI22_X1 port map( A1 => n52467, A2 => n58813, B1 => n53127, B2 => 
                           n59212, ZN => n58535);
   U811 : INV_X1 port map( A => n58535, ZN => n3504);
   U812 : OAI22_X1 port map( A1 => n52448, A2 => n58793, B1 => n53049, B2 => 
                           n59171, ZN => n58536);
   U813 : INV_X1 port map( A => n58536, ZN => n2928);
   U814 : OAI22_X1 port map( A1 => n52440, A2 => n58655, B1 => n53232, B2 => 
                           n59152, ZN => n58537);
   U815 : INV_X1 port map( A => n58537, ZN => n2795);
   U816 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52453, ZN => n59148);
   U817 : OAI22_X1 port map( A1 => n52453, A2 => n58913, B1 => n53350, B2 => 
                           n59148, ZN => n58538);
   U818 : INV_X1 port map( A => n58538, ZN => n2960);
   U819 : OAI22_X1 port map( A1 => n52443, A2 => n58655, B1 => n53349, B2 => 
                           n59158, ZN => n58539);
   U820 : INV_X1 port map( A => n58539, ZN => n2797);
   U821 : OAI22_X1 port map( A1 => n52448, A2 => n58913, B1 => n53048, B2 => 
                           n59171, ZN => n58540);
   U822 : INV_X1 port map( A => n58540, ZN => n2979);
   U823 : OAI22_X1 port map( A1 => n52448, A2 => n58781, B1 => n53047, B2 => 
                           n59171, ZN => n58541);
   U824 : INV_X1 port map( A => n58541, ZN => n3076);
   U825 : OAI22_X1 port map( A1 => n52448, A2 => n59112, B1 => n53046, B2 => 
                           n59171, ZN => n58542);
   U826 : INV_X1 port map( A => n58542, ZN => n3042);
   U827 : OAI22_X1 port map( A1 => n52448, A2 => n58717, B1 => n53045, B2 => 
                           n59171, ZN => n58543);
   U828 : INV_X1 port map( A => n58543, ZN => n3141);
   U829 : OAI22_X1 port map( A1 => n52453, A2 => n59173, B1 => n53244, B2 => 
                           n59148, ZN => n58544);
   U830 : INV_X1 port map( A => n58544, ZN => n3237);
   U831 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52463, ZN => n59146);
   U832 : OAI22_X1 port map( A1 => n52463, A2 => n58721, B1 => n53344, B2 => 
                           n59146, ZN => n58545);
   U833 : INV_X1 port map( A => n58545, ZN => n2863);
   U834 : OAI22_X1 port map( A1 => n52448, A2 => n58789, B1 => n53044, B2 => 
                           n59171, ZN => n58546);
   U835 : INV_X1 port map( A => n58546, ZN => n3108);
   U836 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52438, ZN => n59183);
   U837 : OAI22_X1 port map( A1 => n52438, A2 => n58655, B1 => n53247, B2 => 
                           n59183, ZN => n58547);
   U838 : INV_X1 port map( A => n58547, ZN => n2796);
   U839 : OAI22_X1 port map( A1 => n52437, A2 => n59112, B1 => n53343, B2 => 
                           n59150, ZN => n58548);
   U840 : INV_X1 port map( A => n58548, ZN => n3024);
   U841 : OAI22_X1 port map( A1 => n52457, A2 => n58725, B1 => n53249, B2 => 
                           n59156, ZN => n58549);
   U842 : INV_X1 port map( A => n58549, ZN => n2859);
   U843 : OAI22_X1 port map( A1 => n52437, A2 => n58800, B1 => n53255, B2 => 
                           n59150, ZN => n58550);
   U844 : INV_X1 port map( A => n58550, ZN => n2896);
   U845 : OAI22_X1 port map( A1 => n52447, A2 => n58783, B1 => n53331, B2 => 
                           n59144, ZN => n58551);
   U846 : INV_X1 port map( A => n58551, ZN => n3247);
   U847 : OAI22_X1 port map( A1 => n52467, A2 => n59173, B1 => n53037, B2 => 
                           n59212, ZN => n58552);
   U848 : INV_X1 port map( A => n58552, ZN => n3231);
   U849 : OAI22_X1 port map( A1 => n52438, A2 => n58781, B1 => n53329, B2 => 
                           n59183, ZN => n58553);
   U850 : INV_X1 port map( A => n58553, ZN => n3055);
   U851 : OAI22_X1 port map( A1 => n52447, A2 => n58913, B1 => n53326, B2 => 
                           n59144, ZN => n58554);
   U852 : INV_X1 port map( A => n58554, ZN => n2959);
   U853 : OAI22_X1 port map( A1 => n52435, A2 => n58915, B1 => n52838, B2 => 
                           n59164, ZN => n58555);
   U854 : INV_X1 port map( A => n58555, ZN => n3299);
   U855 : OAI22_X1 port map( A1 => n52435, A2 => n58717, B1 => n52841, B2 => 
                           n59164, ZN => n58556);
   U856 : INV_X1 port map( A => n58556, ZN => n3138);
   U857 : OAI22_X1 port map( A1 => n52457, A2 => n58789, B1 => n52680, B2 => 
                           n59156, ZN => n58557);
   U858 : INV_X1 port map( A => n58557, ZN => n3099);
   U859 : OAI22_X1 port map( A1 => n52457, A2 => n58915, B1 => n52679, B2 => 
                           n59156, ZN => n58558);
   U860 : INV_X1 port map( A => n58558, ZN => n3291);
   U861 : OAI22_X1 port map( A1 => n52447, A2 => n58761, B1 => n52785, B2 => 
                           n59144, ZN => n58559);
   U862 : INV_X1 port map( A => n58559, ZN => n3165);
   U863 : OAI22_X1 port map( A1 => n52457, A2 => n58783, B1 => n52677, B2 => 
                           n59156, ZN => n58560);
   U864 : INV_X1 port map( A => n58560, ZN => n3256);
   U865 : OAI22_X1 port map( A1 => n52457, A2 => n58913, B1 => n52674, B2 => 
                           n59156, ZN => n58561);
   U866 : INV_X1 port map( A => n58561, ZN => n2969);
   U867 : OAI22_X1 port map( A1 => n52435, A2 => n59112, B1 => n52845, B2 => 
                           n59164, ZN => n58562);
   U868 : INV_X1 port map( A => n58562, ZN => n3040);
   U869 : OAI22_X1 port map( A1 => n52457, A2 => n58717, B1 => n52518, B2 => 
                           n59156, ZN => n58563);
   U870 : INV_X1 port map( A => n58563, ZN => n3122);
   U871 : OAI22_X1 port map( A1 => n52463, A2 => n58910, B1 => n52517, B2 => 
                           n59146, ZN => n58564);
   U872 : INV_X1 port map( A => n58564, ZN => n3380);
   U873 : OAI22_X1 port map( A1 => n52437, A2 => n59173, B1 => n52511, B2 => 
                           n59150, ZN => n58565);
   U874 : INV_X1 port map( A => n58565, ZN => n3217);
   U875 : OAI22_X1 port map( A1 => n52463, A2 => n58913, B1 => n52509, B2 => 
                           n59146, ZN => n58566);
   U876 : INV_X1 port map( A => n58566, ZN => n2961);
   U877 : OAI22_X1 port map( A1 => n52438, A2 => n59169, B1 => n52508, B2 => 
                           n59183, ZN => n58567);
   U878 : INV_X1 port map( A => n58567, ZN => n3476);
   U879 : OAI22_X1 port map( A1 => n52439, A2 => n58813, B1 => n52506, B2 => 
                           n59154, ZN => n58568);
   U880 : INV_X1 port map( A => n58568, ZN => n3508);
   U881 : OAI22_X1 port map( A1 => n52447, A2 => n58819, B1 => n52786, B2 => 
                           n59144, ZN => n58569);
   U882 : INV_X1 port map( A => n58569, ZN => n3357);
   U883 : OAI22_X1 port map( A1 => n52447, A2 => n58813, B1 => n52755, B2 => 
                           n59144, ZN => n58570);
   U884 : INV_X1 port map( A => n58570, ZN => n3516);
   U885 : OAI22_X1 port map( A1 => n52439, A2 => n58910, B1 => n52505, B2 => 
                           n59154, ZN => n58571);
   U886 : INV_X1 port map( A => n58571, ZN => n3379);
   U887 : OAI22_X1 port map( A1 => n52440, A2 => n58826, B1 => n52503, B2 => 
                           n59152, ZN => n58572);
   U888 : INV_X1 port map( A => n58572, ZN => n3442);
   U889 : OAI22_X1 port map( A1 => n52440, A2 => n59169, B1 => n52502, B2 => 
                           n59152, ZN => n58573);
   U890 : INV_X1 port map( A => n58573, ZN => n3475);
   U891 : OAI22_X1 port map( A1 => n52443, A2 => n58811, B1 => n52789, B2 => 
                           n59158, ZN => n58574);
   U892 : INV_X1 port map( A => n58574, ZN => n3422);
   U893 : OAI22_X1 port map( A1 => n52447, A2 => n58717, B1 => n52790, B2 => 
                           n59144, ZN => n58575);
   U894 : INV_X1 port map( A => n58575, ZN => n3134);
   U895 : OAI22_X1 port map( A1 => n52443, A2 => n58826, B1 => n52791, B2 => 
                           n59158, ZN => n58576);
   U896 : INV_X1 port map( A => n58576, ZN => n3455);
   U897 : OAI22_X1 port map( A1 => n52447, A2 => n59169, B1 => n52795, B2 => 
                           n59144, ZN => n58577);
   U898 : INV_X1 port map( A => n58577, ZN => n3487);
   U899 : OAI22_X1 port map( A1 => n52463, A2 => n58793, B1 => n52500, B2 => 
                           n59146, ZN => n58578);
   U900 : INV_X1 port map( A => n58578, ZN => n2929);
   U901 : OAI22_X1 port map( A1 => n52439, A2 => n58826, B1 => n52499, B2 => 
                           n59154, ZN => n58579);
   U902 : INV_X1 port map( A => n58579, ZN => n3441);
   U903 : OAI22_X1 port map( A1 => n52440, A2 => n58819, B1 => n52498, B2 => 
                           n59152, ZN => n58580);
   U904 : INV_X1 port map( A => n58580, ZN => n3346);
   U905 : OAI22_X1 port map( A1 => n52437, A2 => n58811, B1 => n52497, B2 => 
                           n59150, ZN => n58581);
   U906 : INV_X1 port map( A => n58581, ZN => n3412);
   U907 : OAI22_X1 port map( A1 => n52439, A2 => n59169, B1 => n52495, B2 => 
                           n59154, ZN => n58582);
   U908 : INV_X1 port map( A => n58582, ZN => n3474);
   U909 : OAI22_X1 port map( A1 => n52437, A2 => n58910, B1 => n52494, B2 => 
                           n59150, ZN => n58583);
   U910 : INV_X1 port map( A => n58583, ZN => n3378);
   U911 : OAI22_X1 port map( A1 => n52439, A2 => n58811, B1 => n52493, B2 => 
                           n59154, ZN => n58584);
   U912 : INV_X1 port map( A => n58584, ZN => n3410);
   U913 : OAI22_X1 port map( A1 => n52438, A2 => n58910, B1 => n52492, B2 => 
                           n59183, ZN => n58585);
   U914 : INV_X1 port map( A => n58585, ZN => n3377);
   U915 : OAI22_X1 port map( A1 => n52438, A2 => n58811, B1 => n52491, B2 => 
                           n59183, ZN => n58586);
   U916 : INV_X1 port map( A => n58586, ZN => n3409);
   U917 : OAI22_X1 port map( A1 => n52463, A2 => n59213, B1 => n52489, B2 => 
                           n59146, ZN => n58587);
   U918 : INV_X1 port map( A => n58587, ZN => n3185);
   U919 : OAI22_X1 port map( A1 => n52435, A2 => n59166, B1 => n52903, B2 => 
                           n59164, ZN => n58588);
   U920 : INV_X1 port map( A => n58588, ZN => n3331);
   U921 : OAI22_X1 port map( A1 => n52438, A2 => n58813, B1 => n52488, B2 => 
                           n59183, ZN => n58589);
   U922 : INV_X1 port map( A => n58589, ZN => n3506);
   U923 : OAI22_X1 port map( A1 => n52437, A2 => n59169, B1 => n52487, B2 => 
                           n59150, ZN => n58590);
   U924 : INV_X1 port map( A => n58590, ZN => n3473);
   U925 : OAI22_X1 port map( A1 => n52437, A2 => n58819, B1 => n53529, B2 => 
                           n59150, ZN => n58591);
   U926 : INV_X1 port map( A => n58591, ZN => n3345);
   U927 : OAI22_X1 port map( A1 => n52437, A2 => n58813, B1 => n52486, B2 => 
                           n59150, ZN => n58592);
   U928 : INV_X1 port map( A => n58592, ZN => n3505);
   U929 : OAI22_X1 port map( A1 => n52463, A2 => n58789, B1 => n52485, B2 => 
                           n59146, ZN => n58593);
   U930 : INV_X1 port map( A => n58593, ZN => n3089);
   U931 : OAI22_X1 port map( A1 => n52435, A2 => n59173, B1 => n52872, B2 => 
                           n59164, ZN => n58594);
   U932 : INV_X1 port map( A => n58594, ZN => n3223);
   U933 : OAI22_X1 port map( A1 => n52435, A2 => n58616, B1 => n52857, B2 => 
                           n59164, ZN => n58595);
   U934 : INV_X1 port map( A => n58595, ZN => n2982);
   U935 : OAI22_X1 port map( A1 => n52435, A2 => n58913, B1 => n52856, B2 => 
                           n59164, ZN => n58596);
   U936 : INV_X1 port map( A => n58596, ZN => n2975);
   U937 : OAI22_X1 port map( A1 => n52435, A2 => n58793, B1 => n52855, B2 => 
                           n59164, ZN => n58597);
   U938 : INV_X1 port map( A => n58597, ZN => n2940);
   U939 : OAI22_X1 port map( A1 => n52463, A2 => n58717, B1 => n52524, B2 => 
                           n59146, ZN => n58598);
   U940 : INV_X1 port map( A => n58598, ZN => n3123);
   U941 : OAI22_X1 port map( A1 => n52443, A2 => n59169, B1 => n52754, B2 => 
                           n59158, ZN => n58599);
   U942 : INV_X1 port map( A => n58599, ZN => n3483);
   U943 : OAI22_X1 port map( A1 => n52453, A2 => n59112, B1 => n52673, B2 => 
                           n59148, ZN => n58600);
   U944 : INV_X1 port map( A => n58600, ZN => n3030);
   U945 : OAI22_X1 port map( A1 => n52447, A2 => n59166, B1 => n52753, B2 => 
                           n59144, ZN => n58601);
   U946 : INV_X1 port map( A => n58601, ZN => n3324);
   U947 : OAI22_X1 port map( A1 => n52457, A2 => n59169, B1 => n52671, B2 => 
                           n59156, ZN => n58602);
   U948 : INV_X1 port map( A => n58602, ZN => n3481);
   U949 : OAI22_X1 port map( A1 => n52457, A2 => n58730, B1 => n52670, B2 => 
                           n59156, ZN => n58603);
   U950 : INV_X1 port map( A => n58603, ZN => n3005);
   U951 : OAI22_X1 port map( A1 => n52457, A2 => n58781, B1 => n52669, B2 => 
                           n59156, ZN => n58604);
   U952 : INV_X1 port map( A => n58604, ZN => n3066);
   U953 : OAI22_X1 port map( A1 => n52453, A2 => n58811, B1 => n52668, B2 => 
                           n59148, ZN => n58605);
   U954 : INV_X1 port map( A => n58605, ZN => n3418);
   U955 : OAI22_X1 port map( A1 => n52443, A2 => n58781, B1 => n52759, B2 => 
                           n59158, ZN => n58606);
   U956 : INV_X1 port map( A => n58606, ZN => n3069);
   U957 : OAI22_X1 port map( A1 => n52453, A2 => n58813, B1 => n52667, B2 => 
                           n59148, ZN => n58607);
   U958 : INV_X1 port map( A => n58607, ZN => n3514);
   U959 : OAI22_X1 port map( A1 => n52453, A2 => n58819, B1 => n52666, B2 => 
                           n59148, ZN => n58608);
   U960 : INV_X1 port map( A => n58608, ZN => n3354);
   U961 : OAI22_X1 port map( A1 => n52441, A2 => n58783, B1 => n53119, B2 => 
                           n59161, ZN => n58609);
   U962 : INV_X1 port map( A => n58609, ZN => n3267);
   U963 : OAI22_X1 port map( A1 => n52447, A2 => n58811, B1 => n52751, B2 => 
                           n59144, ZN => n58610);
   U964 : INV_X1 port map( A => n58610, ZN => n3419);
   U965 : OAI22_X1 port map( A1 => n52438, A2 => n58783, B1 => n52544, B2 => 
                           n59183, ZN => n58611);
   U966 : INV_X1 port map( A => n58611, ZN => n3250);
   U967 : OAI22_X1 port map( A1 => n52453, A2 => n59169, B1 => n52660, B2 => 
                           n59148, ZN => n58612);
   U968 : INV_X1 port map( A => n58612, ZN => n3480);
   U969 : OAI22_X1 port map( A1 => n52443, A2 => n58819, B1 => n52748, B2 => 
                           n59158, ZN => n58613);
   U970 : INV_X1 port map( A => n58613, ZN => n3355);
   U971 : OAI22_X1 port map( A1 => n52435, A2 => n58759, B1 => n52967, B2 => 
                           n59164, ZN => n58614);
   U972 : INV_X1 port map( A => n58614, ZN => n2849);
   U973 : OAI22_X1 port map( A1 => n52438, A2 => n58730, B1 => n52545, B2 => 
                           n59183, ZN => n58615);
   U974 : INV_X1 port map( A => n58615, ZN => n2994);
   U975 : OAI22_X1 port map( A1 => n52453, A2 => n58616, B1 => n52649, B2 => 
                           n59148, ZN => n58617);
   U976 : INV_X1 port map( A => n58617, ZN => n3002);
   U977 : OAI22_X1 port map( A1 => n52443, A2 => n58730, B1 => n52646, B2 => 
                           n59158, ZN => n58618);
   U978 : INV_X1 port map( A => n58618, ZN => n3001);
   U979 : OAI22_X1 port map( A1 => n52453, A2 => n59209, B1 => n52644, B2 => 
                           n59148, ZN => n58619);
   U980 : INV_X1 port map( A => n58619, ZN => n3543);
   U981 : OAI22_X1 port map( A1 => n52443, A2 => n59209, B1 => n52643, B2 => 
                           n59158, ZN => n58620);
   U982 : INV_X1 port map( A => n58620, ZN => n3542);
   U983 : OAI22_X1 port map( A1 => n52453, A2 => n58759, B1 => n52746, B2 => 
                           n59148, ZN => n58621);
   U984 : INV_X1 port map( A => n58621, ZN => n2847);
   U985 : OAI22_X1 port map( A1 => n52457, A2 => n58826, B1 => n52640, B2 => 
                           n59156, ZN => n58622);
   U986 : INV_X1 port map( A => n58622, ZN => n3448);
   U987 : OAI22_X1 port map( A1 => n52447, A2 => n58781, B1 => n52745, B2 => 
                           n59144, ZN => n58623);
   U988 : INV_X1 port map( A => n58623, ZN => n3067);
   U989 : OAI22_X1 port map( A1 => n52443, A2 => n58783, B1 => n52744, B2 => 
                           n59158, ZN => n58624);
   U990 : INV_X1 port map( A => n58624, ZN => n3258);
   U991 : OAI22_X1 port map( A1 => n52438, A2 => n59213, B1 => n52543, B2 => 
                           n59183, ZN => n58625);
   U992 : INV_X1 port map( A => n58625, ZN => n3189);
   U993 : OAI22_X1 port map( A1 => n52457, A2 => n58813, B1 => n52633, B2 => 
                           n59156, ZN => n58626);
   U994 : INV_X1 port map( A => n58626, ZN => n3511);
   U995 : OAI22_X1 port map( A1 => n52437, A2 => n58915, B1 => n52542, B2 => 
                           n59150, ZN => n58627);
   U996 : INV_X1 port map( A => n58627, ZN => n3283);
   U997 : OAI22_X1 port map( A1 => n52463, A2 => n58730, B1 => n52541, B2 => 
                           n59146, ZN => n58628);
   U998 : INV_X1 port map( A => n58628, ZN => n2993);
   U999 : OAI22_X1 port map( A1 => n52443, A2 => n58759, B1 => n52743, B2 => 
                           n59158, ZN => n58629);
   U1000 : INV_X1 port map( A => n58629, ZN => n2846);
   U1001 : OAI22_X1 port map( A1 => n52443, A2 => n58800, B1 => n52742, B2 => 
                           n59158, ZN => n58630);
   U1002 : INV_X1 port map( A => n58630, ZN => n2907);
   U1003 : OAI22_X1 port map( A1 => n52443, A2 => n58913, B1 => n52741, B2 => 
                           n59158, ZN => n58631);
   U1004 : INV_X1 port map( A => n58631, ZN => n2972);
   U1005 : OAI22_X1 port map( A1 => n52457, A2 => n58910, B1 => n52625, B2 => 
                           n59156, ZN => n58632);
   U1006 : INV_X1 port map( A => n58632, ZN => n3382);
   U1007 : OAI22_X1 port map( A1 => n52438, A2 => n58915, B1 => n52546, B2 => 
                           n59183, ZN => n58633);
   U1008 : INV_X1 port map( A => n58633, ZN => n3284);
   U1009 : OAI22_X1 port map( A1 => n52438, A2 => n58913, B1 => n52540, B2 => 
                           n59183, ZN => n58634);
   U1010 : INV_X1 port map( A => n58634, ZN => n2963);
   U1011 : OAI22_X1 port map( A1 => n52438, A2 => n59112, B1 => n52547, B2 => 
                           n59183, ZN => n58635);
   U1012 : INV_X1 port map( A => n58635, ZN => n3027);
   U1013 : OAI22_X1 port map( A1 => n52443, A2 => n58915, B1 => n52740, B2 => 
                           n59158, ZN => n58636);
   U1014 : INV_X1 port map( A => n58636, ZN => n3295);
   U1015 : OAI22_X1 port map( A1 => n52443, A2 => n58789, B1 => n52739, B2 => 
                           n59158, ZN => n58637);
   U1016 : INV_X1 port map( A => n58637, ZN => n3103);
   U1017 : OAI22_X1 port map( A1 => n52438, A2 => n58721, B1 => n52538, B2 => 
                           n59183, ZN => n58638);
   U1018 : INV_X1 port map( A => n58638, ZN => n2866);
   U1019 : OAI22_X1 port map( A1 => n52457, A2 => n59166, B1 => n52622, B2 => 
                           n59156, ZN => n58639);
   U1020 : INV_X1 port map( A => n58639, ZN => n3313);
   U1021 : OAI22_X1 port map( A1 => n52447, A2 => n58915, B1 => n52738, B2 => 
                           n59144, ZN => n58640);
   U1022 : INV_X1 port map( A => n58640, ZN => n3294);
   U1023 : OAI22_X1 port map( A1 => n52439, A2 => n58915, B1 => n52537, B2 => 
                           n59154, ZN => n58641);
   U1024 : INV_X1 port map( A => n58641, ZN => n3282);
   U1025 : OAI22_X1 port map( A1 => n52438, A2 => n58717, B1 => n52549, B2 => 
                           n59183, ZN => n58642);
   U1026 : INV_X1 port map( A => n58642, ZN => n3125);
   U1027 : OAI22_X1 port map( A1 => n52457, A2 => n59112, B1 => n52534, B2 => 
                           n59156, ZN => n58643);
   U1028 : INV_X1 port map( A => n58643, ZN => n3026);
   U1029 : OAI22_X1 port map( A1 => n52439, A2 => n59112, B1 => n52737, B2 => 
                           n59154, ZN => n58644);
   U1030 : INV_X1 port map( A => n58644, ZN => n3036);
   U1031 : OAI22_X1 port map( A1 => n52447, A2 => n58826, B1 => n52763, B2 => 
                           n59144, ZN => n58645);
   U1032 : INV_X1 port map( A => n58645, ZN => n3452);
   U1033 : OAI22_X1 port map( A1 => n52447, A2 => n58759, B1 => n52734, B2 => 
                           n59144, ZN => n58646);
   U1034 : INV_X1 port map( A => n58646, ZN => n2845);
   U1035 : OAI22_X1 port map( A1 => n52463, A2 => n58759, B1 => n52733, B2 => 
                           n59146, ZN => n58647);
   U1036 : INV_X1 port map( A => n58647, ZN => n2844);
   U1037 : OAI22_X1 port map( A1 => n52447, A2 => n58730, B1 => n52620, B2 => 
                           n59144, ZN => n58648);
   U1038 : INV_X1 port map( A => n58648, ZN => n2998);
   U1039 : OAI22_X1 port map( A1 => n52435, A2 => n58741, B1 => n52947, B2 => 
                           n59164, ZN => n58649);
   U1040 : INV_X1 port map( A => n58649, ZN => n2815);
   U1041 : OAI22_X1 port map( A1 => n52463, A2 => n58741, B1 => n52732, B2 => 
                           n59146, ZN => n58650);
   U1042 : INV_X1 port map( A => n58650, ZN => n2812);
   U1043 : OAI22_X1 port map( A1 => n52437, A2 => n58761, B1 => n52550, B2 => 
                           n59150, ZN => n58651);
   U1044 : INV_X1 port map( A => n58651, ZN => n3154);
   U1045 : OAI22_X1 port map( A1 => n52443, A2 => n58910, B1 => n52765, B2 => 
                           n59158, ZN => n58652);
   U1046 : INV_X1 port map( A => n58652, ZN => n3388);
   U1047 : OAI22_X1 port map( A1 => n52453, A2 => n58741, B1 => n52730, B2 => 
                           n59148, ZN => n58653);
   U1048 : INV_X1 port map( A => n58653, ZN => n2811);
   U1049 : OAI22_X1 port map( A1 => n52447, A2 => n58721, B1 => n52613, B2 => 
                           n59144, ZN => n58654);
   U1050 : INV_X1 port map( A => n58654, ZN => n2873);
   U1051 : OAI22_X1 port map( A1 => n52447, A2 => n58655, B1 => n52729, B2 => 
                           n59144, ZN => n58656);
   U1052 : INV_X1 port map( A => n58656, ZN => n2810);
   U1053 : OAI22_X1 port map( A1 => n52453, A2 => n58721, B1 => n52610, B2 => 
                           n59148, ZN => n58657);
   U1054 : INV_X1 port map( A => n58657, ZN => n2870);
   U1055 : OAI22_X1 port map( A1 => n52453, A2 => n58800, B1 => n52766, B2 => 
                           n59148, ZN => n58658);
   U1056 : INV_X1 port map( A => n58658, ZN => n2908);
   U1057 : OAI22_X1 port map( A1 => n52447, A2 => n58800, B1 => n52727, B2 => 
                           n59144, ZN => n58659);
   U1058 : INV_X1 port map( A => n58659, ZN => n2906);
   U1059 : OAI22_X1 port map( A1 => n52443, A2 => n58721, B1 => n52605, B2 => 
                           n59158, ZN => n58660);
   U1060 : INV_X1 port map( A => n58660, ZN => n2869);
   U1061 : OAI22_X1 port map( A1 => n52437, A2 => n58913, B1 => n52551, B2 => 
                           n59150, ZN => n58661);
   U1062 : INV_X1 port map( A => n58661, ZN => n2964);
   U1063 : OAI22_X1 port map( A1 => n52437, A2 => n58826, B1 => n52533, B2 => 
                           n59150, ZN => n58662);
   U1064 : INV_X1 port map( A => n58662, ZN => n3444);
   U1065 : OAI22_X1 port map( A1 => n52453, A2 => n58915, B1 => n52595, B2 => 
                           n59148, ZN => n58663);
   U1066 : INV_X1 port map( A => n58663, ZN => n3288);
   U1067 : OAI22_X1 port map( A1 => n52447, A2 => n58789, B1 => n52726, B2 => 
                           n59144, ZN => n58664);
   U1068 : INV_X1 port map( A => n58664, ZN => n3102);
   U1069 : OAI22_X1 port map( A1 => n52453, A2 => n58761, B1 => n52590, B2 => 
                           n59148, ZN => n58665);
   U1070 : INV_X1 port map( A => n58665, ZN => n3157);
   U1071 : OAI22_X1 port map( A1 => n52453, A2 => n58717, B1 => n52589, B2 => 
                           n59148, ZN => n58666);
   U1072 : INV_X1 port map( A => n58666, ZN => n3129);
   U1073 : OAI22_X1 port map( A1 => n52453, A2 => n58789, B1 => n52588, B2 => 
                           n59148, ZN => n58667);
   U1074 : INV_X1 port map( A => n58667, ZN => n3095);
   U1075 : OAI22_X1 port map( A1 => n52463, A2 => n58800, B1 => n52718, B2 => 
                           n59146, ZN => n58668);
   U1076 : INV_X1 port map( A => n58668, ZN => n2904);
   U1077 : OAI22_X1 port map( A1 => n52437, A2 => n59166, B1 => n52686, B2 => 
                           n59150, ZN => n58669);
   U1078 : INV_X1 port map( A => n58669, ZN => n3320);
   U1079 : OAI22_X1 port map( A1 => n52453, A2 => n58826, B1 => n52665, B2 => 
                           n59148, ZN => n58670);
   U1080 : INV_X1 port map( A => n58670, ZN => n3450);
   U1081 : OAI22_X1 port map( A1 => n52443, A2 => n58813, B1 => n52774, B2 => 
                           n59158, ZN => n58671);
   U1082 : INV_X1 port map( A => n58671, ZN => n3518);
   U1083 : OAI22_X1 port map( A1 => n52457, A2 => n58761, B1 => n52682, B2 => 
                           n59156, ZN => n58672);
   U1084 : INV_X1 port map( A => n58672, ZN => n3161);
   U1085 : OAI22_X1 port map( A1 => n52443, A2 => n59166, B1 => n52779, B2 => 
                           n59158, ZN => n58673);
   U1086 : INV_X1 port map( A => n58673, ZN => n3325);
   U1087 : OAI22_X1 port map( A1 => n52439, A2 => n58721, B1 => n52585, B2 => 
                           n59154, ZN => n58674);
   U1088 : INV_X1 port map( A => n58674, ZN => n2868);
   U1089 : OAI22_X1 port map( A1 => n52439, A2 => n58783, B1 => n52584, B2 => 
                           n59154, ZN => n58675);
   U1090 : INV_X1 port map( A => n58675, ZN => n3252);
   U1091 : OAI22_X1 port map( A1 => n52440, A2 => n58915, B1 => n52566, B2 => 
                           n59152, ZN => n58676);
   U1092 : INV_X1 port map( A => n58676, ZN => n3286);
   U1093 : OAI22_X1 port map( A1 => n52438, A2 => n58761, B1 => n52555, B2 => 
                           n59183, ZN => n58677);
   U1094 : INV_X1 port map( A => n58677, ZN => n3155);
   U1095 : OAI22_X1 port map( A1 => n52437, A2 => n58759, B1 => n52699, B2 => 
                           n59150, ZN => n58678);
   U1096 : INV_X1 port map( A => n58678, ZN => n2841);
   U1097 : OAI22_X1 port map( A1 => n52440, A2 => n58759, B1 => n52698, B2 => 
                           n59152, ZN => n58679);
   U1098 : INV_X1 port map( A => n58679, ZN => n2840);
   U1099 : OAI22_X1 port map( A1 => n52457, A2 => n58793, B1 => n52531, B2 => 
                           n59156, ZN => n58680);
   U1100 : INV_X1 port map( A => n58680, ZN => n2932);
   U1101 : OAI22_X1 port map( A1 => n52439, A2 => n58913, B1 => n52583, B2 => 
                           n59154, ZN => n58681);
   U1102 : INV_X1 port map( A => n58681, ZN => n2966);
   U1103 : OAI22_X1 port map( A1 => n52440, A2 => n58910, B1 => n52530, B2 => 
                           n59152, ZN => n58682);
   U1104 : INV_X1 port map( A => n58682, ZN => n3381);
   U1105 : OAI22_X1 port map( A1 => n52438, A2 => n58759, B1 => n52696, B2 => 
                           n59183, ZN => n58683);
   U1106 : INV_X1 port map( A => n58683, ZN => n2839);
   U1107 : OAI22_X1 port map( A1 => n52439, A2 => n59213, B1 => n52582, B2 => 
                           n59154, ZN => n58684);
   U1108 : INV_X1 port map( A => n58684, ZN => n3192);
   U1109 : OAI22_X1 port map( A1 => n52439, A2 => n58717, B1 => n52581, B2 => 
                           n59154, ZN => n58685);
   U1110 : INV_X1 port map( A => n58685, ZN => n3128);
   U1111 : OAI22_X1 port map( A1 => n52440, A2 => n59166, B1 => n52684, B2 => 
                           n59152, ZN => n58686);
   U1112 : INV_X1 port map( A => n58686, ZN => n3319);
   U1113 : OAI22_X1 port map( A1 => n52447, A2 => n58910, B1 => n52781, B2 => 
                           n59144, ZN => n58687);
   U1114 : INV_X1 port map( A => n58687, ZN => n3390);
   U1115 : OAI22_X1 port map( A1 => n52437, A2 => n58741, B1 => n52709, B2 => 
                           n59150, ZN => n58688);
   U1116 : INV_X1 port map( A => n58688, ZN => n2807);
   U1117 : OAI22_X1 port map( A1 => n52440, A2 => n59213, B1 => n52568, B2 => 
                           n59152, ZN => n58689);
   U1118 : INV_X1 port map( A => n58689, ZN => n3191);
   U1119 : OAI22_X1 port map( A1 => n52457, A2 => n59209, B1 => n52703, B2 => 
                           n59156, ZN => n58690);
   U1120 : INV_X1 port map( A => n58690, ZN => n3544);
   U1121 : OAI22_X1 port map( A1 => n52463, A2 => n58781, B1 => n52565, B2 => 
                           n59146, ZN => n58691);
   U1122 : INV_X1 port map( A => n58691, ZN => n3058);
   U1123 : OAI22_X1 port map( A1 => n52439, A2 => n58730, B1 => n52579, B2 => 
                           n59154, ZN => n58692);
   U1124 : INV_X1 port map( A => n58692, ZN => n2997);
   U1125 : OAI22_X1 port map( A1 => n52463, A2 => n58915, B1 => n52564, B2 => 
                           n59146, ZN => n58693);
   U1126 : INV_X1 port map( A => n58693, ZN => n3285);
   U1127 : OAI22_X1 port map( A1 => n52439, A2 => n58781, B1 => n52578, B2 => 
                           n59154, ZN => n58694);
   U1128 : INV_X1 port map( A => n58694, ZN => n3060);
   U1129 : OAI22_X1 port map( A1 => n52463, A2 => n59173, B1 => n52708, B2 => 
                           n59146, ZN => n58695);
   U1130 : INV_X1 port map( A => n58695, ZN => n3220);
   U1131 : OAI22_X1 port map( A1 => n52440, A2 => n58793, B1 => n52577, B2 => 
                           n59152, ZN => n58696);
   U1132 : INV_X1 port map( A => n58696, ZN => n2935);
   U1133 : OAI22_X1 port map( A1 => n52440, A2 => n58913, B1 => n52576, B2 => 
                           n59152, ZN => n58697);
   U1134 : INV_X1 port map( A => n58697, ZN => n2965);
   U1135 : OAI22_X1 port map( A1 => n52443, A2 => n59112, B1 => n52685, B2 => 
                           n59158, ZN => n58698);
   U1136 : INV_X1 port map( A => n58698, ZN => n3032);
   U1137 : OAI22_X1 port map( A1 => n52437, A2 => n59213, B1 => n52558, B2 => 
                           n59150, ZN => n58699);
   U1138 : INV_X1 port map( A => n58699, ZN => n3190);
   U1139 : OAI22_X1 port map( A1 => n52439, A2 => n58800, B1 => n52706, B2 => 
                           n59154, ZN => n58700);
   U1140 : INV_X1 port map( A => n58700, ZN => n2903);
   U1141 : OAI22_X1 port map( A1 => n52443, A2 => n58761, B1 => n52778, B2 => 
                           n59158, ZN => n58701);
   U1142 : INV_X1 port map( A => n58701, ZN => n3163);
   U1143 : OAI22_X1 port map( A1 => n52440, A2 => n58730, B1 => n52575, B2 => 
                           n59152, ZN => n58702);
   U1144 : INV_X1 port map( A => n58702, ZN => n2996);
   U1145 : OAI22_X1 port map( A1 => n52443, A2 => n58717, B1 => n52782, B2 => 
                           n59158, ZN => n58703);
   U1146 : INV_X1 port map( A => n58703, ZN => n3133);
   U1147 : OAI22_X1 port map( A1 => n52439, A2 => n58759, B1 => n52689, B2 => 
                           n59154, ZN => n58704);
   U1148 : INV_X1 port map( A => n58704, ZN => n2835);
   U1149 : OAI22_X1 port map( A1 => n52437, A2 => n58781, B1 => n52552, B2 => 
                           n59150, ZN => n58705);
   U1150 : INV_X1 port map( A => n58705, ZN => n3057);
   U1151 : OAI22_X1 port map( A1 => n52440, A2 => n59112, B1 => n52574, B2 => 
                           n59152, ZN => n58706);
   U1152 : INV_X1 port map( A => n58706, ZN => n3029);
   U1153 : OAI22_X1 port map( A1 => n52463, A2 => n59169, B1 => n52561, B2 => 
                           n59146, ZN => n58707);
   U1154 : INV_X1 port map( A => n58707, ZN => n3477);
   U1155 : OAI22_X1 port map( A1 => n52439, A2 => n58741, B1 => n52688, B2 => 
                           n59154, ZN => n58708);
   U1156 : INV_X1 port map( A => n58708, ZN => n2803);
   U1157 : OAI22_X1 port map( A1 => n52457, A2 => n58759, B1 => n52693, B2 => 
                           n59156, ZN => n58709);
   U1158 : INV_X1 port map( A => n58709, ZN => n2837);
   U1159 : OAI22_X1 port map( A1 => n52440, A2 => n58761, B1 => n52569, B2 => 
                           n59152, ZN => n58710);
   U1160 : INV_X1 port map( A => n58710, ZN => n3156);
   U1161 : OAI22_X1 port map( A1 => n52457, A2 => n58741, B1 => n52692, B2 => 
                           n59156, ZN => n58711);
   U1162 : INV_X1 port map( A => n58711, ZN => n2805);
   U1163 : OAI22_X1 port map( A1 => n52437, A2 => n58730, B1 => n52572, B2 => 
                           n59150, ZN => n58712);
   U1164 : INV_X1 port map( A => n58712, ZN => n2995);
   U1165 : OAI22_X1 port map( A1 => n52463, A2 => n58819, B1 => n52529, B2 => 
                           n59146, ZN => n58713);
   U1166 : INV_X1 port map( A => n58713, ZN => n3348);
   U1167 : OAI22_X1 port map( A1 => n52439, A2 => n59166, B1 => n52687, B2 => 
                           n59154, ZN => n58714);
   U1168 : INV_X1 port map( A => n58714, ZN => n3321);
   U1169 : OAI22_X1 port map( A1 => n52440, A2 => n58717, B1 => n52570, B2 => 
                           n59152, ZN => n58715);
   U1170 : INV_X1 port map( A => n58715, ZN => n3127);
   U1171 : OAI22_X1 port map( A1 => n52463, A2 => n59112, B1 => n52562, B2 => 
                           n59146, ZN => n58716);
   U1172 : INV_X1 port map( A => n58716, ZN => n3028);
   U1173 : OAI22_X1 port map( A1 => n52437, A2 => n58717, B1 => n52560, B2 => 
                           n59150, ZN => n58718);
   U1174 : INV_X1 port map( A => n58718, ZN => n3126);
   U1175 : OAI22_X1 port map( A1 => n52435, A2 => n58721, B1 => n52854, B2 => 
                           n59164, ZN => n58719);
   U1176 : INV_X1 port map( A => n58719, ZN => n2875);
   U1177 : OAI22_X1 port map( A1 => n52437, A2 => n58789, B1 => n52559, B2 => 
                           n59150, ZN => n58720);
   U1178 : INV_X1 port map( A => n58720, ZN => n3092);
   U1179 : OAI22_X1 port map( A1 => n52437, A2 => n58721, B1 => n52557, B2 => 
                           n59150, ZN => n58722);
   U1180 : INV_X1 port map( A => n58722, ZN => n2867);
   U1181 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n52452, ZN => n59134);
   U1182 : OAI22_X1 port map( A1 => n52452, A2 => n58789, B1 => n53084, B2 => 
                           n59134, ZN => n58723);
   U1183 : INV_X1 port map( A => n58723, ZN => n3109);
   U1184 : OAI22_X1 port map( A1 => n52452, A2 => n58813, B1 => n53036, B2 => 
                           n59134, ZN => n58724);
   U1185 : INV_X1 port map( A => n58724, ZN => n3503);
   U1186 : OAI22_X1 port map( A1 => n52452, A2 => n58725, B1 => n53072, B2 => 
                           n59134, ZN => n58726);
   U1187 : INV_X1 port map( A => n58726, ZN => n2856);
   U1188 : OAI22_X1 port map( A1 => n52452, A2 => n58800, B1 => n53070, B2 => 
                           n59134, ZN => n58727);
   U1189 : INV_X1 port map( A => n58727, ZN => n2917);
   U1190 : OAI22_X1 port map( A1 => n52452, A2 => n58811, B1 => n53039, B2 => 
                           n59134, ZN => n58728);
   U1191 : INV_X1 port map( A => n58728, ZN => n3407);
   U1192 : OAI22_X1 port map( A1 => n52452, A2 => n58793, B1 => n53087, B2 => 
                           n59134, ZN => n58729);
   U1193 : INV_X1 port map( A => n58729, ZN => n2927);
   U1194 : OAI22_X1 port map( A1 => n52452, A2 => n58730, B1 => n53063, B2 => 
                           n59134, ZN => n58731);
   U1195 : INV_X1 port map( A => n58731, ZN => n3013);
   U1196 : OAI22_X1 port map( A1 => n52452, A2 => n58915, B1 => n53080, B2 => 
                           n59134, ZN => n58732);
   U1197 : INV_X1 port map( A => n58732, ZN => n3301);
   U1198 : OAI22_X1 port map( A1 => n52452, A2 => n58826, B1 => n53034, B2 => 
                           n59134, ZN => n58733);
   U1199 : INV_X1 port map( A => n58733, ZN => n3439);
   U1200 : OAI22_X1 port map( A1 => n52452, A2 => n59169, B1 => n53035, B2 => 
                           n59134, ZN => n58734);
   U1201 : INV_X1 port map( A => n58734, ZN => n3471);
   U1202 : OAI22_X1 port map( A1 => n52452, A2 => n58819, B1 => n53042, B2 => 
                           n59134, ZN => n58735);
   U1203 : INV_X1 port map( A => n58735, ZN => n3343);
   U1204 : OAI22_X1 port map( A1 => n52452, A2 => n58736, B1 => n53081, B2 => 
                           n59134, ZN => n58737);
   U1205 : INV_X1 port map( A => n58737, ZN => n3177);
   U1206 : OAI22_X1 port map( A1 => n52452, A2 => n58759, B1 => n52999, B2 => 
                           n59134, ZN => n58738);
   U1207 : INV_X1 port map( A => n58738, ZN => n2851);
   U1208 : OAI22_X1 port map( A1 => n52452, A2 => n58761, B1 => n53082, B2 => 
                           n59134, ZN => n58739);
   U1209 : INV_X1 port map( A => n58739, ZN => n3169);
   U1210 : OAI22_X1 port map( A1 => n52452, A2 => n58910, B1 => n53038, B2 => 
                           n59134, ZN => n58740);
   U1211 : INV_X1 port map( A => n58740, ZN => n3375);
   U1212 : OAI22_X1 port map( A1 => n52452, A2 => n58741, B1 => n53003, B2 => 
                           n59134, ZN => n58742);
   U1213 : INV_X1 port map( A => n58742, ZN => n2816);
   U1214 : OAI22_X1 port map( A1 => n52452, A2 => n59166, B1 => n53040, B2 => 
                           n59134, ZN => n58743);
   U1215 : INV_X1 port map( A => n58743, ZN => n3311);
   U1216 : OAI22_X1 port map( A1 => n52452, A2 => n58781, B1 => n53085, B2 => 
                           n59134, ZN => n58744);
   U1217 : INV_X1 port map( A => n58744, ZN => n3077);
   U1218 : OAI22_X1 port map( A1 => n52452, A2 => n58745, B1 => n53083, B2 => 
                           n59134, ZN => n58746);
   U1219 : INV_X1 port map( A => n58746, ZN => n3113);
   U1220 : OAI22_X1 port map( A1 => n52452, A2 => n58913, B1 => n53086, B2 => 
                           n59134, ZN => n58747);
   U1221 : INV_X1 port map( A => n58747, ZN => n2980);
   U1222 : CLKBUF_X1 port map( A => n59209, Z => n58757);
   U1223 : OAI22_X1 port map( A1 => n52441, A2 => n58757, B1 => n53184, B2 => 
                           n59161, ZN => n58748);
   U1224 : INV_X1 port map( A => n58748, ZN => n3531);
   U1225 : OAI22_X1 port map( A1 => n52448, A2 => n58757, B1 => n53182, B2 => 
                           n59171, ZN => n58749);
   U1226 : INV_X1 port map( A => n58749, ZN => n3529);
   U1227 : OAI22_X1 port map( A1 => n52435, A2 => n58757, B1 => n53185, B2 => 
                           n59164, ZN => n58750);
   U1228 : INV_X1 port map( A => n58750, ZN => n3532);
   U1229 : OAI22_X1 port map( A1 => n52450, A2 => n58757, B1 => n53186, B2 => 
                           n59175, ZN => n58751);
   U1230 : INV_X1 port map( A => n58751, ZN => n3533);
   U1231 : OAI22_X1 port map( A1 => n52463, A2 => n58757, B1 => n52536, B2 => 
                           n59146, ZN => n58752);
   U1232 : INV_X1 port map( A => n58752, ZN => n3539);
   U1233 : OAI22_X1 port map( A1 => n52477, A2 => n58757, B1 => n52893, B2 => 
                           n59126, ZN => n58753);
   U1234 : INV_X1 port map( A => n58753, ZN => n3527);
   U1235 : OAI22_X1 port map( A1 => n52468, A2 => n58757, B1 => n52891, B2 => 
                           n59082, ZN => n58754);
   U1236 : INV_X1 port map( A => n58754, ZN => n3526);
   U1237 : OAI22_X1 port map( A1 => n52447, A2 => n58757, B1 => n53521, B2 => 
                           n59144, ZN => n58755);
   U1238 : INV_X1 port map( A => n58755, ZN => n3541);
   U1239 : OAI22_X1 port map( A1 => n52473, A2 => n58757, B1 => n52897, B2 => 
                           n59130, ZN => n58756);
   U1240 : INV_X1 port map( A => n58756, ZN => n3528);
   U1241 : OAI22_X1 port map( A1 => n52452, A2 => n58757, B1 => n53183, B2 => 
                           n59134, ZN => n58758);
   U1242 : INV_X1 port map( A => n58758, ZN => n3530);
   U1243 : CLKBUF_X1 port map( A => n58759, Z => n58776);
   U1244 : OAI22_X1 port map( A1 => n52455, A2 => n58776, B1 => n52715, B2 => 
                           n58985, ZN => n58760);
   U1245 : INV_X1 port map( A => n58760, ZN => n2842);
   U1246 : CLKBUF_X1 port map( A => n58761, Z => n58779);
   U1247 : OAI22_X1 port map( A1 => n52445, A2 => n58779, B1 => n53113, B2 => 
                           n58967, ZN => n58762);
   U1248 : INV_X1 port map( A => n58762, ZN => n3145);
   U1249 : OAI22_X1 port map( A1 => n52450, A2 => n58776, B1 => n53176, B2 => 
                           n59175, ZN => n58763);
   U1250 : INV_X1 port map( A => n58763, ZN => n2829);
   U1251 : OAI22_X1 port map( A1 => n52442, A2 => n58776, B1 => n53148, B2 => 
                           n59168, ZN => n58764);
   U1252 : INV_X1 port map( A => n58764, ZN => n2826);
   U1253 : OAI22_X1 port map( A1 => n52445, A2 => n58776, B1 => n53166, B2 => 
                           n58967, ZN => n58765);
   U1254 : INV_X1 port map( A => n58765, ZN => n2828);
   U1255 : OAI22_X1 port map( A1 => n52467, A2 => n58779, B1 => n53165, B2 => 
                           n59212, ZN => n58766);
   U1256 : INV_X1 port map( A => n58766, ZN => n3147);
   U1257 : OAI22_X1 port map( A1 => n52444, A2 => n58776, B1 => n53110, B2 => 
                           n59128, ZN => n58767);
   U1258 : INV_X1 port map( A => n58767, ZN => n2825);
   U1259 : OAI22_X1 port map( A1 => n52439, A2 => n58779, B1 => n53201, B2 => 
                           n59154, ZN => n58768);
   U1260 : INV_X1 port map( A => n58768, ZN => n3148);
   U1261 : OAI22_X1 port map( A1 => n52478, A2 => n58779, B1 => n52813, B2 => 
                           n58980, ZN => n58769);
   U1262 : INV_X1 port map( A => n58769, ZN => n3143);
   U1263 : OAI22_X1 port map( A1 => n52441, A2 => n58776, B1 => n53163, B2 => 
                           n59161, ZN => n58770);
   U1264 : INV_X1 port map( A => n58770, ZN => n2827);
   U1265 : OAI22_X1 port map( A1 => n52459, A2 => n58776, B1 => n52860, B2 => 
                           n58993, ZN => n58771);
   U1266 : INV_X1 port map( A => n58771, ZN => n2822);
   U1267 : OAI22_X1 port map( A1 => n52448, A2 => n58779, B1 => n53041, B2 => 
                           n59171, ZN => n58772);
   U1268 : INV_X1 port map( A => n58772, ZN => n3144);
   U1269 : OAI22_X1 port map( A1 => n52469, A2 => n58776, B1 => n52863, B2 => 
                           n58996, ZN => n58773);
   U1270 : INV_X1 port map( A => n58773, ZN => n2823);
   U1271 : OAI22_X1 port map( A1 => n52455, A2 => n58779, B1 => n52711, B2 => 
                           n58985, ZN => n58774);
   U1272 : INV_X1 port map( A => n58774, ZN => n3162);
   U1273 : OAI22_X1 port map( A1 => n52450, A2 => n58779, B1 => n53129, B2 => 
                           n59175, ZN => n58775);
   U1274 : INV_X1 port map( A => n58775, ZN => n3146);
   U1275 : OAI22_X1 port map( A1 => n52478, A2 => n58776, B1 => n52912, B2 => 
                           n58980, ZN => n58777);
   U1276 : INV_X1 port map( A => n58777, ZN => n2824);
   U1277 : OAI22_X1 port map( A1 => n52463, A2 => n58779, B1 => n53238, B2 => 
                           n59146, ZN => n58778);
   U1278 : INV_X1 port map( A => n58778, ZN => n3149);
   U1279 : OAI22_X1 port map( A1 => n52473, A2 => n58779, B1 => n52812, B2 => 
                           n59130, ZN => n58780);
   U1280 : INV_X1 port map( A => n58780, ZN => n3142);
   U1281 : CLKBUF_X1 port map( A => n58781, Z => n58897);
   U1282 : OAI22_X1 port map( A1 => n52442, A2 => n58897, B1 => n53136, B2 => 
                           n59168, ZN => n58782);
   U1283 : INV_X1 port map( A => n58782, ZN => n3053);
   U1284 : CLKBUF_X1 port map( A => n58783, Z => n58904);
   U1285 : OAI22_X1 port map( A1 => n52467, A2 => n58904, B1 => n53139, B2 => 
                           n59212, ZN => n58784);
   U1286 : INV_X1 port map( A => n58784, ZN => n3241);
   U1287 : OAI22_X1 port map( A1 => n52442, A2 => n58904, B1 => n53140, B2 => 
                           n59168, ZN => n58785);
   U1288 : INV_X1 port map( A => n58785, ZN => n3242);
   U1289 : OAI22_X1 port map( A1 => n52450, A2 => n58897, B1 => n53134, B2 => 
                           n59175, ZN => n58786);
   U1290 : INV_X1 port map( A => n58786, ZN => n3052);
   U1291 : OAI22_X1 port map( A1 => n52441, A2 => n58897, B1 => n53133, B2 => 
                           n59161, ZN => n58787);
   U1292 : INV_X1 port map( A => n58787, ZN => n3051);
   U1293 : OAI22_X1 port map( A1 => n52445, A2 => n58897, B1 => n53132, B2 => 
                           n58967, ZN => n58788);
   U1294 : INV_X1 port map( A => n58788, ZN => n3050);
   U1295 : CLKBUF_X1 port map( A => n58789, Z => n58908);
   U1296 : OAI22_X1 port map( A1 => n52450, A2 => n58908, B1 => n53131, B2 => 
                           n59175, ZN => n58790);
   U1297 : INV_X1 port map( A => n58790, ZN => n3083);
   U1298 : OAI22_X1 port map( A1 => n52448, A2 => n58904, B1 => n53141, B2 => 
                           n59171, ZN => n58791);
   U1299 : INV_X1 port map( A => n58791, ZN => n3243);
   U1300 : OAI22_X1 port map( A1 => n52456, A2 => n58904, B1 => n53278, B2 => 
                           n58982, ZN => n58792);
   U1301 : INV_X1 port map( A => n58792, ZN => n3244);
   U1302 : CLKBUF_X1 port map( A => n58793, Z => n58902);
   U1303 : OAI22_X1 port map( A1 => n52446, A2 => n58902, B1 => n53310, B2 => 
                           n58978, ZN => n58794);
   U1304 : INV_X1 port map( A => n58794, ZN => n2924);
   U1305 : OAI22_X1 port map( A1 => n52447, A2 => n58902, B1 => n53317, B2 => 
                           n59144, ZN => n58795);
   U1306 : INV_X1 port map( A => n58795, ZN => n2923);
   U1307 : OAI22_X1 port map( A1 => n52463, A2 => n58904, B1 => n53318, B2 => 
                           n59146, ZN => n58796);
   U1308 : INV_X1 port map( A => n58796, ZN => n3245);
   U1309 : OAI22_X1 port map( A1 => n52455, A2 => n58902, B1 => n53259, B2 => 
                           n58985, ZN => n58797);
   U1310 : INV_X1 port map( A => n58797, ZN => n2925);
   U1311 : OAI22_X1 port map( A1 => n52443, A2 => n58902, B1 => n53333, B2 => 
                           n59158, ZN => n58798);
   U1312 : INV_X1 port map( A => n58798, ZN => n2922);
   U1313 : OAI22_X1 port map( A1 => n52467, A2 => n58908, B1 => n53150, B2 => 
                           n59212, ZN => n58799);
   U1314 : INV_X1 port map( A => n58799, ZN => n3084);
   U1315 : CLKBUF_X1 port map( A => n58800, Z => n58885);
   U1316 : OAI22_X1 port map( A1 => n52450, A2 => n58885, B1 => n53154, B2 => 
                           n59175, ZN => n58801);
   U1317 : INV_X1 port map( A => n58801, ZN => n2890);
   U1318 : OAI22_X1 port map( A1 => n52445, A2 => n58885, B1 => n53155, B2 => 
                           n58967, ZN => n58802);
   U1319 : INV_X1 port map( A => n58802, ZN => n2891);
   U1320 : OAI22_X1 port map( A1 => n52442, A2 => n58885, B1 => n53156, B2 => 
                           n59168, ZN => n58803);
   U1321 : INV_X1 port map( A => n58803, ZN => n2892);
   U1322 : OAI22_X1 port map( A1 => n52442, A2 => n58908, B1 => n53160, B2 => 
                           n59168, ZN => n58804);
   U1323 : INV_X1 port map( A => n58804, ZN => n3085);
   U1324 : OAI22_X1 port map( A1 => n52453, A2 => n58902, B1 => n53354, B2 => 
                           n59148, ZN => n58805);
   U1325 : INV_X1 port map( A => n58805, ZN => n2921);
   U1326 : OAI22_X1 port map( A1 => n52441, A2 => n58885, B1 => n53164, B2 => 
                           n59161, ZN => n58806);
   U1327 : INV_X1 port map( A => n58806, ZN => n2893);
   U1328 : OAI22_X1 port map( A1 => n52473, A2 => n58902, B1 => n53356, B2 => 
                           n59130, ZN => n58807);
   U1329 : INV_X1 port map( A => n58807, ZN => n2920);
   U1330 : OAI22_X1 port map( A1 => n52469, A2 => n58902, B1 => n53358, B2 => 
                           n58996, ZN => n58808);
   U1331 : INV_X1 port map( A => n58808, ZN => n2919);
   U1332 : OAI22_X1 port map( A1 => n52468, A2 => n58902, B1 => n53362, B2 => 
                           n59082, ZN => n58809);
   U1333 : INV_X1 port map( A => n58809, ZN => n2918);
   U1334 : OAI22_X1 port map( A1 => n52445, A2 => n58908, B1 => n53123, B2 => 
                           n58967, ZN => n58810);
   U1335 : INV_X1 port map( A => n58810, ZN => n3082);
   U1336 : CLKBUF_X1 port map( A => n58811, Z => n58894);
   U1337 : OAI22_X1 port map( A1 => n52459, A2 => n58894, B1 => n52911, B2 => 
                           n58993, ZN => n58812);
   U1338 : INV_X1 port map( A => n58812, ZN => n3400);
   U1339 : CLKBUF_X1 port map( A => n58813, Z => n58891);
   U1340 : OAI22_X1 port map( A1 => n52459, A2 => n58891, B1 => n52909, B2 => 
                           n58993, ZN => n58814);
   U1341 : INV_X1 port map( A => n58814, ZN => n3496);
   U1342 : OAI22_X1 port map( A1 => n52473, A2 => n58908, B1 => n52825, B2 => 
                           n59130, ZN => n58815);
   U1343 : INV_X1 port map( A => n58815, ZN => n3080);
   U1344 : OAI22_X1 port map( A1 => n52468, A2 => n58908, B1 => n52822, B2 => 
                           n59082, ZN => n58816);
   U1345 : INV_X1 port map( A => n58816, ZN => n3079);
   U1346 : OAI22_X1 port map( A1 => n52469, A2 => n58908, B1 => n52821, B2 => 
                           n58996, ZN => n58817);
   U1347 : INV_X1 port map( A => n58817, ZN => n3078);
   U1348 : OAI22_X1 port map( A1 => n52438, A2 => n58908, B1 => n52548, B2 => 
                           n59183, ZN => n58818);
   U1349 : INV_X1 port map( A => n58818, ZN => n3091);
   U1350 : CLKBUF_X1 port map( A => n58819, Z => n58887);
   U1351 : OAI22_X1 port map( A1 => n52435, A2 => n58887, B1 => n52888, B2 => 
                           n59164, ZN => n58820);
   U1352 : INV_X1 port map( A => n58820, ZN => n3335);
   U1353 : OAI22_X1 port map( A1 => n52436, A2 => n58891, B1 => n52886, B2 => 
                           n59124, ZN => n58821);
   U1354 : INV_X1 port map( A => n58821, ZN => n3495);
   U1355 : OAI22_X1 port map( A1 => n52437, A2 => n58902, B1 => n52553, B2 => 
                           n59150, ZN => n58822);
   U1356 : INV_X1 port map( A => n58822, ZN => n2934);
   U1357 : OAI22_X1 port map( A1 => n52435, A2 => n58894, B1 => n52884, B2 => 
                           n59164, ZN => n58823);
   U1358 : INV_X1 port map( A => n58823, ZN => n3399);
   U1359 : OAI22_X1 port map( A1 => n52463, A2 => n58891, B1 => n52554, B2 => 
                           n59146, ZN => n58824);
   U1360 : INV_X1 port map( A => n58824, ZN => n3509);
   U1361 : OAI22_X1 port map( A1 => n52435, A2 => n58891, B1 => n52881, B2 => 
                           n59164, ZN => n58825);
   U1362 : INV_X1 port map( A => n58825, ZN => n3494);
   U1363 : CLKBUF_X1 port map( A => n58826, Z => n58900);
   U1364 : OAI22_X1 port map( A1 => n52436, A2 => n58900, B1 => n52879, B2 => 
                           n59124, ZN => n58827);
   U1365 : INV_X1 port map( A => n58827, ZN => n3430);
   U1366 : OAI22_X1 port map( A1 => n52463, A2 => n58900, B1 => n52556, B2 => 
                           n59146, ZN => n58828);
   U1367 : INV_X1 port map( A => n58828, ZN => n3445);
   U1368 : OAI22_X1 port map( A1 => n52436, A2 => n58894, B1 => n52878, B2 => 
                           n59124, ZN => n58829);
   U1369 : INV_X1 port map( A => n58829, ZN => n3398);
   U1370 : OAI22_X1 port map( A1 => n52463, A2 => n58894, B1 => n52563, B2 => 
                           n59146, ZN => n58830);
   U1371 : INV_X1 port map( A => n58830, ZN => n3413);
   U1372 : OAI22_X1 port map( A1 => n52440, A2 => n58904, B1 => n52567, B2 => 
                           n59152, ZN => n58831);
   U1373 : INV_X1 port map( A => n58831, ZN => n3251);
   U1374 : OAI22_X1 port map( A1 => n52440, A2 => n58908, B1 => n52571, B2 => 
                           n59152, ZN => n58832);
   U1375 : INV_X1 port map( A => n58832, ZN => n3093);
   U1376 : OAI22_X1 port map( A1 => n52440, A2 => n58897, B1 => n52573, B2 => 
                           n59152, ZN => n58833);
   U1377 : INV_X1 port map( A => n58833, ZN => n3059);
   U1378 : CLKBUF_X1 port map( A => n59166, Z => n58906);
   U1379 : OAI22_X1 port map( A1 => n52459, A2 => n58906, B1 => n52876, B2 => 
                           n58993, ZN => n58834);
   U1380 : INV_X1 port map( A => n58834, ZN => n3304);
   U1381 : OAI22_X1 port map( A1 => n52436, A2 => n58887, B1 => n52875, B2 => 
                           n59124, ZN => n58835);
   U1382 : INV_X1 port map( A => n58835, ZN => n3334);
   U1383 : OAI22_X1 port map( A1 => n52459, A2 => n58885, B1 => n52870, B2 => 
                           n58993, ZN => n58836);
   U1384 : INV_X1 port map( A => n58836, ZN => n2887);
   U1385 : OAI22_X1 port map( A1 => n52477, A2 => n58885, B1 => n52869, B2 => 
                           n59126, ZN => n58837);
   U1386 : INV_X1 port map( A => n58837, ZN => n2886);
   U1387 : OAI22_X1 port map( A1 => n52473, A2 => n58906, B1 => n52867, B2 => 
                           n59130, ZN => n58838);
   U1388 : INV_X1 port map( A => n58838, ZN => n3303);
   U1389 : OAI22_X1 port map( A1 => n52439, A2 => n58908, B1 => n52580, B2 => 
                           n59154, ZN => n58839);
   U1390 : INV_X1 port map( A => n58839, ZN => n3094);
   U1391 : OAI22_X1 port map( A1 => n52469, A2 => n58906, B1 => n52866, B2 => 
                           n58996, ZN => n58840);
   U1392 : INV_X1 port map( A => n58840, ZN => n3302);
   U1393 : OAI22_X1 port map( A1 => n52453, A2 => n58897, B1 => n52587, B2 => 
                           n59148, ZN => n58841);
   U1394 : INV_X1 port map( A => n58841, ZN => n3061);
   U1395 : OAI22_X1 port map( A1 => n52468, A2 => n58900, B1 => n52927, B2 => 
                           n59082, ZN => n58842);
   U1396 : INV_X1 port map( A => n58842, ZN => n3432);
   U1397 : OAI22_X1 port map( A1 => n52451, A2 => n58904, B1 => n52592, B2 => 
                           n58999, ZN => n58843);
   U1398 : INV_X1 port map( A => n58843, ZN => n3253);
   U1399 : OAI22_X1 port map( A1 => n52453, A2 => n58904, B1 => n52594, B2 => 
                           n59148, ZN => n58844);
   U1400 : INV_X1 port map( A => n58844, ZN => n3254);
   U1401 : OAI22_X1 port map( A1 => n52477, A2 => n58897, B1 => n52932, B2 => 
                           n59126, ZN => n58845);
   U1402 : INV_X1 port map( A => n58845, ZN => n3047);
   U1403 : OAI22_X1 port map( A1 => n52435, A2 => n58897, B1 => n52858, B2 => 
                           n59164, ZN => n58846);
   U1404 : INV_X1 port map( A => n58846, ZN => n3046);
   U1405 : OAI22_X1 port map( A1 => n52477, A2 => n58887, B1 => n52935, B2 => 
                           n59126, ZN => n58847);
   U1406 : INV_X1 port map( A => n58847, ZN => n3336);
   U1407 : OAI22_X1 port map( A1 => n52435, A2 => n58900, B1 => n52883, B2 => 
                           n59164, ZN => n58848);
   U1408 : INV_X1 port map( A => n58848, ZN => n3431);
   U1409 : OAI22_X1 port map( A1 => n52445, A2 => n58891, B1 => n53012, B2 => 
                           n58967, ZN => n58849);
   U1410 : INV_X1 port map( A => n58849, ZN => n3497);
   U1411 : OAI22_X1 port map( A1 => n52449, A2 => n58897, B1 => n52615, B2 => 
                           n58976, ZN => n58850);
   U1412 : INV_X1 port map( A => n58850, ZN => n3062);
   U1413 : OAI22_X1 port map( A1 => n52448, A2 => n58894, B1 => n53022, B2 => 
                           n59171, ZN => n58851);
   U1414 : INV_X1 port map( A => n58851, ZN => n3404);
   U1415 : OAI22_X1 port map( A1 => n52444, A2 => n58900, B1 => n53025, B2 => 
                           n59128, ZN => n58852);
   U1416 : INV_X1 port map( A => n58852, ZN => n3435);
   U1417 : OAI22_X1 port map( A1 => n52442, A2 => n58900, B1 => n53026, B2 => 
                           n59168, ZN => n58853);
   U1418 : INV_X1 port map( A => n58853, ZN => n3436);
   U1419 : OAI22_X1 port map( A1 => n52438, A2 => n58902, B1 => n52539, B2 => 
                           n59183, ZN => n58854);
   U1420 : INV_X1 port map( A => n58854, ZN => n2933);
   U1421 : OAI22_X1 port map( A1 => n52441, A2 => n58900, B1 => n53030, B2 => 
                           n59161, ZN => n58855);
   U1422 : INV_X1 port map( A => n58855, ZN => n3437);
   U1423 : OAI22_X1 port map( A1 => n52438, A2 => n58906, B1 => n52683, B2 => 
                           n59183, ZN => n58856);
   U1424 : INV_X1 port map( A => n58856, ZN => n3318);
   U1425 : OAI22_X1 port map( A1 => n52450, A2 => n58906, B1 => n52996, B2 => 
                           n59175, ZN => n58857);
   U1426 : INV_X1 port map( A => n58857, ZN => n3308);
   U1427 : OAI22_X1 port map( A1 => n52455, A2 => n58885, B1 => n52656, B2 => 
                           n58985, ZN => n58858);
   U1428 : INV_X1 port map( A => n58858, ZN => n2899);
   U1429 : OAI22_X1 port map( A1 => n52439, A2 => n58887, B1 => n52501, B2 => 
                           n59154, ZN => n58859);
   U1430 : INV_X1 port map( A => n58859, ZN => n3347);
   U1431 : OAI22_X1 port map( A1 => n52450, A2 => n58887, B1 => n52993, B2 => 
                           n59175, ZN => n58860);
   U1432 : INV_X1 port map( A => n58860, ZN => n3339);
   U1433 : OAI22_X1 port map( A1 => n52454, A2 => n58887, B1 => n52992, B2 => 
                           n59120, ZN => n58861);
   U1434 : INV_X1 port map( A => n58861, ZN => n3338);
   U1435 : OAI22_X1 port map( A1 => n52458, A2 => n58891, B1 => n52627, B2 => 
                           n59006, ZN => n58862);
   U1436 : INV_X1 port map( A => n58862, ZN => n3510);
   U1437 : OAI22_X1 port map( A1 => n52442, A2 => n58887, B1 => n52997, B2 => 
                           n59168, ZN => n58863);
   U1438 : INV_X1 port map( A => n58863, ZN => n3340);
   U1439 : OAI22_X1 port map( A1 => n52438, A2 => n58887, B1 => n52535, B2 => 
                           n59183, ZN => n58864);
   U1440 : INV_X1 port map( A => n58864, ZN => n3349);
   U1441 : OAI22_X1 port map( A1 => n52444, A2 => n58885, B1 => n53107, B2 => 
                           n59128, ZN => n58865);
   U1442 : INV_X1 port map( A => n58865, ZN => n2889);
   U1443 : OAI22_X1 port map( A1 => n52445, A2 => n58887, B1 => n52998, B2 => 
                           n58967, ZN => n58866);
   U1444 : INV_X1 port map( A => n58866, ZN => n3341);
   U1445 : OAI22_X1 port map( A1 => n52453, A2 => n58906, B1 => n52662, B2 => 
                           n59148, ZN => n58867);
   U1446 : INV_X1 port map( A => n58867, ZN => n3317);
   U1447 : OAI22_X1 port map( A1 => n52445, A2 => n58894, B1 => n53001, B2 => 
                           n58967, ZN => n58868);
   U1448 : INV_X1 port map( A => n58868, ZN => n3401);
   U1449 : OAI22_X1 port map( A1 => n52452, A2 => n58904, B1 => n53079, B2 => 
                           n59134, ZN => n58869);
   U1450 : INV_X1 port map( A => n58869, ZN => n3240);
   U1451 : OAI22_X1 port map( A1 => n52448, A2 => n58906, B1 => n53007, B2 => 
                           n59171, ZN => n58870);
   U1452 : INV_X1 port map( A => n58870, ZN => n3309);
   U1453 : OAI22_X1 port map( A1 => n52445, A2 => n58900, B1 => n53008, B2 => 
                           n58967, ZN => n58871);
   U1454 : INV_X1 port map( A => n58871, ZN => n3433);
   U1455 : OAI22_X1 port map( A1 => n52444, A2 => n58906, B1 => n52989, B2 => 
                           n59128, ZN => n58872);
   U1456 : INV_X1 port map( A => n58872, ZN => n3307);
   U1457 : OAI22_X1 port map( A1 => n52442, A2 => n58891, B1 => n53028, B2 => 
                           n59168, ZN => n58873);
   U1458 : INV_X1 port map( A => n58873, ZN => n3500);
   U1459 : OAI22_X1 port map( A1 => n52440, A2 => n58885, B1 => n52702, B2 => 
                           n59152, ZN => n58874);
   U1460 : INV_X1 port map( A => n58874, ZN => n2902);
   U1461 : OAI22_X1 port map( A1 => n52457, A2 => n58894, B1 => n52621, B2 => 
                           n59156, ZN => n58875);
   U1462 : INV_X1 port map( A => n58875, ZN => n3414);
   U1463 : OAI22_X1 port map( A1 => n52454, A2 => n58894, B1 => n53014, B2 => 
                           n59120, ZN => n58876);
   U1464 : INV_X1 port map( A => n58876, ZN => n3402);
   U1465 : OAI22_X1 port map( A1 => n52454, A2 => n58900, B1 => n53015, B2 => 
                           n59120, ZN => n58877);
   U1466 : INV_X1 port map( A => n58877, ZN => n3434);
   U1467 : OAI22_X1 port map( A1 => n52444, A2 => n58897, B1 => n53103, B2 => 
                           n59128, ZN => n58878);
   U1468 : INV_X1 port map( A => n58878, ZN => n3049);
   U1469 : OAI22_X1 port map( A1 => n52454, A2 => n58891, B1 => n53017, B2 => 
                           n59120, ZN => n58879);
   U1470 : INV_X1 port map( A => n58879, ZN => n3498);
   U1471 : OAI22_X1 port map( A1 => n52440, A2 => n58891, B1 => n52490, B2 => 
                           n59152, ZN => n58880);
   U1472 : INV_X1 port map( A => n58880, ZN => n3507);
   U1473 : OAI22_X1 port map( A1 => n52441, A2 => n58887, B1 => n52986, B2 => 
                           n59161, ZN => n58881);
   U1474 : INV_X1 port map( A => n58881, ZN => n3337);
   U1475 : OAI22_X1 port map( A1 => n52441, A2 => n58894, B1 => n53021, B2 => 
                           n59161, ZN => n58882);
   U1476 : INV_X1 port map( A => n58882, ZN => n3403);
   U1477 : OAI22_X1 port map( A1 => n52435, A2 => n58885, B1 => n52949, B2 => 
                           n59164, ZN => n58883);
   U1478 : INV_X1 port map( A => n58883, ZN => n2888);
   U1479 : OAI22_X1 port map( A1 => n52444, A2 => n58894, B1 => n53023, B2 => 
                           n59128, ZN => n58884);
   U1480 : INV_X1 port map( A => n58884, ZN => n3405);
   U1481 : OAI22_X1 port map( A1 => n52438, A2 => n58885, B1 => n52697, B2 => 
                           n59183, ZN => n58886);
   U1482 : INV_X1 port map( A => n58886, ZN => n2901);
   U1483 : OAI22_X1 port map( A1 => n52457, A2 => n58887, B1 => n52635, B2 => 
                           n59156, ZN => n58888);
   U1484 : INV_X1 port map( A => n58888, ZN => n3350);
   U1485 : OAI22_X1 port map( A1 => n52444, A2 => n58891, B1 => n53027, B2 => 
                           n59128, ZN => n58889);
   U1486 : INV_X1 port map( A => n58889, ZN => n3499);
   U1487 : OAI22_X1 port map( A1 => n52435, A2 => n58904, B1 => n52839, B2 => 
                           n59164, ZN => n58890);
   U1488 : INV_X1 port map( A => n58890, ZN => n3239);
   U1489 : OAI22_X1 port map( A1 => n52441, A2 => n58891, B1 => n53029, B2 => 
                           n59161, ZN => n58892);
   U1490 : INV_X1 port map( A => n58892, ZN => n3501);
   U1491 : OAI22_X1 port map( A1 => n52441, A2 => n58906, B1 => n52982, B2 => 
                           n59161, ZN => n58893);
   U1492 : INV_X1 port map( A => n58893, ZN => n3305);
   U1493 : OAI22_X1 port map( A1 => n52440, A2 => n58894, B1 => n52496, B2 => 
                           n59152, ZN => n58895);
   U1494 : INV_X1 port map( A => n58895, ZN => n3411);
   U1495 : OAI22_X1 port map( A1 => n52458, A2 => n58900, B1 => n52623, B2 => 
                           n59006, ZN => n58896);
   U1496 : INV_X1 port map( A => n58896, ZN => n3446);
   U1497 : OAI22_X1 port map( A1 => n52473, A2 => n58897, B1 => n52955, B2 => 
                           n59130, ZN => n58898);
   U1498 : INV_X1 port map( A => n58898, ZN => n3048);
   U1499 : OAI22_X1 port map( A1 => n52456, A2 => n58906, B1 => n52626, B2 => 
                           n58982, ZN => n58899);
   U1500 : INV_X1 port map( A => n58899, ZN => n3315);
   U1501 : OAI22_X1 port map( A1 => n52438, A2 => n58900, B1 => n52507, B2 => 
                           n59183, ZN => n58901);
   U1502 : INV_X1 port map( A => n58901, ZN => n3443);
   U1503 : OAI22_X1 port map( A1 => n52456, A2 => n58902, B1 => n52528, B2 => 
                           n58982, ZN => n58903);
   U1504 : INV_X1 port map( A => n58903, ZN => n2931);
   U1505 : OAI22_X1 port map( A1 => n52478, A2 => n58904, B1 => n52837, B2 => 
                           n58980, ZN => n58905);
   U1506 : INV_X1 port map( A => n58905, ZN => n3238);
   U1507 : OAI22_X1 port map( A1 => n52442, A2 => n58906, B1 => n52983, B2 => 
                           n59168, ZN => n58907);
   U1508 : INV_X1 port map( A => n58907, ZN => n3306);
   U1509 : OAI22_X1 port map( A1 => n52444, A2 => n58908, B1 => n53102, B2 => 
                           n59128, ZN => n58909);
   U1510 : INV_X1 port map( A => n58909, ZN => n3081);
   U1511 : CLKBUF_X1 port map( A => n58910, Z => n58957);
   U1512 : OAI22_X1 port map( A1 => n52453, A2 => n58957, B1 => n52663, B2 => 
                           n59148, ZN => n58911);
   U1513 : INV_X1 port map( A => n58911, ZN => n3386);
   U1514 : CLKBUF_X1 port map( A => n59169, Z => n58952);
   U1515 : OAI22_X1 port map( A1 => n52456, A2 => n58952, B1 => n52672, B2 => 
                           n58982, ZN => n58912);
   U1516 : INV_X1 port map( A => n58912, ZN => n3482);
   U1517 : CLKBUF_X1 port map( A => n58913, Z => n58954);
   U1518 : OAI22_X1 port map( A1 => n52455, A2 => n58954, B1 => n52719, B2 => 
                           n58985, ZN => n58914);
   U1519 : INV_X1 port map( A => n58914, ZN => n2970);
   U1520 : CLKBUF_X1 port map( A => n58915, Z => n58961);
   U1521 : OAI22_X1 port map( A1 => n52458, A2 => n58961, B1 => n52676, B2 => 
                           n59006, ZN => n58916);
   U1522 : INV_X1 port map( A => n58916, ZN => n3290);
   U1523 : CLKBUF_X1 port map( A => n59173, Z => n58959);
   U1524 : OAI22_X1 port map( A1 => n52458, A2 => n58959, B1 => n53262, B2 => 
                           n59006, ZN => n58917);
   U1525 : INV_X1 port map( A => n58917, ZN => n3210);
   U1526 : OAI22_X1 port map( A1 => n52442, A2 => n58957, B1 => n53005, B2 => 
                           n59168, ZN => n58918);
   U1527 : INV_X1 port map( A => n58918, ZN => n3370);
   U1528 : OAI22_X1 port map( A1 => n52439, A2 => n58959, B1 => n53289, B2 => 
                           n59154, ZN => n58919);
   U1529 : INV_X1 port map( A => n58919, ZN => n3213);
   U1530 : OAI22_X1 port map( A1 => n52438, A2 => n58959, B1 => n53288, B2 => 
                           n59183, ZN => n58920);
   U1531 : INV_X1 port map( A => n58920, ZN => n3212);
   U1532 : OAI22_X1 port map( A1 => n52467, A2 => n58954, B1 => n53173, B2 => 
                           n59212, ZN => n58921);
   U1533 : INV_X1 port map( A => n58921, ZN => n2957);
   U1534 : OAI22_X1 port map( A1 => n52450, A2 => n58954, B1 => n53135, B2 => 
                           n59175, ZN => n58922);
   U1535 : INV_X1 port map( A => n58922, ZN => n2953);
   U1536 : OAI22_X1 port map( A1 => n52448, A2 => n58952, B1 => n52994, B2 => 
                           n59171, ZN => n58923);
   U1537 : INV_X1 port map( A => n58923, ZN => n3468);
   U1538 : OAI22_X1 port map( A1 => n52441, A2 => n58952, B1 => n52991, B2 => 
                           n59161, ZN => n58924);
   U1539 : INV_X1 port map( A => n58924, ZN => n3467);
   U1540 : OAI22_X1 port map( A1 => n52457, A2 => n58959, B1 => n53254, B2 => 
                           n59156, ZN => n58925);
   U1541 : INV_X1 port map( A => n58925, ZN => n3209);
   U1542 : OAI22_X1 port map( A1 => n52445, A2 => n58952, B1 => n52990, B2 => 
                           n58967, ZN => n58926);
   U1543 : INV_X1 port map( A => n58926, ZN => n3466);
   U1544 : OAI22_X1 port map( A1 => n52442, A2 => n58961, B1 => n53142, B2 => 
                           n59168, ZN => n58927);
   U1545 : INV_X1 port map( A => n58927, ZN => n3277);
   U1546 : OAI22_X1 port map( A1 => n52444, A2 => n58952, B1 => n52988, B2 => 
                           n59128, ZN => n58928);
   U1547 : INV_X1 port map( A => n58928, ZN => n3465);
   U1548 : OAI22_X1 port map( A1 => n52478, A2 => n58959, B1 => n52892, B2 => 
                           n58980, ZN => n58929);
   U1549 : INV_X1 port map( A => n58929, ZN => n3226);
   U1550 : OAI22_X1 port map( A1 => n52435, A2 => n58957, B1 => n52885, B2 => 
                           n59164, ZN => n58930);
   U1551 : INV_X1 port map( A => n58930, ZN => n3367);
   U1552 : OAI22_X1 port map( A1 => n52445, A2 => n58961, B1 => n53121, B2 => 
                           n58967, ZN => n58931);
   U1553 : INV_X1 port map( A => n58931, ZN => n3275);
   U1554 : OAI22_X1 port map( A1 => n52469, A2 => n58957, B1 => n52941, B2 => 
                           n58996, ZN => n58932);
   U1555 : INV_X1 port map( A => n58932, ZN => n3368);
   U1556 : OAI22_X1 port map( A1 => n52435, A2 => n58952, B1 => n52882, B2 => 
                           n59164, ZN => n58933);
   U1557 : INV_X1 port map( A => n58933, ZN => n3463);
   U1558 : OAI22_X1 port map( A1 => n52445, A2 => n58957, B1 => n53000, B2 => 
                           n58967, ZN => n58934);
   U1559 : INV_X1 port map( A => n58934, ZN => n3369);
   U1560 : OAI22_X1 port map( A1 => n52445, A2 => n58954, B1 => n53169, B2 => 
                           n58967, ZN => n58935);
   U1561 : INV_X1 port map( A => n58935, ZN => n2955);
   U1562 : OAI22_X1 port map( A1 => n52452, A2 => n58959, B1 => n53078, B2 => 
                           n59134, ZN => n58936);
   U1563 : INV_X1 port map( A => n58936, ZN => n3206);
   U1564 : OAI22_X1 port map( A1 => n52469, A2 => n58961, B1 => n52826, B2 => 
                           n58996, ZN => n58937);
   U1565 : INV_X1 port map( A => n58937, ZN => n3270);
   U1566 : OAI22_X1 port map( A1 => n52477, A2 => n58961, B1 => n52827, B2 => 
                           n59126, ZN => n58938);
   U1567 : INV_X1 port map( A => n58938, ZN => n3271);
   U1568 : OAI22_X1 port map( A1 => n52455, A2 => n58959, B1 => n53269, B2 => 
                           n58985, ZN => n58939);
   U1569 : INV_X1 port map( A => n58939, ZN => n3211);
   U1570 : OAI22_X1 port map( A1 => n52454, A2 => n58957, B1 => n53013, B2 => 
                           n59120, ZN => n58940);
   U1571 : INV_X1 port map( A => n58940, ZN => n3373);
   U1572 : OAI22_X1 port map( A1 => n52477, A2 => n58954, B1 => n52965, B2 => 
                           n59126, ZN => n58941);
   U1573 : INV_X1 port map( A => n58941, ZN => n2952);
   U1574 : OAI22_X1 port map( A1 => n52442, A2 => n58954, B1 => n53153, B2 => 
                           n59168, ZN => n58942);
   U1575 : INV_X1 port map( A => n58942, ZN => n2954);
   U1576 : OAI22_X1 port map( A1 => n52469, A2 => n58952, B1 => n52915, B2 => 
                           n58996, ZN => n58943);
   U1577 : INV_X1 port map( A => n58943, ZN => n3464);
   U1578 : OAI22_X1 port map( A1 => n52454, A2 => n58952, B1 => n53016, B2 => 
                           n59120, ZN => n58944);
   U1579 : INV_X1 port map( A => n58944, ZN => n3469);
   U1580 : OAI22_X1 port map( A1 => n52473, A2 => n58961, B1 => n52829, B2 => 
                           n59130, ZN => n58945);
   U1581 : INV_X1 port map( A => n58945, ZN => n3272);
   U1582 : OAI22_X1 port map( A1 => n52469, A2 => n58954, B1 => n52946, B2 => 
                           n58996, ZN => n58946);
   U1583 : INV_X1 port map( A => n58946, ZN => n2951);
   U1584 : OAI22_X1 port map( A1 => n52442, A2 => n58959, B1 => n53116, B2 => 
                           n59168, ZN => n58947);
   U1585 : INV_X1 port map( A => n58947, ZN => n3208);
   U1586 : OAI22_X1 port map( A1 => n52441, A2 => n58954, B1 => n53172, B2 => 
                           n59161, ZN => n58948);
   U1587 : INV_X1 port map( A => n58948, ZN => n2956);
   U1588 : OAI22_X1 port map( A1 => n52448, A2 => n58957, B1 => n53010, B2 => 
                           n59171, ZN => n58949);
   U1589 : INV_X1 port map( A => n58949, ZN => n3372);
   U1590 : OAI22_X1 port map( A1 => n52454, A2 => n58961, B1 => n53088, B2 => 
                           n59120, ZN => n58950);
   U1591 : INV_X1 port map( A => n58950, ZN => n3273);
   U1592 : OAI22_X1 port map( A1 => n52441, A2 => n58957, B1 => n53009, B2 => 
                           n59161, ZN => n58951);
   U1593 : INV_X1 port map( A => n58951, ZN => n3371);
   U1594 : OAI22_X1 port map( A1 => n52436, A2 => n58952, B1 => n52880, B2 => 
                           n59124, ZN => n58953);
   U1595 : INV_X1 port map( A => n58953, ZN => n3462);
   U1596 : OAI22_X1 port map( A1 => n52473, A2 => n58954, B1 => n52945, B2 => 
                           n59130, ZN => n58955);
   U1597 : INV_X1 port map( A => n58955, ZN => n2950);
   U1598 : OAI22_X1 port map( A1 => n52450, A2 => n58961, B1 => n53124, B2 => 
                           n59175, ZN => n58956);
   U1599 : INV_X1 port map( A => n58956, ZN => n3276);
   U1600 : OAI22_X1 port map( A1 => n52436, A2 => n58957, B1 => n52877, B2 => 
                           n59124, ZN => n58958);
   U1601 : INV_X1 port map( A => n58958, ZN => n3366);
   U1602 : OAI22_X1 port map( A1 => n52454, A2 => n58959, B1 => n53090, B2 => 
                           n59120, ZN => n58960);
   U1603 : INV_X1 port map( A => n58960, ZN => n3207);
   U1604 : OAI22_X1 port map( A1 => n52444, A2 => n58961, B1 => n53094, B2 => 
                           n59128, ZN => n58962);
   U1605 : INV_X1 port map( A => n58962, ZN => n3274);
   U1606 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53620, ZN => n59293);
   U1607 : CLKBUF_X1 port map( A => n59293, Z => n59264);
   U1608 : CLKBUF_X1 port map( A => n59120, Z => n59075);
   U1609 : OAI22_X1 port map( A1 => n52454, A2 => n59264, B1 => n53459, B2 => 
                           n59075, ZN => n58963);
   U1610 : INV_X1 port map( A => n58963, ZN => n2571);
   U1611 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53617, ZN => n59279);
   U1612 : CLKBUF_X1 port map( A => n59279, Z => n59310);
   U1613 : CLKBUF_X1 port map( A => n59128, Z => n59116);
   U1614 : OAI22_X1 port map( A1 => n52444, A2 => n59310, B1 => n53460, B2 => 
                           n59116, ZN => n58964);
   U1615 : INV_X1 port map( A => n58964, ZN => n2667);
   U1616 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53619, ZN => n59319);
   U1617 : CLKBUF_X1 port map( A => n59319, Z => n59277);
   U1618 : OAI22_X1 port map( A1 => n52454, A2 => n59277, B1 => n53470, B2 => 
                           n59075, ZN => n58965);
   U1619 : INV_X1 port map( A => n58965, ZN => n2605);
   U1620 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53616, ZN => n59325);
   U1621 : CLKBUF_X1 port map( A => n59325, Z => n59287);
   U1622 : OAI22_X1 port map( A1 => n52454, A2 => n59287, B1 => n53467, B2 => 
                           n59075, ZN => n58966);
   U1623 : INV_X1 port map( A => n58966, ZN => n2698);
   U1624 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53614, ZN => n59312);
   U1625 : CLKBUF_X1 port map( A => n58967, Z => n59114);
   U1626 : OAI22_X1 port map( A1 => n52445, A2 => n59312, B1 => n53501, B2 => 
                           n59114, ZN => n58968);
   U1627 : INV_X1 port map( A => n58968, ZN => n2766);
   U1628 : CLKBUF_X1 port map( A => n59312, Z => n59295);
   U1629 : OAI22_X1 port map( A1 => n52454, A2 => n59295, B1 => n53490, B2 => 
                           n59075, ZN => n58969);
   U1630 : INV_X1 port map( A => n58969, ZN => n2764);
   U1631 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53621, ZN => n59308);
   U1632 : CLKBUF_X1 port map( A => n59308, Z => n59322);
   U1633 : OAI22_X1 port map( A1 => n52445, A2 => n59322, B1 => n53483, B2 => 
                           n59114, ZN => n58970);
   U1634 : INV_X1 port map( A => n58970, ZN => n2541);
   U1635 : OAI22_X1 port map( A1 => n52444, A2 => n59322, B1 => n53481, B2 => 
                           n59116, ZN => n58971);
   U1636 : INV_X1 port map( A => n58971, ZN => n2540);
   U1637 : OAI22_X1 port map( A1 => n52444, A2 => n59295, B1 => n53479, B2 => 
                           n59116, ZN => n58972);
   U1638 : INV_X1 port map( A => n58972, ZN => n2762);
   U1639 : OAI22_X1 port map( A1 => n52454, A2 => n59322, B1 => n53476, B2 => 
                           n59075, ZN => n58973);
   U1640 : INV_X1 port map( A => n58973, ZN => n2538);
   U1641 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53615, ZN => n59255);
   U1642 : CLKBUF_X1 port map( A => n59255, Z => n59328);
   U1643 : OAI22_X1 port map( A1 => n52445, A2 => n59328, B1 => n53472, B2 => 
                           n59114, ZN => n58974);
   U1644 : INV_X1 port map( A => n58974, ZN => n2728);
   U1645 : OAI22_X1 port map( A1 => n52444, A2 => n59328, B1 => n53473, B2 => 
                           n59116, ZN => n58975);
   U1646 : INV_X1 port map( A => n58975, ZN => n2729);
   U1647 : CLKBUF_X1 port map( A => n58976, Z => n59060);
   U1648 : OAI22_X1 port map( A1 => n52449, A2 => n59279, B1 => n53342, B2 => 
                           n59060, ZN => n58977);
   U1649 : INV_X1 port map( A => n58977, ZN => n2685);
   U1650 : CLKBUF_X1 port map( A => n58978, Z => n59040);
   U1651 : OAI22_X1 port map( A1 => n52446, A2 => n59312, B1 => n53340, B2 => 
                           n59040, ZN => n58979);
   U1652 : INV_X1 port map( A => n58979, ZN => n2782);
   U1653 : CLKBUF_X1 port map( A => n58980, Z => n59032);
   U1654 : OAI22_X1 port map( A1 => n52478, A2 => n59322, B1 => n53392, B2 => 
                           n59032, ZN => n58981);
   U1655 : INV_X1 port map( A => n58981, ZN => n2534);
   U1656 : CLKBUF_X1 port map( A => n58982, Z => n59077);
   U1657 : OAI22_X1 port map( A1 => n52456, A2 => n59287, B1 => n53260, B2 => 
                           n59077, ZN => n58983);
   U1658 : INV_X1 port map( A => n58983, ZN => n2708);
   U1659 : OAI22_X1 port map( A1 => n52478, A2 => n59312, B1 => n53397, B2 => 
                           n59032, ZN => n58984);
   U1660 : INV_X1 port map( A => n58984, ZN => n2787);
   U1661 : CLKBUF_X1 port map( A => n58985, Z => n59118);
   U1662 : OAI22_X1 port map( A1 => n52455, A2 => n59279, B1 => n53257, B2 => 
                           n59118, ZN => n58986);
   U1663 : INV_X1 port map( A => n58986, ZN => n2681);
   U1664 : OAI22_X1 port map( A1 => n52449, A2 => n59319, B1 => n53346, B2 => 
                           n59060, ZN => n58987);
   U1665 : INV_X1 port map( A => n58987, ZN => n2619);
   U1666 : OAI22_X1 port map( A1 => n52456, A2 => n59312, B1 => n53261, B2 => 
                           n59077, ZN => n58988);
   U1667 : INV_X1 port map( A => n58988, ZN => n2773);
   U1668 : OAI22_X1 port map( A1 => n52449, A2 => n59293, B1 => n53335, B2 => 
                           n59060, ZN => n58989);
   U1669 : INV_X1 port map( A => n58989, ZN => n2588);
   U1670 : OAI22_X1 port map( A1 => n52455, A2 => n59293, B1 => n53256, B2 => 
                           n59118, ZN => n58990);
   U1671 : INV_X1 port map( A => n58990, ZN => n2584);
   U1672 : OAI22_X1 port map( A1 => n52456, A2 => n59308, B1 => n53253, B2 => 
                           n59077, ZN => n58991);
   U1673 : INV_X1 port map( A => n58991, ZN => n2547);
   U1674 : CLKBUF_X1 port map( A => n59124, Z => n59048);
   U1675 : OAI22_X1 port map( A1 => n52436, A2 => n59319, B1 => n53398, B2 => 
                           n59048, ZN => n58992);
   U1676 : INV_X1 port map( A => n58992, ZN => n2626);
   U1677 : CLKBUF_X1 port map( A => n58993, Z => n59079);
   U1678 : OAI22_X1 port map( A1 => n52459, A2 => n59328, B1 => n53399, B2 => 
                           n59079, ZN => n58994);
   U1679 : INV_X1 port map( A => n58994, ZN => n2727);
   U1680 : OAI22_X1 port map( A1 => n52446, A2 => n59293, B1 => n53190, B2 => 
                           n59040, ZN => n58995);
   U1681 : INV_X1 port map( A => n58995, ZN => n2576);
   U1682 : CLKBUF_X1 port map( A => n58996, Z => n59110);
   U1683 : OAI22_X1 port map( A1 => n52469, A2 => n59322, B1 => n53400, B2 => 
                           n59110, ZN => n58997);
   U1684 : INV_X1 port map( A => n58997, ZN => n2535);
   U1685 : OAI22_X1 port map( A1 => n52469, A2 => n59310, B1 => n53401, B2 => 
                           n59110, ZN => n58998);
   U1686 : INV_X1 port map( A => n58998, ZN => n2663);
   U1687 : CLKBUF_X1 port map( A => n58999, Z => n59073);
   U1688 : OAI22_X1 port map( A1 => n52451, A2 => n59312, B1 => n53248, B2 => 
                           n59073, ZN => n59000);
   U1689 : INV_X1 port map( A => n59000, ZN => n2771);
   U1690 : OAI22_X1 port map( A1 => n52455, A2 => n59319, B1 => n53264, B2 => 
                           n59118, ZN => n59001);
   U1691 : INV_X1 port map( A => n59001, ZN => n2611);
   U1692 : OAI22_X1 port map( A1 => n52455, A2 => n59328, B1 => n53265, B2 => 
                           n59118, ZN => n59002);
   U1693 : INV_X1 port map( A => n59002, ZN => n2746);
   U1694 : OAI22_X1 port map( A1 => n52469, A2 => n59325, B1 => n53404, B2 => 
                           n59110, ZN => n59003);
   U1695 : INV_X1 port map( A => n59003, ZN => n2722);
   U1696 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n53618, ZN => n59267);
   U1697 : OAI22_X1 port map( A1 => n52446, A2 => n59267, B1 => n53195, B2 => 
                           n59040, ZN => n59004);
   U1698 : INV_X1 port map( A => n59004, ZN => n2640);
   U1699 : OAI22_X1 port map( A1 => n52436, A2 => n59264, B1 => n53408, B2 => 
                           n59048, ZN => n59005);
   U1700 : INV_X1 port map( A => n59005, ZN => n2566);
   U1701 : CLKBUF_X1 port map( A => n59006, Z => n59062);
   U1702 : OAI22_X1 port map( A1 => n52458, A2 => n59312, B1 => n53267, B2 => 
                           n59062, ZN => n59007);
   U1703 : INV_X1 port map( A => n59007, ZN => n2774);
   U1704 : OAI22_X1 port map( A1 => n52451, A2 => n59325, B1 => n53324, B2 => 
                           n59073, ZN => n59008);
   U1705 : INV_X1 port map( A => n59008, ZN => n2716);
   U1706 : OAI22_X1 port map( A1 => n52478, A2 => n59319, B1 => n53410, B2 => 
                           n59032, ZN => n59009);
   U1707 : INV_X1 port map( A => n59009, ZN => n2627);
   U1708 : OAI22_X1 port map( A1 => n52455, A2 => n59312, B1 => n53270, B2 => 
                           n59118, ZN => n59010);
   U1709 : INV_X1 port map( A => n59010, ZN => n2775);
   U1710 : OAI22_X1 port map( A1 => n52478, A2 => n59325, B1 => n53412, B2 => 
                           n59032, ZN => n59011);
   U1711 : INV_X1 port map( A => n59011, ZN => n2723);
   U1712 : OAI22_X1 port map( A1 => n52446, A2 => n59325, B1 => n53323, B2 => 
                           n59040, ZN => n59012);
   U1713 : INV_X1 port map( A => n59012, ZN => n2715);
   U1714 : OAI22_X1 port map( A1 => n52449, A2 => n59312, B1 => n53245, B2 => 
                           n59060, ZN => n59013);
   U1715 : INV_X1 port map( A => n59013, ZN => n2770);
   U1716 : OAI22_X1 port map( A1 => n52446, A2 => n59255, B1 => n53205, B2 => 
                           n59040, ZN => n59014);
   U1717 : INV_X1 port map( A => n59014, ZN => n2738);
   U1718 : OAI22_X1 port map( A1 => n52478, A2 => n59255, B1 => n53414, B2 => 
                           n59032, ZN => n59015);
   U1719 : INV_X1 port map( A => n59015, ZN => n2754);
   U1720 : OAI22_X1 port map( A1 => n52459, A2 => n59308, B1 => n53415, B2 => 
                           n59079, ZN => n59016);
   U1721 : INV_X1 port map( A => n59016, ZN => n2563);
   U1722 : OAI22_X1 port map( A1 => n52446, A2 => n59319, B1 => n53353, B2 => 
                           n59040, ZN => n59017);
   U1723 : INV_X1 port map( A => n59017, ZN => n2622);
   U1724 : OAI22_X1 port map( A1 => n52469, A2 => n59255, B1 => n53383, B2 => 
                           n59110, ZN => n59018);
   U1725 : INV_X1 port map( A => n59018, ZN => n2752);
   U1726 : OAI22_X1 port map( A1 => n52449, A2 => n59267, B1 => n53321, B2 => 
                           n59060, ZN => n59019);
   U1727 : INV_X1 port map( A => n59019, ZN => n2654);
   U1728 : OAI22_X1 port map( A1 => n52455, A2 => n59325, B1 => n53272, B2 => 
                           n59118, ZN => n59020);
   U1729 : INV_X1 port map( A => n59020, ZN => n2709);
   U1730 : OAI22_X1 port map( A1 => n52436, A2 => n59279, B1 => n53417, B2 => 
                           n59048, ZN => n59021);
   U1731 : INV_X1 port map( A => n59021, ZN => n2689);
   U1732 : OAI22_X1 port map( A1 => n52478, A2 => n59279, B1 => n53419, B2 => 
                           n59032, ZN => n59022);
   U1733 : INV_X1 port map( A => n59022, ZN => n2690);
   U1734 : OAI22_X1 port map( A1 => n52436, A2 => n59267, B1 => n53422, B2 => 
                           n59048, ZN => n59023);
   U1735 : INV_X1 port map( A => n59023, ZN => n2658);
   U1736 : OAI22_X1 port map( A1 => n52459, A2 => n59267, B1 => n53423, B2 => 
                           n59079, ZN => n59024);
   U1737 : INV_X1 port map( A => n59024, ZN => n2659);
   U1738 : OAI22_X1 port map( A1 => n52469, A2 => n59293, B1 => n53426, B2 => 
                           n59110, ZN => n59025);
   U1739 : INV_X1 port map( A => n59025, ZN => n2594);
   U1740 : OAI22_X1 port map( A1 => n52436, A2 => n59312, B1 => n53427, B2 => 
                           n59048, ZN => n59026);
   U1741 : INV_X1 port map( A => n59026, ZN => n2788);
   U1742 : OAI22_X1 port map( A1 => n52478, A2 => n59267, B1 => n53428, B2 => 
                           n59032, ZN => n59027);
   U1743 : INV_X1 port map( A => n59027, ZN => n2660);
   U1744 : OAI22_X1 port map( A1 => n52458, A2 => n59293, B1 => n53241, B2 => 
                           n59062, ZN => n59028);
   U1745 : INV_X1 port map( A => n59028, ZN => n2582);
   U1746 : OAI22_X1 port map( A1 => n52446, A2 => n59308, B1 => n53315, B2 => 
                           n59040, ZN => n59029);
   U1747 : INV_X1 port map( A => n59029, ZN => n2557);
   U1748 : OAI22_X1 port map( A1 => n52436, A2 => n59255, B1 => n53433, B2 => 
                           n59048, ZN => n59030);
   U1749 : INV_X1 port map( A => n59030, ZN => n2756);
   U1750 : OAI22_X1 port map( A1 => n52449, A2 => n59308, B1 => n53313, B2 => 
                           n59060, ZN => n59031);
   U1751 : INV_X1 port map( A => n59031, ZN => n2555);
   U1752 : OAI22_X1 port map( A1 => n52478, A2 => n59293, B1 => n53434, B2 => 
                           n59032, ZN => n59033);
   U1753 : INV_X1 port map( A => n59033, ZN => n2596);
   U1754 : OAI22_X1 port map( A1 => n52458, A2 => n59279, B1 => n53240, B2 => 
                           n59062, ZN => n59034);
   U1755 : INV_X1 port map( A => n59034, ZN => n2680);
   U1756 : OAI22_X1 port map( A1 => n52458, A2 => n59255, B1 => n53239, B2 => 
                           n59062, ZN => n59035);
   U1757 : INV_X1 port map( A => n59035, ZN => n2744);
   U1758 : OAI22_X1 port map( A1 => n52459, A2 => n59325, B1 => n53382, B2 => 
                           n59079, ZN => n59036);
   U1759 : INV_X1 port map( A => n59036, ZN => n2720);
   U1760 : OAI22_X1 port map( A1 => n52458, A2 => n59325, B1 => n53279, B2 => 
                           n59062, ZN => n59037);
   U1761 : INV_X1 port map( A => n59037, ZN => n2710);
   U1762 : OAI22_X1 port map( A1 => n52445, A2 => n59277, B1 => n53439, B2 => 
                           n59114, ZN => n59038);
   U1763 : INV_X1 port map( A => n59038, ZN => n2602);
   U1764 : OAI22_X1 port map( A1 => n52456, A2 => n59319, B1 => n53282, B2 => 
                           n59077, ZN => n59039);
   U1765 : INV_X1 port map( A => n59039, ZN => n2613);
   U1766 : OAI22_X1 port map( A1 => n52446, A2 => n59279, B1 => n53191, B2 => 
                           n59040, ZN => n59041);
   U1767 : INV_X1 port map( A => n59041, ZN => n2672);
   U1768 : OAI22_X1 port map( A1 => n52469, A2 => n59277, B1 => n53380, B2 => 
                           n59110, ZN => n59042);
   U1769 : INV_X1 port map( A => n59042, ZN => n2599);
   U1770 : OAI22_X1 port map( A1 => n52454, A2 => n59267, B1 => n53442, B2 => 
                           n59075, ZN => n59043);
   U1771 : INV_X1 port map( A => n59043, ZN => n2661);
   U1772 : OAI22_X1 port map( A1 => n52444, A2 => n59287, B1 => n53443, B2 => 
                           n59116, ZN => n59044);
   U1773 : INV_X1 port map( A => n59044, ZN => n2700);
   U1774 : OAI22_X1 port map( A1 => n52458, A2 => n59319, B1 => n53283, B2 => 
                           n59062, ZN => n59045);
   U1775 : INV_X1 port map( A => n59045, ZN => n2614);
   U1776 : OAI22_X1 port map( A1 => n52436, A2 => n59308, B1 => n53377, B2 => 
                           n59048, ZN => n59046);
   U1777 : INV_X1 port map( A => n59046, ZN => n2560);
   U1778 : OAI22_X1 port map( A1 => n52454, A2 => n59255, B1 => n53458, B2 => 
                           n59075, ZN => n59047);
   U1779 : INV_X1 port map( A => n59047, ZN => n2757);
   U1780 : OAI22_X1 port map( A1 => n52436, A2 => n59325, B1 => n53379, B2 => 
                           n59048, ZN => n59049);
   U1781 : INV_X1 port map( A => n59049, ZN => n2719);
   U1782 : OAI22_X1 port map( A1 => n52445, A2 => n59287, B1 => n53445, B2 => 
                           n59114, ZN => n59050);
   U1783 : INV_X1 port map( A => n59050, ZN => n2699);
   U1784 : OAI22_X1 port map( A1 => n52444, A2 => n59277, B1 => n53446, B2 => 
                           n59116, ZN => n59051);
   U1785 : INV_X1 port map( A => n59051, ZN => n2603);
   U1786 : OAI22_X1 port map( A1 => n52445, A2 => n59279, B1 => n53447, B2 => 
                           n59114, ZN => n59052);
   U1787 : INV_X1 port map( A => n59052, ZN => n2693);
   U1788 : OAI22_X1 port map( A1 => n52456, A2 => n59293, B1 => n53231, B2 => 
                           n59077, ZN => n59053);
   U1789 : INV_X1 port map( A => n59053, ZN => n2580);
   U1790 : OAI22_X1 port map( A1 => n52458, A2 => n59308, B1 => n53287, B2 => 
                           n59062, ZN => n59054);
   U1791 : INV_X1 port map( A => n59054, ZN => n2550);
   U1792 : OAI22_X1 port map( A1 => n52451, A2 => n59322, B1 => n53305, B2 => 
                           n59073, ZN => n59055);
   U1793 : INV_X1 port map( A => n59055, ZN => n2554);
   U1794 : OAI22_X1 port map( A1 => n52455, A2 => n59308, B1 => n53304, B2 => 
                           n59118, ZN => n59056);
   U1795 : INV_X1 port map( A => n59056, ZN => n2553);
   U1796 : OAI22_X1 port map( A1 => n52449, A2 => n59325, B1 => n53303, B2 => 
                           n59060, ZN => n59057);
   U1797 : INV_X1 port map( A => n59057, ZN => n2713);
   U1798 : OAI22_X1 port map( A1 => n52451, A2 => n59319, B1 => n53307, B2 => 
                           n59073, ZN => n59058);
   U1799 : INV_X1 port map( A => n59058, ZN => n2617);
   U1800 : OAI22_X1 port map( A1 => n52456, A2 => n59279, B1 => n53229, B2 => 
                           n59077, ZN => n59059);
   U1801 : INV_X1 port map( A => n59059, ZN => n2678);
   U1802 : OAI22_X1 port map( A1 => n52449, A2 => n59255, B1 => n53297, B2 => 
                           n59060, ZN => n59061);
   U1803 : INV_X1 port map( A => n59061, ZN => n2749);
   U1804 : OAI22_X1 port map( A1 => n52458, A2 => n59267, B1 => n53223, B2 => 
                           n59062, ZN => n59063);
   U1805 : INV_X1 port map( A => n59063, ZN => n2645);
   U1806 : OAI22_X1 port map( A1 => n52459, A2 => n59293, B1 => n53374, B2 => 
                           n59079, ZN => n59064);
   U1807 : INV_X1 port map( A => n59064, ZN => n2591);
   U1808 : OAI22_X1 port map( A1 => n52456, A2 => n59267, B1 => n53230, B2 => 
                           n59077, ZN => n59065);
   U1809 : INV_X1 port map( A => n59065, ZN => n2647);
   U1810 : OAI22_X1 port map( A1 => n52451, A2 => n59310, B1 => n53311, B2 => 
                           n59073, ZN => n59066);
   U1811 : INV_X1 port map( A => n59066, ZN => n2682);
   U1812 : OAI22_X1 port map( A1 => n52451, A2 => n59267, B1 => n53309, B2 => 
                           n59073, ZN => n59067);
   U1813 : INV_X1 port map( A => n59067, ZN => n2652);
   U1814 : OAI22_X1 port map( A1 => n52459, A2 => n59319, B1 => n53373, B2 => 
                           n59079, ZN => n59068);
   U1815 : INV_X1 port map( A => n59068, ZN => n2623);
   U1816 : OAI22_X1 port map( A1 => n52459, A2 => n59279, B1 => n53376, B2 => 
                           n59079, ZN => n59069);
   U1817 : INV_X1 port map( A => n59069, ZN => n2687);
   U1818 : OAI22_X1 port map( A1 => n52469, A2 => n59295, B1 => n53363, B2 => 
                           n59110, ZN => n59070);
   U1819 : INV_X1 port map( A => n59070, ZN => n2758);
   U1820 : OAI22_X1 port map( A1 => n52444, A2 => n59264, B1 => n53457, B2 => 
                           n59116, ZN => n59071);
   U1821 : INV_X1 port map( A => n59071, ZN => n2570);
   U1822 : OAI22_X1 port map( A1 => n52451, A2 => n59255, B1 => n53294, B2 => 
                           n59073, ZN => n59072);
   U1823 : INV_X1 port map( A => n59072, ZN => n2747);
   U1824 : OAI22_X1 port map( A1 => n52451, A2 => n59293, B1 => n53306, B2 => 
                           n59073, ZN => n59074);
   U1825 : INV_X1 port map( A => n59074, ZN => n2585);
   U1826 : OAI22_X1 port map( A1 => n52454, A2 => n59310, B1 => n53453, B2 => 
                           n59075, ZN => n59076);
   U1827 : INV_X1 port map( A => n59076, ZN => n2665);
   U1828 : OAI22_X1 port map( A1 => n52456, A2 => n59255, B1 => n53224, B2 => 
                           n59077, ZN => n59078);
   U1829 : INV_X1 port map( A => n59078, ZN => n2741);
   U1830 : OAI22_X1 port map( A1 => n52459, A2 => n59312, B1 => n53369, B2 => 
                           n59079, ZN => n59080);
   U1831 : INV_X1 port map( A => n59080, ZN => n2784);
   U1832 : OAI22_X1 port map( A1 => n52445, A2 => n59264, B1 => n53456, B2 => 
                           n59114, ZN => n59081);
   U1833 : INV_X1 port map( A => n59081, ZN => n2569);
   U1834 : CLKBUF_X1 port map( A => n59082, Z => n59108);
   U1835 : OAI22_X1 port map( A1 => n52468, A2 => n59293, B1 => n53429, B2 => 
                           n59108, ZN => n59083);
   U1836 : INV_X1 port map( A => n59083, ZN => n2595);
   U1837 : OAI22_X1 port map( A1 => n52468, A2 => n59277, B1 => n53378, B2 => 
                           n59108, ZN => n59084);
   U1838 : INV_X1 port map( A => n59084, ZN => n2598);
   U1839 : CLKBUF_X1 port map( A => n59130, Z => n59106);
   U1840 : OAI22_X1 port map( A1 => n52473, A2 => n59319, B1 => n53381, B2 => 
                           n59106, ZN => n59085);
   U1841 : INV_X1 port map( A => n59085, ZN => n2624);
   U1842 : CLKBUF_X1 port map( A => n59126, Z => n59102);
   U1843 : OAI22_X1 port map( A1 => n52477, A2 => n59279, B1 => n53431, B2 => 
                           n59102, ZN => n59086);
   U1844 : INV_X1 port map( A => n59086, ZN => n2691);
   U1845 : OAI22_X1 port map( A1 => n52473, A2 => n59293, B1 => n53407, B2 => 
                           n59106, ZN => n59087);
   U1846 : INV_X1 port map( A => n59087, ZN => n2592);
   U1847 : OAI22_X1 port map( A1 => n52473, A2 => n59308, B1 => n53406, B2 => 
                           n59106, ZN => n59088);
   U1848 : INV_X1 port map( A => n59088, ZN => n2562);
   U1849 : OAI22_X1 port map( A1 => n52477, A2 => n59319, B1 => n53411, B2 => 
                           n59102, ZN => n59089);
   U1850 : INV_X1 port map( A => n59089, ZN => n2628);
   U1851 : OAI22_X1 port map( A1 => n52473, A2 => n59325, B1 => n53403, B2 => 
                           n59106, ZN => n59090);
   U1852 : INV_X1 port map( A => n59090, ZN => n2721);
   U1853 : OAI22_X1 port map( A1 => n52477, A2 => n59325, B1 => n53395, B2 => 
                           n59102, ZN => n59091);
   U1854 : INV_X1 port map( A => n59091, ZN => n2702);
   U1855 : OAI22_X1 port map( A1 => n52468, A2 => n59325, B1 => n53413, B2 => 
                           n59108, ZN => n59092);
   U1856 : INV_X1 port map( A => n59092, ZN => n2724);
   U1857 : OAI22_X1 port map( A1 => n52468, A2 => n59312, B1 => n53371, B2 => 
                           n59108, ZN => n59093);
   U1858 : INV_X1 port map( A => n59093, ZN => n2785);
   U1859 : OAI22_X1 port map( A1 => n52468, A2 => n59308, B1 => n53418, B2 => 
                           n59108, ZN => n59094);
   U1860 : INV_X1 port map( A => n59094, ZN => n2564);
   U1861 : OAI22_X1 port map( A1 => n52477, A2 => n59312, B1 => n53355, B2 => 
                           n59102, ZN => n59095);
   U1862 : INV_X1 port map( A => n59095, ZN => n2783);
   U1863 : OAI22_X1 port map( A1 => n52473, A2 => n59267, B1 => n53365, B2 => 
                           n59106, ZN => n59096);
   U1864 : INV_X1 port map( A => n59096, ZN => n2655);
   U1865 : OAI22_X1 port map( A1 => n52477, A2 => n59267, B1 => n53420, B2 => 
                           n59102, ZN => n59097);
   U1866 : INV_X1 port map( A => n59097, ZN => n2657);
   U1867 : OAI22_X1 port map( A1 => n52477, A2 => n59264, B1 => n53409, B2 => 
                           n59102, ZN => n59098);
   U1868 : INV_X1 port map( A => n59098, ZN => n2567);
   U1869 : OAI22_X1 port map( A1 => n52473, A2 => n59310, B1 => n53396, B2 => 
                           n59106, ZN => n59099);
   U1870 : INV_X1 port map( A => n59099, ZN => n2662);
   U1871 : OAI22_X1 port map( A1 => n52468, A2 => n59328, B1 => n53393, B2 => 
                           n59108, ZN => n59100);
   U1872 : INV_X1 port map( A => n59100, ZN => n2726);
   U1873 : OAI22_X1 port map( A1 => n52477, A2 => n59308, B1 => n53405, B2 => 
                           n59102, ZN => n59101);
   U1874 : INV_X1 port map( A => n59101, ZN => n2561);
   U1875 : OAI22_X1 port map( A1 => n52477, A2 => n59255, B1 => n53430, B2 => 
                           n59102, ZN => n59103);
   U1876 : INV_X1 port map( A => n59103, ZN => n2755);
   U1877 : OAI22_X1 port map( A1 => n52468, A2 => n59279, B1 => n53391, B2 => 
                           n59108, ZN => n59104);
   U1878 : INV_X1 port map( A => n59104, ZN => n2688);
   U1879 : OAI22_X1 port map( A1 => n52473, A2 => n59255, B1 => n53368, B2 => 
                           n59106, ZN => n59105);
   U1880 : INV_X1 port map( A => n59105, ZN => n2751);
   U1881 : OAI22_X1 port map( A1 => n52473, A2 => n59295, B1 => n53366, B2 => 
                           n59106, ZN => n59107);
   U1882 : INV_X1 port map( A => n59107, ZN => n2759);
   U1883 : OAI22_X1 port map( A1 => n52468, A2 => n59267, B1 => n53367, B2 => 
                           n59108, ZN => n59109);
   U1884 : INV_X1 port map( A => n59109, ZN => n2656);
   U1885 : CLKBUF_X1 port map( A => n59267, Z => n59302);
   U1886 : OAI22_X1 port map( A1 => n52469, A2 => n59302, B1 => n53364, B2 => 
                           n59110, ZN => n59111);
   U1887 : INV_X1 port map( A => n59111, ZN => n2630);
   U1888 : CLKBUF_X1 port map( A => n59112, Z => n59132);
   U1889 : OAI22_X1 port map( A1 => n52447, A2 => n59132, B1 => n52701, B2 => 
                           n59144, ZN => n59113);
   U1890 : INV_X1 port map( A => n59113, ZN => n3034);
   U1891 : OAI22_X1 port map( A1 => n52445, A2 => n59302, B1 => n53451, B2 => 
                           n59114, ZN => n59115);
   U1892 : INV_X1 port map( A => n59115, ZN => n2633);
   U1893 : OAI22_X1 port map( A1 => n52444, A2 => n59302, B1 => n53455, B2 => 
                           n59116, ZN => n59117);
   U1894 : INV_X1 port map( A => n59117, ZN => n2635);
   U1895 : OAI22_X1 port map( A1 => n52455, A2 => n59302, B1 => n53273, B2 => 
                           n59118, ZN => n59119);
   U1896 : INV_X1 port map( A => n59119, ZN => n2650);
   U1897 : OAI22_X1 port map( A1 => n52454, A2 => n59132, B1 => n53061, B2 => 
                           n59120, ZN => n59121);
   U1898 : INV_X1 port map( A => n59121, ZN => n3020);
   U1899 : OAI22_X1 port map( A1 => n52452, A2 => n59132, B1 => n53060, B2 => 
                           n59134, ZN => n59122);
   U1900 : INV_X1 port map( A => n59122, ZN => n3019);
   U1901 : OAI22_X1 port map( A1 => n52450, A2 => n59132, B1 => n53058, B2 => 
                           n59175, ZN => n59123);
   U1902 : INV_X1 port map( A => n59123, ZN => n3017);
   U1903 : OAI22_X1 port map( A1 => n52436, A2 => n59132, B1 => n52847, B2 => 
                           n59124, ZN => n59125);
   U1904 : INV_X1 port map( A => n59125, ZN => n3016);
   U1905 : OAI22_X1 port map( A1 => n52477, A2 => n59132, B1 => n52801, B2 => 
                           n59126, ZN => n59127);
   U1906 : INV_X1 port map( A => n59127, ZN => n3015);
   U1907 : OAI22_X1 port map( A1 => n52444, A2 => n59132, B1 => n53059, B2 => 
                           n59128, ZN => n59129);
   U1908 : INV_X1 port map( A => n59129, ZN => n3018);
   U1909 : OAI22_X1 port map( A1 => n52473, A2 => n59132, B1 => n52800, B2 => 
                           n59130, ZN => n59131);
   U1910 : INV_X1 port map( A => n59131, ZN => n3014);
   U1911 : OAI22_X1 port map( A1 => n52467, A2 => n59132, B1 => n53174, B2 => 
                           n59212, ZN => n59133);
   U1912 : INV_X1 port map( A => n59133, ZN => n3021);
   U1913 : CLKBUF_X1 port map( A => n59134, Z => n59142);
   U1914 : OAI22_X1 port map( A1 => n52452, A2 => n59322, B1 => n53475, B2 => 
                           n59142, ZN => n59135);
   U1915 : INV_X1 port map( A => n59135, ZN => n2537);
   U1916 : OAI22_X1 port map( A1 => n52452, A2 => n59302, B1 => n53466, B2 => 
                           n59142, ZN => n59136);
   U1917 : INV_X1 port map( A => n59136, ZN => n2636);
   U1918 : OAI22_X1 port map( A1 => n52452, A2 => n59264, B1 => n53463, B2 => 
                           n59142, ZN => n59137);
   U1919 : INV_X1 port map( A => n59137, ZN => n2572);
   U1920 : OAI22_X1 port map( A1 => n52452, A2 => n59310, B1 => n53468, B2 => 
                           n59142, ZN => n59138);
   U1921 : INV_X1 port map( A => n59138, ZN => n2668);
   U1922 : OAI22_X1 port map( A1 => n52452, A2 => n59277, B1 => n53464, B2 => 
                           n59142, ZN => n59139);
   U1923 : INV_X1 port map( A => n59139, ZN => n2604);
   U1924 : OAI22_X1 port map( A1 => n52452, A2 => n59287, B1 => n53469, B2 => 
                           n59142, ZN => n59140);
   U1925 : INV_X1 port map( A => n59140, ZN => n2697);
   U1926 : OAI22_X1 port map( A1 => n52452, A2 => n59295, B1 => n53486, B2 => 
                           n59142, ZN => n59141);
   U1927 : INV_X1 port map( A => n59141, ZN => n2763);
   U1928 : OAI22_X1 port map( A1 => n52452, A2 => n59328, B1 => n53484, B2 => 
                           n59142, ZN => n59143);
   U1929 : INV_X1 port map( A => n59143, ZN => n2731);
   U1930 : CLKBUF_X1 port map( A => n59144, Z => n59314);
   U1931 : OAI22_X1 port map( A1 => n52447, A2 => n59255, B1 => n53296, B2 => 
                           n59314, ZN => n59145);
   U1932 : INV_X1 port map( A => n59145, ZN => n2748);
   U1933 : CLKBUF_X1 port map( A => n59146, Z => n59324);
   U1934 : OAI22_X1 port map( A1 => n52463, A2 => n59319, B1 => n53293, B2 => 
                           n59324, ZN => n59147);
   U1935 : INV_X1 port map( A => n59147, ZN => n2615);
   U1936 : CLKBUF_X1 port map( A => n59148, Z => n59305);
   U1937 : OAI22_X1 port map( A1 => n52453, A2 => n59325, B1 => n53298, B2 => 
                           n59305, ZN => n59149);
   U1938 : INV_X1 port map( A => n59149, ZN => n2712);
   U1939 : CLKBUF_X1 port map( A => n59150, Z => n59297);
   U1940 : OAI22_X1 port map( A1 => n52437, A2 => n59209, B1 => n52586, B2 => 
                           n59297, ZN => n59151);
   U1941 : INV_X1 port map( A => n59151, ZN => n3540);
   U1942 : CLKBUF_X1 port map( A => n59152, Z => n59284);
   U1943 : OAI22_X1 port map( A1 => n52440, A2 => n59209, B1 => n52504, B2 => 
                           n59284, ZN => n59153);
   U1944 : INV_X1 port map( A => n59153, ZN => n3537);
   U1945 : CLKBUF_X1 port map( A => n59154, Z => n59269);
   U1946 : OAI22_X1 port map( A1 => n52439, A2 => n59209, B1 => n52510, B2 => 
                           n59269, ZN => n59155);
   U1947 : INV_X1 port map( A => n59155, ZN => n3538);
   U1948 : CLKBUF_X1 port map( A => n59156, Z => n59318);
   U1949 : OAI22_X1 port map( A1 => n52457, A2 => n59213, B1 => n52516, B2 => 
                           n59318, ZN => n59157);
   U1950 : INV_X1 port map( A => n59157, ZN => n3186);
   U1951 : CLKBUF_X1 port map( A => n59158, Z => n59299);
   U1952 : OAI22_X1 port map( A1 => n52443, A2 => n59267, B1 => n53299, B2 => 
                           n59299, ZN => n59159);
   U1953 : INV_X1 port map( A => n59159, ZN => n2651);
   U1954 : OAI22_X1 port map( A1 => n52453, A2 => n59213, B1 => n52593, B2 => 
                           n59305, ZN => n59160);
   U1955 : INV_X1 port map( A => n59160, ZN => n3193);
   U1956 : CLKBUF_X1 port map( A => n59161, Z => n59327);
   U1957 : OAI22_X1 port map( A1 => n52441, A2 => n59308, B1 => n53461, B2 => 
                           n59327, ZN => n59162);
   U1958 : INV_X1 port map( A => n59162, ZN => n2565);
   U1959 : OAI22_X1 port map( A1 => n52447, A2 => n59213, B1 => n52775, B2 => 
                           n59314, ZN => n59163);
   U1960 : INV_X1 port map( A => n59163, ZN => n3199);
   U1961 : CLKBUF_X1 port map( A => n59164, Z => n59244);
   U1962 : OAI22_X1 port map( A1 => n52435, A2 => n59213, B1 => n52840, B2 => 
                           n59244, ZN => n59165);
   U1963 : INV_X1 port map( A => n59165, ZN => n3203);
   U1964 : OAI22_X1 port map( A1 => n52463, A2 => n59166, B1 => n52714, B2 => 
                           n59324, ZN => n59167);
   U1965 : INV_X1 port map( A => n59167, ZN => n3322);
   U1966 : CLKBUF_X1 port map( A => n59168, Z => n59321);
   U1967 : OAI22_X1 port map( A1 => n52442, A2 => n59169, B1 => n52987, B2 => 
                           n59321, ZN => n59170);
   U1968 : INV_X1 port map( A => n59170, ZN => n3493);
   U1969 : CLKBUF_X1 port map( A => n59171, Z => n59286);
   U1970 : OAI22_X1 port map( A1 => n52448, A2 => n59213, B1 => n53069, B2 => 
                           n59286, ZN => n59172);
   U1971 : INV_X1 port map( A => n59172, ZN => n3205);
   U1972 : OAI22_X1 port map( A1 => n52441, A2 => n59173, B1 => n53118, B2 => 
                           n59327, ZN => n59174);
   U1973 : INV_X1 port map( A => n59174, ZN => n3233);
   U1974 : CLKBUF_X1 port map( A => n59175, Z => n59301);
   U1975 : OAI22_X1 port map( A1 => n52450, A2 => n59213, B1 => n53128, B2 => 
                           n59301, ZN => n59176);
   U1976 : INV_X1 port map( A => n59176, ZN => n3183);
   U1977 : OAI22_X1 port map( A1 => n52443, A2 => n59213, B1 => n52761, B2 => 
                           n59299, ZN => n59177);
   U1978 : INV_X1 port map( A => n59177, ZN => n3197);
   U1979 : OAI22_X1 port map( A1 => n52440, A2 => n59319, B1 => n53222, B2 => 
                           n59284, ZN => n59178);
   U1980 : INV_X1 port map( A => n59178, ZN => n2610);
   U1981 : OAI22_X1 port map( A1 => n52440, A2 => n59325, B1 => n53221, B2 => 
                           n59284, ZN => n59179);
   U1982 : INV_X1 port map( A => n59179, ZN => n2706);
   U1983 : OAI22_X1 port map( A1 => n52437, A2 => n59293, B1 => n53220, B2 => 
                           n59297, ZN => n59180);
   U1984 : INV_X1 port map( A => n59180, ZN => n2578);
   U1985 : OAI22_X1 port map( A1 => n52437, A2 => n59267, B1 => n53219, B2 => 
                           n59297, ZN => n59181);
   U1986 : INV_X1 port map( A => n59181, ZN => n2644);
   U1987 : OAI22_X1 port map( A1 => n52437, A2 => n59255, B1 => n53218, B2 => 
                           n59297, ZN => n59182);
   U1988 : INV_X1 port map( A => n59182, ZN => n2740);
   U1989 : CLKBUF_X1 port map( A => n59183, Z => n59307);
   U1990 : OAI22_X1 port map( A1 => n52438, A2 => n59279, B1 => n53217, B2 => 
                           n59307, ZN => n59184);
   U1991 : INV_X1 port map( A => n59184, ZN => n2676);
   U1992 : OAI22_X1 port map( A1 => n52438, A2 => n59312, B1 => n53216, B2 => 
                           n59307, ZN => n59185);
   U1993 : INV_X1 port map( A => n59185, ZN => n2769);
   U1994 : OAI22_X1 port map( A1 => n52438, A2 => n59325, B1 => n53215, B2 => 
                           n59307, ZN => n59186);
   U1995 : INV_X1 port map( A => n59186, ZN => n2705);
   U1996 : OAI22_X1 port map( A1 => n52437, A2 => n59308, B1 => n53225, B2 => 
                           n59297, ZN => n59187);
   U1997 : INV_X1 port map( A => n59187, ZN => n2545);
   U1998 : OAI22_X1 port map( A1 => n52435, A2 => n59325, B1 => n53385, B2 => 
                           n59244, ZN => n59188);
   U1999 : INV_X1 port map( A => n59188, ZN => n2703);
   U2000 : OAI22_X1 port map( A1 => n52439, A2 => n59319, B1 => n53213, B2 => 
                           n59269, ZN => n59189);
   U2001 : INV_X1 port map( A => n59189, ZN => n2609);
   U2002 : OAI22_X1 port map( A1 => n52438, A2 => n59319, B1 => n53212, B2 => 
                           n59307, ZN => n59190);
   U2003 : INV_X1 port map( A => n59190, ZN => n2608);
   U2004 : OAI22_X1 port map( A1 => n52439, A2 => n59293, B1 => n53226, B2 => 
                           n59269, ZN => n59191);
   U2005 : INV_X1 port map( A => n59191, ZN => n2579);
   U2006 : OAI22_X1 port map( A1 => n52439, A2 => n59267, B1 => n53227, B2 => 
                           n59269, ZN => n59192);
   U2007 : INV_X1 port map( A => n59192, ZN => n2646);
   U2008 : OAI22_X1 port map( A1 => n52435, A2 => n59312, B1 => n53386, B2 => 
                           n59244, ZN => n59193);
   U2009 : INV_X1 port map( A => n59193, ZN => n2786);
   U2010 : OAI22_X1 port map( A1 => n52439, A2 => n59325, B1 => n53210, B2 => 
                           n59269, ZN => n59194);
   U2011 : INV_X1 port map( A => n59194, ZN => n2704);
   U2012 : OAI22_X1 port map( A1 => n52453, A2 => n59279, B1 => n53209, B2 => 
                           n59305, ZN => n59195);
   U2013 : INV_X1 port map( A => n59195, ZN => n2675);
   U2014 : OAI22_X1 port map( A1 => n52439, A2 => n59312, B1 => n53208, B2 => 
                           n59269, ZN => n59196);
   U2015 : INV_X1 port map( A => n59196, ZN => n2768);
   U2016 : OAI22_X1 port map( A1 => n52463, A2 => n59279, B1 => n53207, B2 => 
                           n59324, ZN => n59197);
   U2017 : INV_X1 port map( A => n59197, ZN => n2674);
   U2018 : OAI22_X1 port map( A1 => n52440, A2 => n59255, B1 => n53206, B2 => 
                           n59284, ZN => n59198);
   U2019 : INV_X1 port map( A => n59198, ZN => n2739);
   U2020 : OAI22_X1 port map( A1 => n52463, A2 => n59255, B1 => n53204, B2 => 
                           n59324, ZN => n59199);
   U2021 : INV_X1 port map( A => n59199, ZN => n2737);
   U2022 : OAI22_X1 port map( A1 => n52463, A2 => n59308, B1 => n53202, B2 => 
                           n59324, ZN => n59200);
   U2023 : INV_X1 port map( A => n59200, ZN => n2544);
   U2024 : OAI22_X1 port map( A1 => n52463, A2 => n59267, B1 => n53199, B2 => 
                           n59324, ZN => n59201);
   U2025 : INV_X1 port map( A => n59201, ZN => n2643);
   U2026 : OAI22_X1 port map( A1 => n52448, A2 => n59295, B1 => n53462, B2 => 
                           n59286, ZN => n59202);
   U2027 : INV_X1 port map( A => n59202, ZN => n2760);
   U2028 : OAI22_X1 port map( A1 => n52440, A2 => n59267, B1 => n53198, B2 => 
                           n59284, ZN => n59203);
   U2029 : INV_X1 port map( A => n59203, ZN => n2642);
   U2030 : OAI22_X1 port map( A1 => n52453, A2 => n59267, B1 => n53197, B2 => 
                           n59305, ZN => n59204);
   U2031 : INV_X1 port map( A => n59204, ZN => n2641);
   U2032 : OAI22_X1 port map( A1 => n52440, A2 => n59279, B1 => n53194, B2 => 
                           n59284, ZN => n59205);
   U2033 : INV_X1 port map( A => n59205, ZN => n2673);
   U2034 : OAI22_X1 port map( A1 => n52439, A2 => n59279, B1 => n53228, B2 => 
                           n59269, ZN => n59206);
   U2035 : INV_X1 port map( A => n59206, ZN => n2677);
   U2036 : OAI22_X1 port map( A1 => n52453, A2 => n59293, B1 => n53193, B2 => 
                           n59305, ZN => n59207);
   U2037 : INV_X1 port map( A => n59207, ZN => n2577);
   U2038 : OAI22_X1 port map( A1 => n52453, A2 => n59255, B1 => n53192, B2 => 
                           n59305, ZN => n59208);
   U2039 : INV_X1 port map( A => n59208, ZN => n2736);
   U2040 : OAI22_X1 port map( A1 => n52438, A2 => n59209, B1 => n53189, B2 => 
                           n59307, ZN => n59210);
   U2041 : INV_X1 port map( A => n59210, ZN => n3536);
   U2042 : OAI22_X1 port map( A1 => n52435, A2 => n59255, B1 => n53402, B2 => 
                           n59244, ZN => n59211);
   U2043 : INV_X1 port map( A => n59211, ZN => n2753);
   U2044 : CLKBUF_X1 port map( A => n59212, Z => n59316);
   U2045 : OAI22_X1 port map( A1 => n52467, A2 => n59213, B1 => n53175, B2 => 
                           n59316, ZN => n59214);
   U2046 : INV_X1 port map( A => n59214, ZN => n3184);
   U2047 : OAI22_X1 port map( A1 => n52435, A2 => n59302, B1 => n53416, B2 => 
                           n59244, ZN => n59215);
   U2048 : INV_X1 port map( A => n59215, ZN => n2631);
   U2049 : OAI22_X1 port map( A1 => n52435, A2 => n59293, B1 => n53424, B2 => 
                           n59244, ZN => n59216);
   U2050 : INV_X1 port map( A => n59216, ZN => n2593);
   U2051 : OAI22_X1 port map( A1 => n52435, A2 => n59279, B1 => n53432, B2 => 
                           n59244, ZN => n59217);
   U2052 : INV_X1 port map( A => n59217, ZN => n2692);
   U2053 : OAI22_X1 port map( A1 => n52467, A2 => n59312, B1 => n53435, B2 => 
                           n59316, ZN => n59218);
   U2054 : INV_X1 port map( A => n59218, ZN => n2789);
   U2055 : OAI22_X1 port map( A1 => n52442, A2 => n59319, B1 => n53436, B2 => 
                           n59321, ZN => n59219);
   U2056 : INV_X1 port map( A => n59219, ZN => n2629);
   U2057 : OAI22_X1 port map( A1 => n52441, A2 => n59277, B1 => n53437, B2 => 
                           n59327, ZN => n59220);
   U2058 : INV_X1 port map( A => n59220, ZN => n2600);
   U2059 : OAI22_X1 port map( A1 => n52450, A2 => n59277, B1 => n53438, B2 => 
                           n59301, ZN => n59221);
   U2060 : INV_X1 port map( A => n59221, ZN => n2601);
   U2061 : OAI22_X1 port map( A1 => n52441, A2 => n59325, B1 => n53440, B2 => 
                           n59327, ZN => n59222);
   U2062 : INV_X1 port map( A => n59222, ZN => n2725);
   U2063 : OAI22_X1 port map( A1 => n52442, A2 => n59287, B1 => n53441, B2 => 
                           n59321, ZN => n59223);
   U2064 : INV_X1 port map( A => n59223, ZN => n2701);
   U2065 : OAI22_X1 port map( A1 => n52439, A2 => n59255, B1 => n53233, B2 => 
                           n59269, ZN => n59224);
   U2066 : INV_X1 port map( A => n59224, ZN => n2742);
   U2067 : OAI22_X1 port map( A1 => n52441, A2 => n59302, B1 => n53444, B2 => 
                           n59327, ZN => n59225);
   U2068 : INV_X1 port map( A => n59225, ZN => n2632);
   U2069 : OAI22_X1 port map( A1 => n52467, A2 => n59255, B1 => n53506, B2 => 
                           n59316, ZN => n59226);
   U2070 : INV_X1 port map( A => n59226, ZN => n2735);
   U2071 : OAI22_X1 port map( A1 => n52467, A2 => n59279, B1 => n53505, B2 => 
                           n59316, ZN => n59227);
   U2072 : INV_X1 port map( A => n59227, ZN => n2671);
   U2073 : OAI22_X1 port map( A1 => n52448, A2 => n59319, B1 => n53504, B2 => 
                           n59286, ZN => n59228);
   U2074 : INV_X1 port map( A => n59228, ZN => n2607);
   U2075 : OAI22_X1 port map( A1 => n52442, A2 => n59312, B1 => n53503, B2 => 
                           n59321, ZN => n59229);
   U2076 : INV_X1 port map( A => n59229, ZN => n2767);
   U2077 : OAI22_X1 port map( A1 => n52448, A2 => n59267, B1 => n53502, B2 => 
                           n59286, ZN => n59230);
   U2078 : INV_X1 port map( A => n59230, ZN => n2639);
   U2079 : OAI22_X1 port map( A1 => n52450, A2 => n59310, B1 => n53448, B2 => 
                           n59301, ZN => n59231);
   U2080 : INV_X1 port map( A => n59231, ZN => n2664);
   U2081 : OAI22_X1 port map( A1 => n52448, A2 => n59308, B1 => n53500, B2 => 
                           n59286, ZN => n59232);
   U2082 : INV_X1 port map( A => n59232, ZN => n2543);
   U2083 : OAI22_X1 port map( A1 => n52450, A2 => n59308, B1 => n53499, B2 => 
                           n59301, ZN => n59233);
   U2084 : INV_X1 port map( A => n59233, ZN => n2542);
   U2085 : OAI22_X1 port map( A1 => n52435, A2 => n59308, B1 => n53359, B2 => 
                           n59244, ZN => n59234);
   U2086 : INV_X1 port map( A => n59234, ZN => n2559);
   U2087 : OAI22_X1 port map( A1 => n52448, A2 => n59293, B1 => n53498, B2 => 
                           n59286, ZN => n59235);
   U2088 : INV_X1 port map( A => n59235, ZN => n2575);
   U2089 : OAI22_X1 port map( A1 => n52442, A2 => n59267, B1 => n53497, B2 => 
                           n59321, ZN => n59236);
   U2090 : INV_X1 port map( A => n59236, ZN => n2638);
   U2091 : OAI22_X1 port map( A1 => n52442, A2 => n59255, B1 => n53496, B2 => 
                           n59321, ZN => n59237);
   U2092 : INV_X1 port map( A => n59237, ZN => n2734);
   U2093 : OAI22_X1 port map( A1 => n52450, A2 => n59328, B1 => n53495, B2 => 
                           n59301, ZN => n59238);
   U2094 : INV_X1 port map( A => n59238, ZN => n2733);
   U2095 : OAI22_X1 port map( A1 => n52448, A2 => n59328, B1 => n53494, B2 => 
                           n59286, ZN => n59239);
   U2096 : INV_X1 port map( A => n59239, ZN => n2732);
   U2097 : OAI22_X1 port map( A1 => n52448, A2 => n59279, B1 => n53493, B2 => 
                           n59286, ZN => n59240);
   U2098 : INV_X1 port map( A => n59240, ZN => n2670);
   U2099 : OAI22_X1 port map( A1 => n52457, A2 => n59255, B1 => n53234, B2 => 
                           n59318, ZN => n59241);
   U2100 : INV_X1 port map( A => n59241, ZN => n2743);
   U2101 : OAI22_X1 port map( A1 => n52457, A2 => n59279, B1 => n53235, B2 => 
                           n59318, ZN => n59242);
   U2102 : INV_X1 port map( A => n59242, ZN => n2679);
   U2103 : OAI22_X1 port map( A1 => n52443, A2 => n59293, B1 => n53348, B2 => 
                           n59299, ZN => n59243);
   U2104 : INV_X1 port map( A => n59243, ZN => n2589);
   U2105 : OAI22_X1 port map( A1 => n52435, A2 => n59319, B1 => n53384, B2 => 
                           n59244, ZN => n59245);
   U2106 : INV_X1 port map( A => n59245, ZN => n2625);
   U2107 : OAI22_X1 port map( A1 => n52457, A2 => n59267, B1 => n53236, B2 => 
                           n59318, ZN => n59246);
   U2108 : INV_X1 port map( A => n59246, ZN => n2648);
   U2109 : OAI22_X1 port map( A1 => n52442, A2 => n59264, B1 => n53488, B2 => 
                           n59321, ZN => n59247);
   U2110 : INV_X1 port map( A => n59247, ZN => n2573);
   U2111 : OAI22_X1 port map( A1 => n52467, A2 => n59287, B1 => n53487, B2 => 
                           n59316, ZN => n59248);
   U2112 : INV_X1 port map( A => n59248, ZN => n2694);
   U2113 : OAI22_X1 port map( A1 => n52457, A2 => n59293, B1 => n53237, B2 => 
                           n59318, ZN => n59249);
   U2114 : INV_X1 port map( A => n59249, ZN => n2581);
   U2115 : OAI22_X1 port map( A1 => n52443, A2 => n59255, B1 => n53301, B2 => 
                           n59299, ZN => n59250);
   U2116 : INV_X1 port map( A => n59250, ZN => n2750);
   U2117 : OAI22_X1 port map( A1 => n52438, A2 => n59293, B1 => n53246, B2 => 
                           n59307, ZN => n59251);
   U2118 : INV_X1 port map( A => n59251, ZN => n2583);
   U2119 : OAI22_X1 port map( A1 => n52447, A2 => n59267, B1 => n53320, B2 => 
                           n59314, ZN => n59252);
   U2120 : INV_X1 port map( A => n59252, ZN => n2653);
   U2121 : OAI22_X1 port map( A1 => n52443, A2 => n59319, B1 => n53352, B2 => 
                           n59299, ZN => n59253);
   U2122 : INV_X1 port map( A => n59253, ZN => n2621);
   U2123 : OAI22_X1 port map( A1 => n52441, A2 => n59295, B1 => n53492, B2 => 
                           n59327, ZN => n59254);
   U2124 : INV_X1 port map( A => n59254, ZN => n2765);
   U2125 : OAI22_X1 port map( A1 => n52438, A2 => n59255, B1 => n53252, B2 => 
                           n59307, ZN => n59256);
   U2126 : INV_X1 port map( A => n59256, ZN => n2745);
   U2127 : OAI22_X1 port map( A1 => n52447, A2 => n59293, B1 => n53351, B2 => 
                           n59314, ZN => n59257);
   U2128 : INV_X1 port map( A => n59257, ZN => n2590);
   U2129 : OAI22_X1 port map( A1 => n52467, A2 => n59302, B1 => n53491, B2 => 
                           n59316, ZN => n59258);
   U2130 : INV_X1 port map( A => n59258, ZN => n2637);
   U2131 : OAI22_X1 port map( A1 => n52447, A2 => n59308, B1 => n53314, B2 => 
                           n59314, ZN => n59259);
   U2132 : INV_X1 port map( A => n59259, ZN => n2556);
   U2133 : OAI22_X1 port map( A1 => n52440, A2 => n59312, B1 => n53312, B2 => 
                           n59284, ZN => n59260);
   U2134 : INV_X1 port map( A => n59260, ZN => n2779);
   U2135 : OAI22_X1 port map( A1 => n52457, A2 => n59308, B1 => n53274, B2 => 
                           n59318, ZN => n59261);
   U2136 : INV_X1 port map( A => n59261, ZN => n2549);
   U2137 : OAI22_X1 port map( A1 => n52463, A2 => n59312, B1 => n53316, B2 => 
                           n59324, ZN => n59262);
   U2138 : INV_X1 port map( A => n59262, ZN => n2780);
   U2139 : OAI22_X1 port map( A1 => n52443, A2 => n59312, B1 => n53275, B2 => 
                           n59299, ZN => n59263);
   U2140 : INV_X1 port map( A => n59263, ZN => n2776);
   U2141 : OAI22_X1 port map( A1 => n52441, A2 => n59264, B1 => n53450, B2 => 
                           n59327, ZN => n59265);
   U2142 : INV_X1 port map( A => n59265, ZN => n2568);
   U2143 : OAI22_X1 port map( A1 => n52447, A2 => n59319, B1 => n53347, B2 => 
                           n59314, ZN => n59266);
   U2144 : INV_X1 port map( A => n59266, ZN => n2620);
   U2145 : OAI22_X1 port map( A1 => n52438, A2 => n59267, B1 => n53242, B2 => 
                           n59307, ZN => n59268);
   U2146 : INV_X1 port map( A => n59268, ZN => n2649);
   U2147 : OAI22_X1 port map( A1 => n52439, A2 => n59308, B1 => n53243, B2 => 
                           n59269, ZN => n59270);
   U2148 : INV_X1 port map( A => n59270, ZN => n2546);
   U2149 : OAI22_X1 port map( A1 => n52443, A2 => n59279, B1 => n53345, B2 => 
                           n59299, ZN => n59271);
   U2150 : INV_X1 port map( A => n59271, ZN => n2686);
   U2151 : OAI22_X1 port map( A1 => n52450, A2 => n59287, B1 => n53482, B2 => 
                           n59301, ZN => n59272);
   U2152 : INV_X1 port map( A => n59272, ZN => n2695);
   U2153 : OAI22_X1 port map( A1 => n52437, A2 => n59279, B1 => n53341, B2 => 
                           n59297, ZN => n59273);
   U2154 : INV_X1 port map( A => n59273, ZN => n2684);
   U2155 : OAI22_X1 port map( A1 => n52453, A2 => n59312, B1 => n53250, B2 => 
                           n59305, ZN => n59274);
   U2156 : INV_X1 port map( A => n59274, ZN => n2772);
   U2157 : OAI22_X1 port map( A1 => n52437, A2 => n59325, B1 => n53339, B2 => 
                           n59297, ZN => n59275);
   U2158 : INV_X1 port map( A => n59275, ZN => n2718);
   U2159 : OAI22_X1 port map( A1 => n52467, A2 => n59319, B1 => n53478, B2 => 
                           n59316, ZN => n59276);
   U2160 : INV_X1 port map( A => n59276, ZN => n2606);
   U2161 : OAI22_X1 port map( A1 => n52453, A2 => n59277, B1 => n53336, B2 => 
                           n59305, ZN => n59278);
   U2162 : INV_X1 port map( A => n59278, ZN => n2618);
   U2163 : OAI22_X1 port map( A1 => n52447, A2 => n59279, B1 => n53334, B2 => 
                           n59314, ZN => n59280);
   U2164 : INV_X1 port map( A => n59280, ZN => n2683);
   U2165 : OAI22_X1 port map( A1 => n52440, A2 => n59293, B1 => n53332, B2 => 
                           n59284, ZN => n59281);
   U2166 : INV_X1 port map( A => n59281, ZN => n2587);
   U2167 : OAI22_X1 port map( A1 => n52463, A2 => n59293, B1 => n53330, B2 => 
                           n59324, ZN => n59282);
   U2168 : INV_X1 port map( A => n59282, ZN => n2586);
   U2169 : OAI22_X1 port map( A1 => n52457, A2 => n59287, B1 => n53258, B2 => 
                           n59318, ZN => n59283);
   U2170 : INV_X1 port map( A => n59283, ZN => n2707);
   U2171 : OAI22_X1 port map( A1 => n52440, A2 => n59308, B1 => n53290, B2 => 
                           n59284, ZN => n59285);
   U2172 : INV_X1 port map( A => n59285, ZN => n2551);
   U2173 : OAI22_X1 port map( A1 => n52448, A2 => n59287, B1 => n53471, B2 => 
                           n59286, ZN => n59288);
   U2174 : INV_X1 port map( A => n59288, ZN => n2696);
   U2175 : OAI22_X1 port map( A1 => n52443, A2 => n59325, B1 => n53328, B2 => 
                           n59299, ZN => n59289);
   U2176 : INV_X1 port map( A => n59289, ZN => n2717);
   U2177 : OAI22_X1 port map( A1 => n52450, A2 => n59293, B1 => n53449, B2 => 
                           n59301, ZN => n59290);
   U2178 : INV_X1 port map( A => n59290, ZN => n2597);
   U2179 : OAI22_X1 port map( A1 => n52450, A2 => n59295, B1 => n53474, B2 => 
                           n59301, ZN => n59291);
   U2180 : INV_X1 port map( A => n59291, ZN => n2761);
   U2181 : OAI22_X1 port map( A1 => n52437, A2 => n59312, B1 => n53327, B2 => 
                           n59297, ZN => n59292);
   U2182 : INV_X1 port map( A => n59292, ZN => n2781);
   U2183 : OAI22_X1 port map( A1 => n52467, A2 => n59293, B1 => n53489, B2 => 
                           n59316, ZN => n59294);
   U2184 : INV_X1 port map( A => n59294, ZN => n2574);
   U2185 : OAI22_X1 port map( A1 => n52457, A2 => n59295, B1 => n53286, B2 => 
                           n59318, ZN => n59296);
   U2186 : INV_X1 port map( A => n59296, ZN => n2778);
   U2187 : OAI22_X1 port map( A1 => n52437, A2 => n59319, B1 => n53302, B2 => 
                           n59297, ZN => n59298);
   U2188 : INV_X1 port map( A => n59298, ZN => n2616);
   U2189 : OAI22_X1 port map( A1 => n52443, A2 => n59308, B1 => n53322, B2 => 
                           n59299, ZN => n59300);
   U2190 : INV_X1 port map( A => n59300, ZN => n2558);
   U2191 : OAI22_X1 port map( A1 => n52450, A2 => n59302, B1 => n53452, B2 => 
                           n59301, ZN => n59303);
   U2192 : INV_X1 port map( A => n59303, ZN => n2634);
   U2193 : OAI22_X1 port map( A1 => n52442, A2 => n59310, B1 => n53485, B2 => 
                           n59321, ZN => n59304);
   U2194 : INV_X1 port map( A => n59304, ZN => n2669);
   U2195 : OAI22_X1 port map( A1 => n52453, A2 => n59308, B1 => n53300, B2 => 
                           n59305, ZN => n59306);
   U2196 : INV_X1 port map( A => n59306, ZN => n2552);
   U2197 : OAI22_X1 port map( A1 => n52438, A2 => n59308, B1 => n53266, B2 => 
                           n59307, ZN => n59309);
   U2198 : INV_X1 port map( A => n59309, ZN => n2548);
   U2199 : OAI22_X1 port map( A1 => n52441, A2 => n59310, B1 => n53454, B2 => 
                           n59327, ZN => n59311);
   U2200 : INV_X1 port map( A => n59311, ZN => n2666);
   U2201 : OAI22_X1 port map( A1 => n52447, A2 => n59312, B1 => n53277, B2 => 
                           n59314, ZN => n59313);
   U2202 : INV_X1 port map( A => n59313, ZN => n2777);
   U2203 : OAI22_X1 port map( A1 => n52447, A2 => n59325, B1 => n53319, B2 => 
                           n59314, ZN => n59315);
   U2204 : INV_X1 port map( A => n59315, ZN => n2714);
   U2205 : OAI22_X1 port map( A1 => n52467, A2 => n59322, B1 => n53465, B2 => 
                           n59316, ZN => n59317);
   U2206 : INV_X1 port map( A => n59317, ZN => n2536);
   U2207 : OAI22_X1 port map( A1 => n52457, A2 => n59319, B1 => n53276, B2 => 
                           n59318, ZN => n59320);
   U2208 : INV_X1 port map( A => n59320, ZN => n2612);
   U2209 : OAI22_X1 port map( A1 => n52442, A2 => n59322, B1 => n53480, B2 => 
                           n59321, ZN => n59323);
   U2210 : INV_X1 port map( A => n59323, ZN => n2539);
   U2211 : OAI22_X1 port map( A1 => n52463, A2 => n59325, B1 => n53281, B2 => 
                           n59324, ZN => n59326);
   U2212 : INV_X1 port map( A => n59326, ZN => n2711);
   U2213 : OAI22_X1 port map( A1 => n52441, A2 => n59328, B1 => n53477, B2 => 
                           n59327, ZN => n59329);
   U2214 : INV_X1 port map( A => n59329, ZN => n2730);
   U2215 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1),
                           ZN => n40561);
   U2216 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n53531, ZN => 
                           n59336);
   U2217 : NOR2_X1 port map( A1 => n53511, A2 => n59336, ZN => n59334);
   U2218 : NAND2_X1 port map( A1 => n52397, A2 => n59334, ZN => n40647);
   U2219 : INV_X1 port map( A => ADD_WR(0), ZN => n59330);
   U2220 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n59330, ZN
                           => n40558);
   U2221 : NAND2_X1 port map( A1 => n59334, A2 => n52394, ZN => n40646);
   U2222 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n59330, ZN => n59331);
   U2223 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n59331, ZN => n40643);
   U2224 : NAND2_X1 port map( A1 => n59334, A2 => n52474, ZN => n40642);
   U2225 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n59332);
   U2226 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n59332, ZN => n40639);
   U2227 : NAND2_X1 port map( A1 => n59334, A2 => n52470, ZN => n40638);
   U2228 : INV_X1 port map( A => ADD_WR(2), ZN => n59333);
   U2229 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n59333, ZN
                           => n40555);
   U2230 : NAND2_X1 port map( A1 => n59334, A2 => n52391, ZN => n40637);
   U2231 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n59330, A3 => n59333, ZN =>
                           n40552);
   U2232 : NAND2_X1 port map( A1 => n59334, A2 => n52388, ZN => n40636);
   U2233 : NOR2_X1 port map( A1 => n59333, A2 => n59331, ZN => n40633);
   U2234 : NAND2_X1 port map( A1 => n59334, A2 => n52464, ZN => n40632);
   U2235 : NOR2_X1 port map( A1 => n59333, A2 => n59332, ZN => n40629);
   U2236 : NAND2_X1 port map( A1 => n59334, A2 => n52460, ZN => n40628);
   U2237 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n53530, ZN => 
                           n59338);
   U2238 : NOR2_X1 port map( A1 => n53511, A2 => n59338, ZN => n59335);
   U2239 : NAND2_X1 port map( A1 => n52397, A2 => n59335, ZN => n40627);
   U2240 : NAND2_X1 port map( A1 => n52394, A2 => n59335, ZN => n40626);
   U2241 : NAND2_X1 port map( A1 => n52474, A2 => n59335, ZN => n40625);
   U2242 : NAND2_X1 port map( A1 => n52470, A2 => n59335, ZN => n40624);
   U2243 : NAND2_X1 port map( A1 => n52391, A2 => n59335, ZN => n40623);
   U2244 : NAND2_X1 port map( A1 => n52388, A2 => n59335, ZN => n40622);
   U2245 : NAND2_X1 port map( A1 => n52464, A2 => n59335, ZN => n40621);
   U2246 : NAND2_X1 port map( A1 => n52460, A2 => n59335, ZN => n40620);
   U2247 : NOR2_X1 port map( A1 => n53509, A2 => n59336, ZN => n59337);
   U2248 : NAND2_X1 port map( A1 => n52397, A2 => n59337, ZN => n40619);
   U2249 : NAND2_X1 port map( A1 => n52394, A2 => n59337, ZN => n40618);
   U2250 : NAND2_X1 port map( A1 => n52474, A2 => n59337, ZN => n40617);
   U2251 : NAND2_X1 port map( A1 => n52470, A2 => n59337, ZN => n40616);
   U2252 : NAND2_X1 port map( A1 => n52391, A2 => n59337, ZN => n40615);
   U2253 : NAND2_X1 port map( A1 => n52388, A2 => n59337, ZN => n40614);
   U2254 : NAND2_X1 port map( A1 => n52464, A2 => n59337, ZN => n40613);
   U2255 : NAND2_X1 port map( A1 => n52460, A2 => n59337, ZN => n40612);
   U2256 : NOR2_X1 port map( A1 => n53509, A2 => n59338, ZN => n59339);
   U2257 : NAND2_X1 port map( A1 => n52397, A2 => n59339, ZN => n40611);
   U2258 : NAND2_X1 port map( A1 => n52394, A2 => n59339, ZN => n40610);
   U2259 : NAND2_X1 port map( A1 => n52474, A2 => n59339, ZN => n40609);
   U2260 : NAND2_X1 port map( A1 => n52470, A2 => n59339, ZN => n40608);
   U2261 : NAND2_X1 port map( A1 => n52391, A2 => n59339, ZN => n40607);
   U2262 : NAND2_X1 port map( A1 => n52388, A2 => n59339, ZN => n40606);
   U2263 : NAND2_X1 port map( A1 => n52464, A2 => n59339, ZN => n40605);
   U2264 : NAND2_X1 port map( A1 => n52460, A2 => n59339, ZN => n40604);
   U2265 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n3567, ZN => n59348);
   U2266 : INV_X1 port map( A => n3573, ZN => n59341);
   U2267 : NOR2_X1 port map( A1 => n59348, A2 => n59341, ZN => n47429);
   U2268 : INV_X1 port map( A => n3571, ZN => n59346);
   U2269 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n59343)
                           ;
   U2270 : NOR2_X1 port map( A1 => n59346, A2 => n59343, ZN => n49092);
   U2271 : NOR2_X1 port map( A1 => n59343, A2 => n3572, ZN => n49093);
   U2272 : INV_X1 port map( A => n3574, ZN => n59340);
   U2273 : NOR2_X1 port map( A1 => n59343, A2 => n59340, ZN => n49094);
   U2274 : NOR2_X1 port map( A1 => n59348, A2 => n3572, ZN => n49087);
   U2275 : INV_X1 port map( A => n3570, ZN => n59345);
   U2276 : NOR2_X1 port map( A1 => n59343, A2 => n59345, ZN => n49089);
   U2277 : INV_X1 port map( A => n3569, ZN => n59347);
   U2278 : NOR2_X1 port map( A1 => n59343, A2 => n59347, ZN => n49091);
   U2279 : NOR2_X1 port map( A1 => n59348, A2 => n59340, ZN => n49090);
   U2280 : INV_X1 port map( A => n3568, ZN => n59342);
   U2281 : NOR2_X1 port map( A1 => n59348, A2 => n59342, ZN => n49086);
   U2282 : NOR2_X1 port map( A1 => n59341, A2 => n59343, ZN => n49088);
   U2283 : NOR2_X1 port map( A1 => n59343, A2 => n59342, ZN => n47428);
   U2284 : INV_X1 port map( A => n3575, ZN => n59344);
   U2285 : NOR2_X1 port map( A1 => n59343, A2 => n59344, ZN => n40592);
   U2286 : NOR2_X1 port map( A1 => n59348, A2 => n59344, ZN => n40591);
   U2287 : NOR2_X1 port map( A1 => n59348, A2 => n59345, ZN => n49085);
   U2288 : NOR2_X1 port map( A1 => n59348, A2 => n59346, ZN => n40589);
   U2289 : NOR2_X1 port map( A1 => n59348, A2 => n59347, ZN => n40588);
   U2290 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n53629, A3 => n53626, ZN 
                           => n60059);
   U2291 : AOI22_X1 port map( A1 => n51548, A2 => n53585, B1 => n51556, B2 => 
                           n52421, ZN => n59352);
   U2292 : AOI22_X1 port map( A1 => n51604, A2 => n52425, B1 => n51409, B2 => 
                           n52428, ZN => n59351);
   U2293 : AOI22_X1 port map( A1 => n51557, A2 => n53588, B1 => n51371, B2 => 
                           n52426, ZN => n59350);
   U2294 : AOI22_X1 port map( A1 => n51370, A2 => n52430, B1 => n51390, B2 => 
                           n52424, ZN => n59349);
   U2295 : NAND4_X1 port map( A1 => n59352, A2 => n59351, A3 => n59350, A4 => 
                           n59349, ZN => n59358);
   U2296 : AOI22_X1 port map( A1 => n51645, A2 => n52423, B1 => n51580, B2 => 
                           n52432, ZN => n59356);
   U2297 : AOI22_X1 port map( A1 => n51555, A2 => n53586, B1 => n51387, B2 => 
                           n52422, ZN => n59355);
   U2298 : AOI22_X1 port map( A1 => n51389, A2 => n53589, B1 => n51511, B2 => 
                           n52431, ZN => n59354);
   U2299 : AOI22_X1 port map( A1 => n51493, A2 => n53587, B1 => n51627, B2 => 
                           n52429, ZN => n59353);
   U2300 : NAND4_X1 port map( A1 => n59356, A2 => n59355, A3 => n59354, A4 => 
                           n59353, ZN => n59357);
   U2301 : NOR2_X1 port map( A1 => n59358, A2 => n59357, ZN => n59370);
   U2302 : NOR3_X1 port map( A1 => n53622, A2 => n53623, A3 => n59857, ZN => 
                           n59810);
   U2303 : CLKBUF_X1 port map( A => n59810, Z => n59878);
   U2304 : AOI22_X1 port map( A1 => n51465, A2 => n53580, B1 => n51405, B2 => 
                           n53514, ZN => n59362);
   U2305 : AOI22_X1 port map( A1 => n51470, A2 => n53581, B1 => n51452, B2 => 
                           n53519, ZN => n59361);
   U2306 : AOI22_X1 port map( A1 => n51478, A2 => n53584, B1 => n51668, B2 => 
                           n53582, ZN => n59360);
   U2307 : AOI22_X1 port map( A1 => n51464, A2 => n53583, B1 => n51455, B2 => 
                           n53513, ZN => n59359);
   U2308 : NAND4_X1 port map( A1 => n59362, A2 => n59361, A3 => n59360, A4 => 
                           n59359, ZN => n59368);
   U2309 : NOR3_X1 port map( A1 => n53623, A2 => n52484, A3 => n59857, ZN => 
                           n59588);
   U2310 : CLKBUF_X1 port map( A => n59588, Z => n60054);
   U2311 : AOI22_X1 port map( A1 => n51565, A2 => n53577, B1 => n51566, B2 => 
                           n53515, ZN => n59366);
   U2312 : AOI22_X1 port map( A1 => n53519, A2 => n51394, B1 => n51596, B2 => 
                           n53579, ZN => n59365);
   U2313 : AOI22_X1 port map( A1 => n53582, A2 => n51395, B1 => n51617, B2 => 
                           n52400, ZN => n59364);
   U2314 : AOI22_X1 port map( A1 => n51570, A2 => n53578, B1 => n51583, B2 => 
                           n53516, ZN => n59363);
   U2315 : NAND4_X1 port map( A1 => n59366, A2 => n59365, A3 => n59364, A4 => 
                           n59363, ZN => n59367);
   U2316 : AOI22_X1 port map( A1 => n59878, A2 => n59368, B1 => n60054, B2 => 
                           n59367, ZN => n59369);
   U2317 : OAI21_X1 port map( B1 => n59857, B2 => n59370, A => n59369, ZN => 
                           OUT2(31));
   U2318 : AOI22_X1 port map( A1 => n52428, A2 => n51420, B1 => n51382, B2 => 
                           n53575, ZN => n59374);
   U2319 : AOI22_X1 port map( A1 => n52422, A2 => n51414, B1 => n52432, B2 => 
                           n51538, ZN => n59373);
   U2320 : AOI22_X1 port map( A1 => n53587, A2 => n51462, B1 => n51624, B2 => 
                           n53576, ZN => n59372);
   U2321 : AOI22_X1 port map( A1 => n53589, A2 => n51413, B1 => n52421, B2 => 
                           n51519, ZN => n59371);
   U2322 : NAND4_X1 port map( A1 => n59374, A2 => n59373, A3 => n59372, A4 => 
                           n59371, ZN => n59380);
   U2323 : AOI22_X1 port map( A1 => n52430, A2 => n51372, B1 => n51644, B2 => 
                           n53573, ZN => n59378);
   U2324 : AOI22_X1 port map( A1 => n52423, A2 => n51650, B1 => n51421, B2 => 
                           n53572, ZN => n59377);
   U2325 : AOI22_X1 port map( A1 => n53588, A2 => n51535, B1 => n51522, B2 => 
                           n52427, ZN => n59376);
   U2326 : AOI22_X1 port map( A1 => n51446, A2 => n53574, B1 => n51680, B2 => 
                           n52434, ZN => n59375);
   U2327 : NAND4_X1 port map( A1 => n59378, A2 => n59377, A3 => n59376, A4 => 
                           n59375, ZN => n59379);
   U2328 : NOR2_X1 port map( A1 => n59380, A2 => n59379, ZN => n59392);
   U2329 : AOI22_X1 port map( A1 => n53577, A2 => n51496, B1 => n52400, B2 => 
                           n51463, ZN => n59384);
   U2330 : AOI22_X1 port map( A1 => n51461, A2 => n53512, B1 => n51540, B2 => 
                           n53520, ZN => n59383);
   U2331 : AOI22_X1 port map( A1 => n53519, A2 => n51441, B1 => n53516, B2 => 
                           n51436, ZN => n59382);
   U2332 : AOI22_X1 port map( A1 => n53515, A2 => n51444, B1 => n51381, B2 => 
                           n53571, ZN => n59381);
   U2333 : NAND4_X1 port map( A1 => n59384, A2 => n59383, A3 => n59382, A4 => 
                           n59381, ZN => n59390);
   U2334 : AOI22_X1 port map( A1 => n53519, A2 => n51411, B1 => n51407, B2 => 
                           n53570, ZN => n59388);
   U2335 : AOI22_X1 port map( A1 => n53516, A2 => n51629, B1 => n53571, B2 => 
                           n51677, ZN => n59387);
   U2336 : AOI22_X1 port map( A1 => n53513, A2 => n51564, B1 => n51639, B2 => 
                           n53523, ZN => n59386);
   U2337 : AOI22_X1 port map( A1 => n53515, A2 => n51614, B1 => n53579, B2 => 
                           n51633, ZN => n59385);
   U2338 : NAND4_X1 port map( A1 => n59388, A2 => n59387, A3 => n59386, A4 => 
                           n59385, ZN => n59389);
   U2339 : AOI22_X1 port map( A1 => n59878, A2 => n59390, B1 => n60054, B2 => 
                           n59389, ZN => n59391);
   U2340 : OAI21_X1 port map( B1 => n59857, B2 => n59392, A => n59391, ZN => 
                           OUT2(30));
   U2341 : AOI22_X1 port map( A1 => n53573, A2 => n51657, B1 => n52427, B2 => 
                           n51518, ZN => n59396);
   U2342 : AOI22_X1 port map( A1 => n52422, A2 => n51431, B1 => n52425, B2 => 
                           n51658, ZN => n59395);
   U2343 : AOI22_X1 port map( A1 => n52432, A2 => n51648, B1 => n52426, B2 => 
                           n51432, ZN => n59394);
   U2344 : AOI22_X1 port map( A1 => n53586, A2 => n51517, B1 => n53587, B2 => 
                           n51472, ZN => n59393);
   U2345 : NAND4_X1 port map( A1 => n59396, A2 => n59395, A3 => n59394, A4 => 
                           n59393, ZN => n59402);
   U2346 : AOI22_X1 port map( A1 => n53589, A2 => n51424, B1 => n51433, B2 => 
                           n53569, ZN => n59400);
   U2347 : AOI22_X1 port map( A1 => n52430, A2 => n51366, B1 => n52424, B2 => 
                           n51434, ZN => n59399);
   U2348 : AOI22_X1 port map( A1 => n52431, A2 => n51486, B1 => n51568, B2 => 
                           n53568, ZN => n59398);
   U2349 : AOI22_X1 port map( A1 => n51524, A2 => n52419, B1 => n51523, B2 => 
                           n53567, ZN => n59397);
   U2350 : NAND4_X1 port map( A1 => n59400, A2 => n59399, A3 => n59398, A4 => 
                           n59397, ZN => n59401);
   U2351 : NOR2_X1 port map( A1 => n59402, A2 => n59401, ZN => n59414);
   U2352 : AOI22_X1 port map( A1 => n53519, A2 => n51492, B1 => n53520, B2 => 
                           n51577, ZN => n59406);
   U2353 : AOI22_X1 port map( A1 => n53577, A2 => n51497, B1 => n51490, B2 => 
                           n53566, ZN => n59405);
   U2354 : AOI22_X1 port map( A1 => n52400, A2 => n51489, B1 => n53571, B2 => 
                           n51392, ZN => n59404);
   U2355 : AOI22_X1 port map( A1 => n53579, A2 => n51459, B1 => n53516, B2 => 
                           n51460, ZN => n59403);
   U2356 : NAND4_X1 port map( A1 => n59406, A2 => n59405, A3 => n59404, A4 => 
                           n59403, ZN => n59412);
   U2357 : AOI22_X1 port map( A1 => n53584, A2 => n51587, B1 => n53577, B2 => 
                           n51563, ZN => n59410);
   U2358 : AOI22_X1 port map( A1 => n53570, A2 => n51406, B1 => n53523, B2 => 
                           n51588, ZN => n59409);
   U2359 : AOI22_X1 port map( A1 => n53512, A2 => n51594, B1 => n53571, B2 => 
                           n51534, ZN => n59408);
   U2360 : AOI22_X1 port map( A1 => n53581, A2 => n51606, B1 => n53519, B2 => 
                           n51400, ZN => n59407);
   U2361 : NAND4_X1 port map( A1 => n59410, A2 => n59409, A3 => n59408, A4 => 
                           n59407, ZN => n59411);
   U2362 : AOI22_X1 port map( A1 => n59878, A2 => n59412, B1 => n60054, B2 => 
                           n59411, ZN => n59413);
   U2363 : OAI21_X1 port map( B1 => n59857, B2 => n59414, A => n59413, ZN => 
                           OUT2(29));
   U2364 : AOI22_X1 port map( A1 => n53576, A2 => n51628, B1 => n53569, B2 => 
                           n51426, ZN => n59418);
   U2365 : AOI22_X1 port map( A1 => n52430, A2 => n51368, B1 => n51415, B2 => 
                           n52420, ZN => n59417);
   U2366 : AOI22_X1 port map( A1 => n52424, A2 => n51373, B1 => n52427, B2 => 
                           n51571, ZN => n59416);
   U2367 : AOI22_X1 port map( A1 => n53586, A2 => n51675, B1 => n53573, B2 => 
                           n51643, ZN => n59415);
   U2368 : NAND4_X1 port map( A1 => n59418, A2 => n59417, A3 => n59416, A4 => 
                           n59415, ZN => n59424);
   U2369 : AOI22_X1 port map( A1 => n52422, A2 => n51419, B1 => n53567, B2 => 
                           n51550, ZN => n59422);
   U2370 : AOI22_X1 port map( A1 => n52432, A2 => n51672, B1 => n53572, B2 => 
                           n51418, ZN => n59421);
   U2371 : AOI22_X1 port map( A1 => n53587, A2 => n51448, B1 => n53568, B2 => 
                           n51651, ZN => n59420);
   U2372 : AOI22_X1 port map( A1 => n52431, A2 => n51454, B1 => n52419, B2 => 
                           n51549, ZN => n59419);
   U2373 : NAND4_X1 port map( A1 => n59422, A2 => n59421, A3 => n59420, A4 => 
                           n59419, ZN => n59423);
   U2374 : NOR2_X1 port map( A1 => n59424, A2 => n59423, ZN => n59436);
   U2375 : AOI22_X1 port map( A1 => n53519, A2 => n51503, B1 => n53523, B2 => 
                           n51505, ZN => n59428);
   U2376 : AOI22_X1 port map( A1 => n53584, A2 => n51442, B1 => n53512, B2 => 
                           n51450, ZN => n59427);
   U2377 : AOI22_X1 port map( A1 => n53514, A2 => n51379, B1 => n53577, B2 => 
                           n51447, ZN => n59426);
   U2378 : AOI22_X1 port map( A1 => n53515, A2 => n51506, B1 => n53570, B2 => 
                           n51671, ZN => n59425);
   U2379 : NAND4_X1 port map( A1 => n59428, A2 => n59427, A3 => n59426, A4 => 
                           n59425, ZN => n59434);
   U2380 : AOI22_X1 port map( A1 => n53515, A2 => n51597, B1 => n52400, B2 => 
                           n51640, ZN => n59432);
   U2381 : AOI22_X1 port map( A1 => n53512, A2 => n51634, B1 => n51647, B2 => 
                           n53565, ZN => n59431);
   U2382 : AOI22_X1 port map( A1 => n53519, A2 => n51428, B1 => n53571, B2 => 
                           n51673, ZN => n59430);
   U2383 : AOI22_X1 port map( A1 => n53577, A2 => n51561, B1 => n53570, B2 => 
                           n51404, ZN => n59429);
   U2384 : NAND4_X1 port map( A1 => n59432, A2 => n59431, A3 => n59430, A4 => 
                           n59429, ZN => n59433);
   U2385 : AOI22_X1 port map( A1 => n59878, A2 => n59434, B1 => n60054, B2 => 
                           n59433, ZN => n59435);
   U2386 : OAI21_X1 port map( B1 => n59857, B2 => n59436, A => n59435, ZN => 
                           OUT2(28));
   U2387 : AOI22_X1 port map( A1 => n52427, A2 => n51525, B1 => n51377, B2 => 
                           n53563, ZN => n59440);
   U2388 : AOI22_X1 port map( A1 => n52432, A2 => n51676, B1 => n53569, B2 => 
                           n51416, ZN => n59439);
   U2389 : AOI22_X1 port map( A1 => n52423, A2 => n51529, B1 => n52434, B2 => 
                           n51679, ZN => n59438);
   U2390 : AOI22_X1 port map( A1 => n52420, A2 => n51410, B1 => n51423, B2 => 
                           n53564, ZN => n59437);
   U2391 : NAND4_X1 port map( A1 => n59440, A2 => n59439, A3 => n59438, A4 => 
                           n59437, ZN => n59446);
   U2392 : AOI22_X1 port map( A1 => n53587, A2 => n51453, B1 => n53572, B2 => 
                           n51422, ZN => n59444);
   U2393 : AOI22_X1 port map( A1 => n53588, A2 => n51528, B1 => n53573, B2 => 
                           n51642, ZN => n59443);
   U2394 : AOI22_X1 port map( A1 => n52431, A2 => n51438, B1 => n53575, B2 => 
                           n51385, ZN => n59442);
   U2395 : AOI22_X1 port map( A1 => n52425, A2 => n51653, B1 => n53567, B2 => 
                           n51536, ZN => n59441);
   U2396 : NAND4_X1 port map( A1 => n59444, A2 => n59443, A3 => n59442, A4 => 
                           n59441, ZN => n59445);
   U2397 : NOR2_X1 port map( A1 => n59446, A2 => n59445, ZN => n59458);
   U2398 : AOI22_X1 port map( A1 => n53513, A2 => n51494, B1 => n53565, B2 => 
                           n51451, ZN => n59450);
   U2399 : AOI22_X1 port map( A1 => n53514, A2 => n51365, B1 => n53519, B2 => 
                           n51479, ZN => n59449);
   U2400 : AOI22_X1 port map( A1 => n53515, A2 => n51469, B1 => n53520, B2 => 
                           n51663, ZN => n59448);
   U2401 : AOI22_X1 port map( A1 => n52400, A2 => n51474, B1 => n53512, B2 => 
                           n51439, ZN => n59447);
   U2402 : NAND4_X1 port map( A1 => n59450, A2 => n59449, A3 => n59448, A4 => 
                           n59447, ZN => n59456);
   U2403 : AOI22_X1 port map( A1 => n53520, A2 => n51402, B1 => n51559, B2 => 
                           n53562, ZN => n59454);
   U2404 : AOI22_X1 port map( A1 => n53519, A2 => n51417, B1 => n53523, B2 => 
                           n51641, ZN => n59453);
   U2405 : AOI22_X1 port map( A1 => n53515, A2 => n51613, B1 => n53512, B2 => 
                           n51635, ZN => n59452);
   U2406 : AOI22_X1 port map( A1 => n53584, A2 => n51630, B1 => n53578, B2 => 
                           n51661, ZN => n59451);
   U2407 : NAND4_X1 port map( A1 => n59454, A2 => n59453, A3 => n59452, A4 => 
                           n59451, ZN => n59455);
   U2408 : AOI22_X1 port map( A1 => n59878, A2 => n59456, B1 => n59588, B2 => 
                           n59455, ZN => n59457);
   U2409 : OAI21_X1 port map( B1 => n59857, B2 => n59458, A => n59457, ZN => 
                           OUT2(27));
   U2410 : AOI22_X1 port map( A1 => n52423, A2 => n51531, B1 => n53569, B2 => 
                           n51430, ZN => n59462);
   U2411 : AOI22_X1 port map( A1 => n52424, A2 => n51429, B1 => n53576, B2 => 
                           n51655, ZN => n59461);
   U2412 : AOI22_X1 port map( A1 => n53587, A2 => n51491, B1 => n52430, B2 => 
                           n51399, ZN => n59460);
   U2413 : AOI22_X1 port map( A1 => n52431, A2 => n51485, B1 => n52434, B2 => 
                           n51547, ZN => n59459);
   U2414 : NAND4_X1 port map( A1 => n59462, A2 => n59461, A3 => n59460, A4 => 
                           n59459, ZN => n59468);
   U2415 : AOI22_X1 port map( A1 => n52422, A2 => n51425, B1 => n52427, B2 => 
                           n51542, ZN => n59466);
   U2416 : AOI22_X1 port map( A1 => n52420, A2 => n51427, B1 => n51649, B2 => 
                           n53561, ZN => n59465);
   U2417 : AOI22_X1 port map( A1 => n53573, A2 => n51660, B1 => n53567, B2 => 
                           n51551, ZN => n59464);
   U2418 : AOI22_X1 port map( A1 => n53588, A2 => n51567, B1 => n52426, B2 => 
                           n51388, ZN => n59463);
   U2419 : NAND4_X1 port map( A1 => n59466, A2 => n59465, A3 => n59464, A4 => 
                           n59463, ZN => n59467);
   U2420 : NOR2_X1 port map( A1 => n59468, A2 => n59467, ZN => n59480);
   U2421 : AOI22_X1 port map( A1 => n53584, A2 => n51458, B1 => n53515, B2 => 
                           n51466, ZN => n59472);
   U2422 : AOI22_X1 port map( A1 => n53512, A2 => n51475, B1 => n53520, B2 => 
                           n51589, ZN => n59471);
   U2423 : AOI22_X1 port map( A1 => n53523, A2 => n51467, B1 => n53562, B2 => 
                           n51488, ZN => n59470);
   U2424 : AOI22_X1 port map( A1 => n53514, A2 => n51383, B1 => n53519, B2 => 
                           n51457, ZN => n59469);
   U2425 : NAND4_X1 port map( A1 => n59472, A2 => n59471, A3 => n59470, A4 => 
                           n59469, ZN => n59478);
   U2426 : AOI22_X1 port map( A1 => n53519, A2 => n51403, B1 => n53512, B2 => 
                           n51612, ZN => n59476);
   U2427 : AOI22_X1 port map( A1 => n53584, A2 => n51591, B1 => n53562, B2 => 
                           n51546, ZN => n59475);
   U2428 : AOI22_X1 port map( A1 => n53581, A2 => n51598, B1 => n52400, B2 => 
                           n51610, ZN => n59474);
   U2429 : AOI22_X1 port map( A1 => n53514, A2 => n51572, B1 => n53582, B2 => 
                           n51401, ZN => n59473);
   U2430 : NAND4_X1 port map( A1 => n59476, A2 => n59475, A3 => n59474, A4 => 
                           n59473, ZN => n59477);
   U2431 : AOI22_X1 port map( A1 => n59878, A2 => n59478, B1 => n59588, B2 => 
                           n59477, ZN => n59479);
   U2432 : OAI21_X1 port map( B1 => n59857, B2 => n59480, A => n59479, ZN => 
                           OUT2(26));
   U2433 : AOI22_X1 port map( A1 => n52425, A2 => n51618, B1 => n53573, B2 => 
                           n51637, ZN => n59484);
   U2434 : AOI22_X1 port map( A1 => n52430, A2 => n51376, B1 => n52426, B2 => 
                           n51375, ZN => n59483);
   U2435 : AOI22_X1 port map( A1 => n53569, A2 => n51393, B1 => n52419, B2 => 
                           n51573, ZN => n59482);
   U2436 : AOI22_X1 port map( A1 => n53587, A2 => n51437, B1 => n53575, B2 => 
                           n51374, ZN => n59481);
   U2437 : NAND4_X1 port map( A1 => n59484, A2 => n59483, A3 => n59482, A4 => 
                           n59481, ZN => n59490);
   U2438 : AOI22_X1 port map( A1 => n53589, A2 => n51397, B1 => n53568, B2 => 
                           n51652, ZN => n59488);
   U2439 : AOI22_X1 port map( A1 => n52434, A2 => n51665, B1 => n53567, B2 => 
                           n51574, ZN => n59487);
   U2440 : AOI22_X1 port map( A1 => n52431, A2 => n51468, B1 => n53564, B2 => 
                           n51398, ZN => n59486);
   U2441 : AOI22_X1 port map( A1 => n52427, A2 => n51569, B1 => n53561, B2 => 
                           n51664, ZN => n59485);
   U2442 : NAND4_X1 port map( A1 => n59488, A2 => n59487, A3 => n59486, A4 => 
                           n59485, ZN => n59489);
   U2443 : NOR2_X1 port map( A1 => n59490, A2 => n59489, ZN => n59502);
   U2444 : AOI22_X1 port map( A1 => n53512, A2 => n51440, B1 => n51477, B2 => 
                           n53559, ZN => n59494);
   U2445 : AOI22_X1 port map( A1 => n53514, A2 => n51364, B1 => n52400, B2 => 
                           n51502, ZN => n59493);
   U2446 : AOI22_X1 port map( A1 => n53516, A2 => n51456, B1 => n53566, B2 => 
                           n51487, ZN => n59492);
   U2447 : AOI22_X1 port map( A1 => n53520, A2 => n51666, B1 => n53562, B2 => 
                           n51471, ZN => n59491);
   U2448 : NAND4_X1 port map( A1 => n59494, A2 => n59493, A3 => n59492, A4 => 
                           n59491, ZN => n59500);
   U2449 : AOI22_X1 port map( A1 => n53570, A2 => n51386, B1 => n53562, B2 => 
                           n51576, ZN => n59498);
   U2450 : AOI22_X1 port map( A1 => n53578, A2 => n51678, B1 => n53565, B2 => 
                           n51631, ZN => n59497);
   U2451 : AOI22_X1 port map( A1 => n53512, A2 => n51636, B1 => n53523, B2 => 
                           n51646, ZN => n59496);
   U2452 : AOI22_X1 port map( A1 => n53581, A2 => n51605, B1 => n53559, B2 => 
                           n51412, ZN => n59495);
   U2453 : NAND4_X1 port map( A1 => n59498, A2 => n59497, A3 => n59496, A4 => 
                           n59495, ZN => n59499);
   U2454 : AOI22_X1 port map( A1 => n59878, A2 => n59500, B1 => n59588, B2 => 
                           n59499, ZN => n59501);
   U2455 : OAI21_X1 port map( B1 => n59857, B2 => n59502, A => n59501, ZN => 
                           OUT2(25));
   U2456 : AOI22_X1 port map( A1 => n52431, A2 => n51484, B1 => n53575, B2 => 
                           n51367, ZN => n59506);
   U2457 : AOI22_X1 port map( A1 => n53586, A2 => n51530, B1 => n52422, B2 => 
                           n51369, ZN => n59505);
   U2458 : AOI22_X1 port map( A1 => n53569, A2 => n51378, B1 => n52420, B2 => 
                           n51391, ZN => n59504);
   U2459 : AOI22_X1 port map( A1 => n52425, A2 => n51654, B1 => n53563, B2 => 
                           n51408, ZN => n59503);
   U2460 : NAND4_X1 port map( A1 => n59506, A2 => n59505, A3 => n59504, A4 => 
                           n59503, ZN => n59512);
   U2461 : AOI22_X1 port map( A1 => n52427, A2 => n51595, B1 => n52419, B2 => 
                           n51625, ZN => n59510);
   U2462 : AOI22_X1 port map( A1 => n52432, A2 => n51558, B1 => n52426, B2 => 
                           n51396, ZN => n59509);
   U2463 : AOI22_X1 port map( A1 => n52423, A2 => n51543, B1 => n53587, B2 => 
                           n51443, ZN => n59508);
   U2464 : AOI22_X1 port map( A1 => n52421, A2 => n51593, B1 => n53573, B2 => 
                           n51662, ZN => n59507);
   U2465 : NAND4_X1 port map( A1 => n59510, A2 => n59509, A3 => n59508, A4 => 
                           n59507, ZN => n59511);
   U2466 : NOR2_X1 port map( A1 => n59512, A2 => n59511, ZN => n59524);
   U2467 : AOI22_X1 port map( A1 => n53516, A2 => n51473, B1 => n53559, B2 => 
                           n51499, ZN => n59516);
   U2468 : AOI22_X1 port map( A1 => n53514, A2 => n51435, B1 => n53513, B2 => 
                           n51501, ZN => n59515);
   U2469 : AOI22_X1 port map( A1 => n53583, A2 => n51504, B1 => n53570, B2 => 
                           n51554, ZN => n59514);
   U2470 : AOI22_X1 port map( A1 => n53515, A2 => n51507, B1 => n53579, B2 => 
                           n51515, ZN => n59513);
   U2471 : NAND4_X1 port map( A1 => n59516, A2 => n59515, A3 => n59514, A4 => 
                           n59513, ZN => n59522);
   U2472 : AOI22_X1 port map( A1 => n53515, A2 => n51600, B1 => n53565, B2 => 
                           n51603, ZN => n59520);
   U2473 : AOI22_X1 port map( A1 => n53579, A2 => n51584, B1 => n53559, B2 => 
                           n51380, ZN => n59519);
   U2474 : AOI22_X1 port map( A1 => n53514, A2 => n51620, B1 => n53513, B2 => 
                           n51622, ZN => n59518);
   U2475 : AOI22_X1 port map( A1 => n53582, A2 => n51384, B1 => n53583, B2 => 
                           n51609, ZN => n59517);
   U2476 : NAND4_X1 port map( A1 => n59520, A2 => n59519, A3 => n59518, A4 => 
                           n59517, ZN => n59521);
   U2477 : AOI22_X1 port map( A1 => n59878, A2 => n59522, B1 => n59588, B2 => 
                           n59521, ZN => n59523);
   U2478 : OAI21_X1 port map( B1 => n59857, B2 => n59524, A => n59523, ZN => 
                           OUT2(24));
   U2479 : AOI22_X1 port map( A1 => n52425, A2 => n51623, B1 => n53563, B2 => 
                           n51817, ZN => n59528);
   U2480 : AOI22_X1 port map( A1 => n53564, A2 => n51699, B1 => n53561, B2 => 
                           n51638, ZN => n59527);
   U2481 : AOI22_X1 port map( A1 => n52424, A2 => n51723, B1 => n53569, B2 => 
                           n51709, ZN => n59526);
   U2482 : AOI22_X1 port map( A1 => n53573, A2 => n52182, B1 => n52434, B2 => 
                           n52142, ZN => n59525);
   U2483 : NAND4_X1 port map( A1 => n59528, A2 => n59527, A3 => n59526, A4 => 
                           n59525, ZN => n59534);
   U2484 : AOI22_X1 port map( A1 => n52423, A2 => n52161, B1 => n52427, B2 => 
                           n51521, ZN => n59532);
   U2485 : AOI22_X1 port map( A1 => n53588, A2 => n52265, B1 => n53572, B2 => 
                           n51777, ZN => n59531);
   U2486 : AOI22_X1 port map( A1 => n53589, A2 => n51756, B1 => n53567, B2 => 
                           n52141, ZN => n59530);
   U2487 : AOI22_X1 port map( A1 => n53587, A2 => n51906, B1 => n53574, B2 => 
                           n51923, ZN => n59529);
   U2488 : NAND4_X1 port map( A1 => n59532, A2 => n59531, A3 => n59530, A4 => 
                           n59529, ZN => n59533);
   U2489 : NOR2_X1 port map( A1 => n59534, A2 => n59533, ZN => n59546);
   U2490 : AOI22_X1 port map( A1 => n53578, A2 => n51864, B1 => n53516, B2 => 
                           n51481, ZN => n59538);
   U2491 : AOI22_X1 port map( A1 => n53513, A2 => n51498, B1 => n53566, B2 => 
                           n51900, ZN => n59537);
   U2492 : AOI22_X1 port map( A1 => n53520, A2 => n52138, B1 => n53559, B2 => 
                           n52011, ZN => n59536);
   U2493 : AOI22_X1 port map( A1 => n52400, A2 => n51940, B1 => n53512, B2 => 
                           n51480, ZN => n59535);
   U2494 : NAND4_X1 port map( A1 => n59538, A2 => n59537, A3 => n59536, A4 => 
                           n59535, ZN => n59544);
   U2495 : AOI22_X1 port map( A1 => n53514, A2 => n52140, B1 => n53512, B2 => 
                           n52178, ZN => n59542);
   U2496 : AOI22_X1 port map( A1 => n53570, A2 => n51867, B1 => n53559, B2 => 
                           n51692, ZN => n59541);
   U2497 : AOI22_X1 port map( A1 => n53515, A2 => n52149, B1 => n52400, B2 => 
                           n52176, ZN => n59540);
   U2498 : AOI22_X1 port map( A1 => n53565, A2 => n52180, B1 => n53562, B2 => 
                           n52267, ZN => n59539);
   U2499 : NAND4_X1 port map( A1 => n59542, A2 => n59541, A3 => n59540, A4 => 
                           n59539, ZN => n59543);
   U2500 : AOI22_X1 port map( A1 => n59878, A2 => n59544, B1 => n59588, B2 => 
                           n59543, ZN => n59545);
   U2501 : OAI21_X1 port map( B1 => n60059, B2 => n59546, A => n59545, ZN => 
                           OUT2(23));
   U2502 : AOI22_X1 port map( A1 => n52431, A2 => n51903, B1 => n52424, B2 => 
                           n51722, ZN => n59550);
   U2503 : AOI22_X1 port map( A1 => n53569, A2 => n51707, B1 => n52420, B2 => 
                           n51760, ZN => n59549);
   U2504 : AOI22_X1 port map( A1 => n52432, A2 => n52172, B1 => n53588, B2 => 
                           n52264, ZN => n59548);
   U2505 : AOI22_X1 port map( A1 => n52434, A2 => n52139, B1 => n53563, B2 => 
                           n51818, ZN => n59547);
   U2506 : NAND4_X1 port map( A1 => n59550, A2 => n59549, A3 => n59548, A4 => 
                           n59547, ZN => n59556);
   U2507 : AOI22_X1 port map( A1 => n52422, A2 => n51704, B1 => n53567, B2 => 
                           n52136, ZN => n59554);
   U2508 : AOI22_X1 port map( A1 => n52423, A2 => n52171, B1 => n53587, B2 => 
                           n51445, ZN => n59553);
   U2509 : AOI22_X1 port map( A1 => n52429, A2 => n52181, B1 => n52426, B2 => 
                           n51694, ZN => n59552);
   U2510 : AOI22_X1 port map( A1 => n52425, A2 => n52174, B1 => n52427, B2 => 
                           n52127, ZN => n59551);
   U2511 : NAND4_X1 port map( A1 => n59554, A2 => n59553, A3 => n59552, A4 => 
                           n59551, ZN => n59555);
   U2512 : NOR2_X1 port map( A1 => n59556, A2 => n59555, ZN => n59568);
   U2513 : AOI22_X1 port map( A1 => n53579, A2 => n52002, B1 => n53520, B2 => 
                           n52137, ZN => n59560);
   U2514 : AOI22_X1 port map( A1 => n53514, A2 => n51866, B1 => n53565, B2 => 
                           n51958, ZN => n59559);
   U2515 : AOI22_X1 port map( A1 => n53515, A2 => n52007, B1 => n53559, B2 => 
                           n51500, ZN => n59558);
   U2516 : AOI22_X1 port map( A1 => n53513, A2 => n52010, B1 => n52400, B2 => 
                           n51495, ZN => n59557);
   U2517 : NAND4_X1 port map( A1 => n59560, A2 => n59559, A3 => n59558, A4 => 
                           n59557, ZN => n59566);
   U2518 : AOI22_X1 port map( A1 => n53514, A2 => n52124, B1 => n53583, B2 => 
                           n52175, ZN => n59564);
   U2519 : AOI22_X1 port map( A1 => n53579, A2 => n52177, B1 => n53559, B2 => 
                           n51892, ZN => n59563);
   U2520 : AOI22_X1 port map( A1 => n53584, A2 => n52179, B1 => n53577, B2 => 
                           n52268, ZN => n59562);
   U2521 : AOI22_X1 port map( A1 => n53582, A2 => n51871, B1 => n53515, B2 => 
                           n52155, ZN => n59561);
   U2522 : NAND4_X1 port map( A1 => n59564, A2 => n59563, A3 => n59562, A4 => 
                           n59561, ZN => n59565);
   U2523 : AOI22_X1 port map( A1 => n59878, A2 => n59566, B1 => n59588, B2 => 
                           n59565, ZN => n59567);
   U2524 : OAI21_X1 port map( B1 => n60059, B2 => n59568, A => n59567, ZN => 
                           OUT2(22));
   U2525 : AOI22_X1 port map( A1 => n52431, A2 => n52016, B1 => n52427, B2 => 
                           n52266, ZN => n59572);
   U2526 : AOI22_X1 port map( A1 => n52429, A2 => n52286, B1 => n52425, B2 => 
                           n52333, ZN => n59571);
   U2527 : AOI22_X1 port map( A1 => n52419, A2 => n52259, B1 => n53564, B2 => 
                           n51793, ZN => n59570);
   U2528 : AOI22_X1 port map( A1 => n53587, A2 => n52028, B1 => n52426, B2 => 
                           n51799, ZN => n59569);
   U2529 : NAND4_X1 port map( A1 => n59572, A2 => n59571, A3 => n59570, A4 => 
                           n59569, ZN => n59578);
   U2530 : AOI22_X1 port map( A1 => n52424, A2 => n51795, B1 => n52434, B2 => 
                           n51575, ZN => n59576);
   U2531 : AOI22_X1 port map( A1 => n53568, A2 => n52314, B1 => n53563, B2 => 
                           n51819, ZN => n59575);
   U2532 : AOI22_X1 port map( A1 => n53589, A2 => n51794, B1 => n52428, B2 => 
                           n51796, ZN => n59574);
   U2533 : AOI22_X1 port map( A1 => n53567, A2 => n52258, B1 => n53561, B2 => 
                           n51670, ZN => n59573);
   U2534 : NAND4_X1 port map( A1 => n59576, A2 => n59575, A3 => n59574, A4 => 
                           n59573, ZN => n59577);
   U2535 : NOR2_X1 port map( A1 => n59578, A2 => n59577, ZN => n59591);
   U2536 : AOI22_X1 port map( A1 => n53515, A2 => n51913, B1 => n53570, B2 => 
                           n51526, ZN => n59582);
   U2537 : AOI22_X1 port map( A1 => n53583, A2 => n51918, B1 => n53559, B2 => 
                           n51909, ZN => n59581);
   U2538 : AOI22_X1 port map( A1 => n53512, A2 => n51919, B1 => n53562, B2 => 
                           n51927, ZN => n59580);
   U2539 : AOI22_X1 port map( A1 => n53514, A2 => n51702, B1 => n53565, B2 => 
                           n51509, ZN => n59579);
   U2540 : NAND4_X1 port map( A1 => n59582, A2 => n59581, A3 => n59580, A4 => 
                           n59579, ZN => n59589);
   U2541 : AOI22_X1 port map( A1 => n53579, A2 => n51621, B1 => n53562, B2 => 
                           n52260, ZN => n59586);
   U2542 : AOI22_X1 port map( A1 => n53514, A2 => n52261, B1 => n53584, B2 => 
                           n52350, ZN => n59585);
   U2543 : AOI22_X1 port map( A1 => n53582, A2 => n51798, B1 => n53559, B2 => 
                           n51797, ZN => n59584);
   U2544 : AOI22_X1 port map( A1 => n53515, A2 => n51602, B1 => n52400, B2 => 
                           n51607, ZN => n59583);
   U2545 : NAND4_X1 port map( A1 => n59586, A2 => n59585, A3 => n59584, A4 => 
                           n59583, ZN => n59587);
   U2546 : AOI22_X1 port map( A1 => n59878, A2 => n59589, B1 => n59588, B2 => 
                           n59587, ZN => n59590);
   U2547 : OAI21_X1 port map( B1 => n60059, B2 => n59591, A => n59590, ZN => 
                           OUT2(21));
   U2548 : AOI22_X1 port map( A1 => n52422, A2 => n51715, B1 => n53568, B2 => 
                           n51615, ZN => n59595);
   U2549 : AOI22_X1 port map( A1 => n52419, A2 => n52263, B1 => n53561, B2 => 
                           n52168, ZN => n59594);
   U2550 : AOI22_X1 port map( A1 => n52426, A2 => n51716, B1 => n52420, B2 => 
                           n51763, ZN => n59593);
   U2551 : AOI22_X1 port map( A1 => n52425, A2 => n52173, B1 => n52427, B2 => 
                           n52128, ZN => n59592);
   U2552 : NAND4_X1 port map( A1 => n59595, A2 => n59594, A3 => n59593, A4 => 
                           n59592, ZN => n59601);
   U2553 : AOI22_X1 port map( A1 => n53587, A2 => n51920, B1 => n52431, B2 => 
                           n51921, ZN => n59599);
   U2554 : AOI22_X1 port map( A1 => n52429, A2 => n52164, B1 => n53563, B2 => 
                           n51820, ZN => n59598);
   U2555 : AOI22_X1 port map( A1 => n52421, A2 => n52143, B1 => n53575, B2 => 
                           n51714, ZN => n59597);
   U2556 : AOI22_X1 port map( A1 => n53586, A2 => n52145, B1 => n52428, B2 => 
                           n51706, ZN => n59596);
   U2557 : NAND4_X1 port map( A1 => n59599, A2 => n59598, A3 => n59597, A4 => 
                           n59596, ZN => n59600);
   U2558 : NOR2_X1 port map( A1 => n59601, A2 => n59600, ZN => n59613);
   U2559 : AOI22_X1 port map( A1 => n53562, A2 => n52000, B1 => n53559, B2 => 
                           n51999, ZN => n59605);
   U2560 : AOI22_X1 port map( A1 => n53514, A2 => n51852, B1 => n52400, B2 => 
                           n52009, ZN => n59604);
   U2561 : AOI22_X1 port map( A1 => n53516, A2 => n52006, B1 => n53570, B2 => 
                           n52152, ZN => n59603);
   U2562 : AOI22_X1 port map( A1 => n53512, A2 => n52001, B1 => n53566, B2 => 
                           n52005, ZN => n59602);
   U2563 : NAND4_X1 port map( A1 => n59605, A2 => n59604, A3 => n59603, A4 => 
                           n59602, ZN => n59611);
   U2564 : AOI22_X1 port map( A1 => n53578, A2 => n52104, B1 => n53565, B2 => 
                           n51656, ZN => n59609);
   U2565 : AOI22_X1 port map( A1 => n53523, A2 => n52206, B1 => n53562, B2 => 
                           n52269, ZN => n59608);
   U2566 : AOI22_X1 port map( A1 => n53515, A2 => n52214, B1 => n53512, B2 => 
                           n51667, ZN => n59607);
   U2567 : AOI22_X1 port map( A1 => n53570, A2 => n51800, B1 => n53559, B2 => 
                           n51893, ZN => n59606);
   U2568 : NAND4_X1 port map( A1 => n59609, A2 => n59608, A3 => n59607, A4 => 
                           n59606, ZN => n59610);
   U2569 : AOI22_X1 port map( A1 => n59878, A2 => n59611, B1 => n60054, B2 => 
                           n59610, ZN => n59612);
   U2570 : OAI21_X1 port map( B1 => n60059, B2 => n59613, A => n59612, ZN => 
                           OUT2(20));
   U2571 : AOI22_X1 port map( A1 => n52428, A2 => n51711, B1 => n53561, B2 => 
                           n52294, ZN => n59617);
   U2572 : AOI22_X1 port map( A1 => n52426, A2 => n51718, B1 => n53564, B2 => 
                           n51691, ZN => n59616);
   U2573 : AOI22_X1 port map( A1 => n52420, A2 => n51764, B1 => n53563, B2 => 
                           n51821, ZN => n59615);
   U2574 : AOI22_X1 port map( A1 => n52429, A2 => n51659, B1 => n52421, B2 => 
                           n51553, ZN => n59614);
   U2575 : NAND4_X1 port map( A1 => n59617, A2 => n59616, A3 => n59615, A4 => 
                           n59614, ZN => n59623);
   U2576 : AOI22_X1 port map( A1 => n52425, A2 => n52332, B1 => n53574, B2 => 
                           n52015, ZN => n59621);
   U2577 : AOI22_X1 port map( A1 => n52423, A2 => n52318, B1 => n52027, B2 => 
                           n52433, ZN => n59620);
   U2578 : AOI22_X1 port map( A1 => n53586, A2 => n51560, B1 => n53588, B2 => 
                           n52262, ZN => n59619);
   U2579 : AOI22_X1 port map( A1 => n53585, A2 => n51537, B1 => n52424, B2 => 
                           n51713, ZN => n59618);
   U2580 : NAND4_X1 port map( A1 => n59621, A2 => n59620, A3 => n59619, A4 => 
                           n59618, ZN => n59622);
   U2581 : NOR2_X1 port map( A1 => n59623, A2 => n59622, ZN => n59635);
   U2582 : CLKBUF_X1 port map( A => n59810, Z => n60056);
   U2583 : AOI22_X1 port map( A1 => n53512, A2 => n51926, B1 => n53565, B2 => 
                           n52067, ZN => n59627);
   U2584 : AOI22_X1 port map( A1 => n53519, A2 => n51508, B1 => n53583, B2 => 
                           n51514, ZN => n59626);
   U2585 : AOI22_X1 port map( A1 => n53515, A2 => n51512, B1 => n53570, B2 => 
                           n52371, ZN => n59625);
   U2586 : AOI22_X1 port map( A1 => n53514, A2 => n51700, B1 => n53562, B2 => 
                           n51916, ZN => n59624);
   U2587 : NAND4_X1 port map( A1 => n59627, A2 => n59626, A3 => n59625, A4 => 
                           n59624, ZN => n59633);
   U2588 : AOI22_X1 port map( A1 => n53515, A2 => n51611, B1 => n53570, B2 => 
                           n51783, ZN => n59631);
   U2589 : AOI22_X1 port map( A1 => n53519, A2 => n51894, B1 => n53512, B2 => 
                           n52340, ZN => n59630);
   U2590 : AOI22_X1 port map( A1 => n53514, A2 => n51516, B1 => n53565, B2 => 
                           n52345, ZN => n59629);
   U2591 : AOI22_X1 port map( A1 => n53523, A2 => n52343, B1 => n53562, B2 => 
                           n52270, ZN => n59628);
   U2592 : NAND4_X1 port map( A1 => n59631, A2 => n59630, A3 => n59629, A4 => 
                           n59628, ZN => n59632);
   U2593 : AOI22_X1 port map( A1 => n60056, A2 => n59633, B1 => n60054, B2 => 
                           n59632, ZN => n59634);
   U2594 : OAI21_X1 port map( B1 => n60059, B2 => n59635, A => n59634, ZN => 
                           OUT2(19));
   U2595 : AOI22_X1 port map( A1 => n53574, A2 => n52014, B1 => n52420, B2 => 
                           n51765, ZN => n59639);
   U2596 : AOI22_X1 port map( A1 => n52425, A2 => n52331, B1 => n53568, B2 => 
                           n52320, ZN => n59638);
   U2597 : AOI22_X1 port map( A1 => n53585, A2 => n52129, B1 => n52433, B2 => 
                           n52026, ZN => n59637);
   U2598 : AOI22_X1 port map( A1 => n52424, A2 => n51717, B1 => n53563, B2 => 
                           n51822, ZN => n59636);
   U2599 : NAND4_X1 port map( A1 => n59639, A2 => n59638, A3 => n59637, A4 => 
                           n59636, ZN => n59645);
   U2600 : AOI22_X1 port map( A1 => n52422, A2 => n51701, B1 => n52419, B2 => 
                           n52257, ZN => n59643);
   U2601 : AOI22_X1 port map( A1 => n52429, A2 => n52288, B1 => n52428, B2 => 
                           n51698, ZN => n59642);
   U2602 : AOI22_X1 port map( A1 => n53572, A2 => n51735, B1 => n52434, B2 => 
                           n52135, ZN => n59641);
   U2603 : AOI22_X1 port map( A1 => n52421, A2 => n51544, B1 => n53561, B2 => 
                           n52295, ZN => n59640);
   U2604 : NAND4_X1 port map( A1 => n59643, A2 => n59642, A3 => n59641, A4 => 
                           n59640, ZN => n59644);
   U2605 : NOR2_X1 port map( A1 => n59645, A2 => n59644, ZN => n59657);
   U2606 : AOI22_X1 port map( A1 => n53512, A2 => n51905, B1 => n53565, B2 => 
                           n52056, ZN => n59649);
   U2607 : AOI22_X1 port map( A1 => n53578, A2 => n51697, B1 => n53562, B2 => 
                           n51904, ZN => n59648);
   U2608 : AOI22_X1 port map( A1 => n53583, A2 => n51925, B1 => n51922, B2 => 
                           n53560, ZN => n59647);
   U2609 : AOI22_X1 port map( A1 => n53515, A2 => n51924, B1 => n53570, B2 => 
                           n52362, ZN => n59646);
   U2610 : NAND4_X1 port map( A1 => n59649, A2 => n59648, A3 => n59647, A4 => 
                           n59646, ZN => n59655);
   U2611 : AOI22_X1 port map( A1 => n53578, A2 => n51520, B1 => n53565, B2 => 
                           n51586, ZN => n59653);
   U2612 : AOI22_X1 port map( A1 => n53512, A2 => n52196, B1 => n53566, B2 => 
                           n52151, ZN => n59652);
   U2613 : AOI22_X1 port map( A1 => n53570, A2 => n51784, B1 => n53562, B2 => 
                           n52271, ZN => n59651);
   U2614 : AOI22_X1 port map( A1 => n53519, A2 => n51895, B1 => n53523, B2 => 
                           n52344, ZN => n59650);
   U2615 : NAND4_X1 port map( A1 => n59653, A2 => n59652, A3 => n59651, A4 => 
                           n59650, ZN => n59654);
   U2616 : AOI22_X1 port map( A1 => n59878, A2 => n59655, B1 => n60054, B2 => 
                           n59654, ZN => n59656);
   U2617 : OAI21_X1 port map( B1 => n60059, B2 => n59657, A => n59656, ZN => 
                           OUT2(18));
   U2618 : AOI22_X1 port map( A1 => n53561, A2 => n52296, B1 => n52433, B2 => 
                           n52024, ZN => n59661);
   U2619 : AOI22_X1 port map( A1 => n52421, A2 => n52251, B1 => n52434, B2 => 
                           n52225, ZN => n59660);
   U2620 : AOI22_X1 port map( A1 => n52423, A2 => n52299, B1 => n52427, B2 => 
                           n52224, ZN => n59659);
   U2621 : AOI22_X1 port map( A1 => n52422, A2 => n51802, B1 => n52430, B2 => 
                           n51814, ZN => n59658);
   U2622 : NAND4_X1 port map( A1 => n59661, A2 => n59660, A3 => n59659, A4 => 
                           n59658, ZN => n59667);
   U2623 : AOI22_X1 port map( A1 => n53589, A2 => n51803, B1 => n52431, B2 => 
                           n52013, ZN => n59665);
   U2624 : AOI22_X1 port map( A1 => n52429, A2 => n52292, B1 => n52424, B2 => 
                           n51804, ZN => n59664);
   U2625 : AOI22_X1 port map( A1 => n52425, A2 => n52326, B1 => n52428, B2 => 
                           n51805, ZN => n59663);
   U2626 : AOI22_X1 port map( A1 => n52426, A2 => n51808, B1 => n52419, B2 => 
                           n51590, ZN => n59662);
   U2627 : NAND4_X1 port map( A1 => n59665, A2 => n59664, A3 => n59663, A4 => 
                           n59662, ZN => n59666);
   U2628 : NOR2_X1 port map( A1 => n59667, A2 => n59666, ZN => n59679);
   U2629 : AOI22_X1 port map( A1 => n53570, A2 => n52330, B1 => n53566, B2 => 
                           n51960, ZN => n59671);
   U2630 : AOI22_X1 port map( A1 => n53583, A2 => n51971, B1 => n53513, B2 => 
                           n51965, ZN => n59670);
   U2631 : AOI22_X1 port map( A1 => n53519, A2 => n51962, B1 => n53578, B2 => 
                           n51766, ZN => n59669);
   U2632 : AOI22_X1 port map( A1 => n53516, A2 => n52061, B1 => n53512, B2 => 
                           n51970, ZN => n59668);
   U2633 : NAND4_X1 port map( A1 => n59671, A2 => n59670, A3 => n59669, A4 => 
                           n59668, ZN => n59677);
   U2634 : AOI22_X1 port map( A1 => n53515, A2 => n52213, B1 => n53523, B2 => 
                           n52209, ZN => n59675);
   U2635 : AOI22_X1 port map( A1 => n53513, A2 => n51585, B1 => n53512, B2 => 
                           n52200, ZN => n59674);
   U2636 : AOI22_X1 port map( A1 => n53519, A2 => n51806, B1 => n53570, B2 => 
                           n51807, ZN => n59673);
   U2637 : AOI22_X1 port map( A1 => n53578, A2 => n52221, B1 => n53565, B2 => 
                           n52240, ZN => n59672);
   U2638 : NAND4_X1 port map( A1 => n59675, A2 => n59674, A3 => n59673, A4 => 
                           n59672, ZN => n59676);
   U2639 : AOI22_X1 port map( A1 => n60056, A2 => n59677, B1 => n60054, B2 => 
                           n59676, ZN => n59678);
   U2640 : OAI21_X1 port map( B1 => n60059, B2 => n59679, A => n59678, ZN => 
                           OUT2(17));
   U2641 : AOI22_X1 port map( A1 => n52421, A2 => n52169, B1 => n52433, B2 => 
                           n52023, ZN => n59683);
   U2642 : AOI22_X1 port map( A1 => n52432, A2 => n52297, B1 => n53589, B2 => 
                           n51811, ZN => n59682);
   U2643 : AOI22_X1 port map( A1 => n52422, A2 => n51813, B1 => n52430, B2 => 
                           n51824, ZN => n59681);
   U2644 : AOI22_X1 port map( A1 => n52425, A2 => n52324, B1 => n53574, B2 => 
                           n52025, ZN => n59680);
   U2645 : NAND4_X1 port map( A1 => n59683, A2 => n59682, A3 => n59681, A4 => 
                           n59680, ZN => n59689);
   U2646 : AOI22_X1 port map( A1 => n53585, A2 => n52185, B1 => n53572, B2 => 
                           n51812, ZN => n59687);
   U2647 : AOI22_X1 port map( A1 => n52429, A2 => n52133, B1 => n53575, B2 => 
                           n51815, ZN => n59686);
   U2648 : AOI22_X1 port map( A1 => n52423, A2 => n51527, B1 => n52434, B2 => 
                           n52170, ZN => n59685);
   U2649 : AOI22_X1 port map( A1 => n52428, A2 => n51816, B1 => n53588, B2 => 
                           n51619, ZN => n59684);
   U2650 : NAND4_X1 port map( A1 => n59687, A2 => n59686, A3 => n59685, A4 => 
                           n59684, ZN => n59688);
   U2651 : NOR2_X1 port map( A1 => n59689, A2 => n59688, ZN => n59701);
   U2652 : AOI22_X1 port map( A1 => n53512, A2 => n52069, B1 => n53570, B2 => 
                           n52309, ZN => n59693);
   U2653 : AOI22_X1 port map( A1 => n52400, A2 => n52070, B1 => n53565, B2 => 
                           n51964, ZN => n59692);
   U2654 : AOI22_X1 port map( A1 => n53515, A2 => n52071, B1 => n53578, B2 => 
                           n51696, ZN => n59691);
   U2655 : AOI22_X1 port map( A1 => n53519, A2 => n52072, B1 => n53513, B2 => 
                           n52073, ZN => n59690);
   U2656 : NAND4_X1 port map( A1 => n59693, A2 => n59692, A3 => n59691, A4 => 
                           n59690, ZN => n59699);
   U2657 : AOI22_X1 port map( A1 => n53583, A2 => n51599, B1 => n53562, B2 => 
                           n52195, ZN => n59697);
   U2658 : AOI22_X1 port map( A1 => n53519, A2 => n51809, B1 => n53520, B2 => 
                           n51810, ZN => n59696);
   U2659 : AOI22_X1 port map( A1 => n53578, A2 => n52197, B1 => n53565, B2 => 
                           n52349, ZN => n59695);
   U2660 : AOI22_X1 port map( A1 => n53515, A2 => n52154, B1 => n53512, B2 => 
                           n52337, ZN => n59694);
   U2661 : NAND4_X1 port map( A1 => n59697, A2 => n59696, A3 => n59695, A4 => 
                           n59694, ZN => n59698);
   U2662 : AOI22_X1 port map( A1 => n60056, A2 => n59699, B1 => n60054, B2 => 
                           n59698, ZN => n59700);
   U2663 : OAI21_X1 port map( B1 => n60059, B2 => n59701, A => n59700, ZN => 
                           OUT2(16));
   U2664 : AOI22_X1 port map( A1 => n52430, A2 => n51823, B1 => n52426, B2 => 
                           n51736, ZN => n59705);
   U2665 : AOI22_X1 port map( A1 => n52423, A2 => n52319, B1 => n52429, B2 => 
                           n52293, ZN => n59704);
   U2666 : AOI22_X1 port map( A1 => n52432, A2 => n52298, B1 => n52427, B2 => 
                           n52111, ZN => n59703);
   U2667 : AOI22_X1 port map( A1 => n53564, A2 => n51738, B1 => n52433, B2 => 
                           n52022, ZN => n59702);
   U2668 : NAND4_X1 port map( A1 => n59705, A2 => n59704, A3 => n59703, A4 => 
                           n59702, ZN => n59711);
   U2669 : AOI22_X1 port map( A1 => n52425, A2 => n51541, B1 => n52420, B2 => 
                           n51767, ZN => n59709);
   U2670 : AOI22_X1 port map( A1 => n52421, A2 => n52125, B1 => n53588, B2 => 
                           n52256, ZN => n59708);
   U2671 : AOI22_X1 port map( A1 => n52428, A2 => n51737, B1 => n52434, B2 => 
                           n52121, ZN => n59707);
   U2672 : AOI22_X1 port map( A1 => n52431, A2 => n52012, B1 => n53575, B2 => 
                           n51734, ZN => n59706);
   U2673 : NAND4_X1 port map( A1 => n59709, A2 => n59708, A3 => n59707, A4 => 
                           n59706, ZN => n59710);
   U2674 : NOR2_X1 port map( A1 => n59711, A2 => n59710, ZN => n59723);
   U2675 : AOI22_X1 port map( A1 => n53566, A2 => n51899, B1 => n53565, B2 => 
                           n52047, ZN => n59715);
   U2676 : AOI22_X1 port map( A1 => n53578, A2 => n51725, B1 => n53523, B2 => 
                           n51915, ZN => n59714);
   U2677 : AOI22_X1 port map( A1 => n53580, A2 => n51938, B1 => n53577, B2 => 
                           n51928, ZN => n59713);
   U2678 : AOI22_X1 port map( A1 => n53520, A2 => n52306, B1 => n53559, B2 => 
                           n51914, ZN => n59712);
   U2679 : NAND4_X1 port map( A1 => n59715, A2 => n59714, A3 => n59713, A4 => 
                           n59712, ZN => n59721);
   U2680 : AOI22_X1 port map( A1 => n53515, A2 => n52217, B1 => n53562, B2 => 
                           n51532, ZN => n59719);
   U2681 : AOI22_X1 port map( A1 => n53578, A2 => n52284, B1 => n53565, B2 => 
                           n52243, ZN => n59718);
   U2682 : AOI22_X1 port map( A1 => n53579, A2 => n52201, B1 => n53570, B2 => 
                           n51785, ZN => n59717);
   U2683 : AOI22_X1 port map( A1 => n53519, A2 => n51896, B1 => n53523, B2 => 
                           n52241, ZN => n59716);
   U2684 : NAND4_X1 port map( A1 => n59719, A2 => n59718, A3 => n59717, A4 => 
                           n59716, ZN => n59720);
   U2685 : AOI22_X1 port map( A1 => n59878, A2 => n59721, B1 => n60054, B2 => 
                           n59720, ZN => n59722);
   U2686 : OAI21_X1 port map( B1 => n60059, B2 => n59723, A => n59722, ZN => 
                           OUT2(15));
   U2687 : AOI22_X1 port map( A1 => n52422, A2 => n51747, B1 => n52421, B2 => 
                           n52144, ZN => n59727);
   U2688 : AOI22_X1 port map( A1 => n52432, A2 => n52300, B1 => n52427, B2 => 
                           n52131, ZN => n59726);
   U2689 : AOI22_X1 port map( A1 => n53576, A2 => n52323, B1 => n52419, B2 => 
                           n52255, ZN => n59725);
   U2690 : AOI22_X1 port map( A1 => n53586, A2 => n52146, B1 => n52429, B2 => 
                           n52291, ZN => n59724);
   U2691 : NAND4_X1 port map( A1 => n59727, A2 => n59726, A3 => n59725, A4 => 
                           n59724, ZN => n59733);
   U2692 : AOI22_X1 port map( A1 => n53589, A2 => n51768, B1 => n52433, B2 => 
                           n52021, ZN => n59731);
   U2693 : AOI22_X1 port map( A1 => n52431, A2 => n51482, B1 => n52424, B2 => 
                           n51710, ZN => n59730);
   U2694 : AOI22_X1 port map( A1 => n52423, A2 => n52312, B1 => n52426, B2 => 
                           n51739, ZN => n59729);
   U2695 : AOI22_X1 port map( A1 => n52428, A2 => n51703, B1 => n52430, B2 => 
                           n51826, ZN => n59728);
   U2696 : NAND4_X1 port map( A1 => n59731, A2 => n59730, A3 => n59729, A4 => 
                           n59728, ZN => n59732);
   U2697 : NOR2_X1 port map( A1 => n59733, A2 => n59732, ZN => n59745);
   U2698 : AOI22_X1 port map( A1 => n53520, A2 => n52387, B1 => n53566, B2 => 
                           n52049, ZN => n59737);
   U2699 : AOI22_X1 port map( A1 => n53579, A2 => n52046, B1 => n53562, B2 => 
                           n51483, ZN => n59736);
   U2700 : AOI22_X1 port map( A1 => n53584, A2 => n51956, B1 => n53523, B2 => 
                           n52045, ZN => n59735);
   U2701 : AOI22_X1 port map( A1 => n53578, A2 => n51720, B1 => n53559, B2 => 
                           n52048, ZN => n59734);
   U2702 : NAND4_X1 port map( A1 => n59737, A2 => n59736, A3 => n59735, A4 => 
                           n59734, ZN => n59743);
   U2703 : AOI22_X1 port map( A1 => n53519, A2 => n51897, B1 => n53520, B2 => 
                           n51786, ZN => n59741);
   U2704 : AOI22_X1 port map( A1 => n53512, A2 => n52190, B1 => n53565, B2 => 
                           n52192, ZN => n59740);
   U2705 : AOI22_X1 port map( A1 => n53578, A2 => n52283, B1 => n53523, B2 => 
                           n52348, ZN => n59739);
   U2706 : AOI22_X1 port map( A1 => n53577, A2 => n52272, B1 => n53566, B2 => 
                           n52147, ZN => n59738);
   U2707 : NAND4_X1 port map( A1 => n59741, A2 => n59740, A3 => n59739, A4 => 
                           n59738, ZN => n59742);
   U2708 : AOI22_X1 port map( A1 => n59878, A2 => n59743, B1 => n60054, B2 => 
                           n59742, ZN => n59744);
   U2709 : OAI21_X1 port map( B1 => n60059, B2 => n59745, A => n59744, ZN => 
                           OUT2(14));
   U2710 : AOI22_X1 port map( A1 => n52423, A2 => n52311, B1 => n52421, B2 => 
                           n52080, ZN => n59749);
   U2711 : AOI22_X1 port map( A1 => n53589, A2 => n51769, B1 => n53564, B2 => 
                           n51750, ZN => n59748);
   U2712 : AOI22_X1 port map( A1 => n52431, A2 => n52029, B1 => n52426, B2 => 
                           n51740, ZN => n59747);
   U2713 : AOI22_X1 port map( A1 => n52429, A2 => n52290, B1 => n52427, B2 => 
                           n52088, ZN => n59746);
   U2714 : NAND4_X1 port map( A1 => n59749, A2 => n59748, A3 => n59747, A4 => 
                           n59746, ZN => n59755);
   U2715 : AOI22_X1 port map( A1 => n52430, A2 => n51825, B1 => n52424, B2 => 
                           n51753, ZN => n59753);
   U2716 : AOI22_X1 port map( A1 => n52434, A2 => n52076, B1 => n52433, B2 => 
                           n52020, ZN => n59752);
   U2717 : AOI22_X1 port map( A1 => n52432, A2 => n52301, B1 => n52428, B2 => 
                           n51755, ZN => n59751);
   U2718 : AOI22_X1 port map( A1 => n53576, A2 => n52322, B1 => n52419, B2 => 
                           n52254, ZN => n59750);
   U2719 : NAND4_X1 port map( A1 => n59753, A2 => n59752, A3 => n59751, A4 => 
                           n59750, ZN => n59754);
   U2720 : NOR2_X1 port map( A1 => n59755, A2 => n59754, ZN => n59767);
   U2721 : AOI22_X1 port map( A1 => n53581, A2 => n51510, B1 => n53583, B2 => 
                           n52053, ZN => n59759);
   U2722 : AOI22_X1 port map( A1 => n53582, A2 => n52347, B1 => n53513, B2 => 
                           n52050, ZN => n59758);
   U2723 : AOI22_X1 port map( A1 => n53516, A2 => n52051, B1 => n53560, B2 => 
                           n52054, ZN => n59757);
   U2724 : AOI22_X1 port map( A1 => n53580, A2 => n52052, B1 => n53514, B2 => 
                           n51712, ZN => n59756);
   U2725 : NAND4_X1 port map( A1 => n59759, A2 => n59758, A3 => n59757, A4 => 
                           n59756, ZN => n59765);
   U2726 : AOI22_X1 port map( A1 => n53582, A2 => n51787, B1 => n53571, B2 => 
                           n52282, ZN => n59763);
   U2727 : AOI22_X1 port map( A1 => n53577, A2 => n52273, B1 => n53515, B2 => 
                           n52153, ZN => n59762);
   U2728 : AOI22_X1 port map( A1 => n53580, A2 => n52353, B1 => n53565, B2 => 
                           n52346, ZN => n59761);
   U2729 : AOI22_X1 port map( A1 => n53523, A2 => n52357, B1 => n53560, B2 => 
                           n51898, ZN => n59760);
   U2730 : NAND4_X1 port map( A1 => n59763, A2 => n59762, A3 => n59761, A4 => 
                           n59760, ZN => n59764);
   U2731 : AOI22_X1 port map( A1 => n59878, A2 => n59765, B1 => n60054, B2 => 
                           n59764, ZN => n59766);
   U2732 : OAI21_X1 port map( B1 => n60059, B2 => n59767, A => n59766, ZN => 
                           OUT2(13));
   U2733 : AOI22_X1 port map( A1 => n53574, A2 => n51476, B1 => n52420, B2 => 
                           n51770, ZN => n59771);
   U2734 : AOI22_X1 port map( A1 => n52430, A2 => n51829, B1 => n52433, B2 => 
                           n51449, ZN => n59770);
   U2735 : AOI22_X1 port map( A1 => n52428, A2 => n51759, B1 => n53568, B2 => 
                           n52321, ZN => n59769);
   U2736 : AOI22_X1 port map( A1 => n52429, A2 => n51669, B1 => n53588, B2 => 
                           n52253, ZN => n59768);
   U2737 : NAND4_X1 port map( A1 => n59771, A2 => n59770, A3 => n59769, A4 => 
                           n59768, ZN => n59777);
   U2738 : AOI22_X1 port map( A1 => n52421, A2 => n52085, B1 => n52427, B2 => 
                           n52092, ZN => n59775);
   U2739 : AOI22_X1 port map( A1 => n53586, A2 => n52090, B1 => n53576, B2 => 
                           n52316, ZN => n59774);
   U2740 : AOI22_X1 port map( A1 => n52422, A2 => n51757, B1 => n52432, B2 => 
                           n52302, ZN => n59773);
   U2741 : AOI22_X1 port map( A1 => n52424, A2 => n51758, B1 => n53572, B2 => 
                           n51741, ZN => n59772);
   U2742 : NAND4_X1 port map( A1 => n59775, A2 => n59774, A3 => n59773, A4 => 
                           n59772, ZN => n59776);
   U2743 : NOR2_X1 port map( A1 => n59777, A2 => n59776, ZN => n59789);
   U2744 : AOI22_X1 port map( A1 => n53513, A2 => n52055, B1 => n53566, B2 => 
                           n52059, ZN => n59781);
   U2745 : AOI22_X1 port map( A1 => n53580, A2 => n51513, B1 => n53560, B2 => 
                           n52060, ZN => n59780);
   U2746 : AOI22_X1 port map( A1 => n53583, A2 => n52058, B1 => n53578, B2 => 
                           n51705, ZN => n59779);
   U2747 : AOI22_X1 port map( A1 => n53516, A2 => n52057, B1 => n53520, B2 => 
                           n51632, ZN => n59778);
   U2748 : NAND4_X1 port map( A1 => n59781, A2 => n59780, A3 => n59779, A4 => 
                           n59778, ZN => n59787);
   U2749 : AOI22_X1 port map( A1 => n53580, A2 => n52188, B1 => n53571, B2 => 
                           n52281, ZN => n59785);
   U2750 : AOI22_X1 port map( A1 => n53583, A2 => n52351, B1 => n53516, B2 => 
                           n52189, ZN => n59784);
   U2751 : AOI22_X1 port map( A1 => n53582, A2 => n51788, B1 => n53560, B2 => 
                           n51778, ZN => n59783);
   U2752 : AOI22_X1 port map( A1 => n53581, A2 => n52159, B1 => n53513, B2 => 
                           n52274, ZN => n59782);
   U2753 : NAND4_X1 port map( A1 => n59785, A2 => n59784, A3 => n59783, A4 => 
                           n59782, ZN => n59786);
   U2754 : AOI22_X1 port map( A1 => n59878, A2 => n59787, B1 => n60054, B2 => 
                           n59786, ZN => n59788);
   U2755 : OAI21_X1 port map( B1 => n60059, B2 => n59789, A => n59788, ZN => 
                           OUT2(12));
   U2756 : AOI22_X1 port map( A1 => n52423, A2 => n52313, B1 => n52432, B2 => 
                           n52303, ZN => n59793);
   U2757 : AOI22_X1 port map( A1 => n52425, A2 => n52328, B1 => n53575, B2 => 
                           n51773, ZN => n59792);
   U2758 : AOI22_X1 port map( A1 => n53574, A2 => n52030, B1 => n52420, B2 => 
                           n51772, ZN => n59791);
   U2759 : AOI22_X1 port map( A1 => n52421, A2 => n52095, B1 => n53572, B2 => 
                           n51742, ZN => n59790);
   U2760 : NAND4_X1 port map( A1 => n59793, A2 => n59792, A3 => n59791, A4 => 
                           n59790, ZN => n59799);
   U2761 : AOI22_X1 port map( A1 => n52434, A2 => n52098, B1 => n52419, B2 => 
                           n52252, ZN => n59797);
   U2762 : AOI22_X1 port map( A1 => n53564, A2 => n51771, B1 => n52433, B2 => 
                           n52019, ZN => n59796);
   U2763 : AOI22_X1 port map( A1 => n52429, A2 => n52289, B1 => n52430, B2 => 
                           n51801, ZN => n59795);
   U2764 : AOI22_X1 port map( A1 => n52428, A2 => n51774, B1 => n53585, B2 => 
                           n52109, ZN => n59794);
   U2765 : NAND4_X1 port map( A1 => n59797, A2 => n59796, A3 => n59795, A4 => 
                           n59794, ZN => n59798);
   U2766 : NOR2_X1 port map( A1 => n59799, A2 => n59798, ZN => n59812);
   U2767 : AOI22_X1 port map( A1 => n53579, A2 => n52064, B1 => n53560, B2 => 
                           n52068, ZN => n59803);
   U2768 : AOI22_X1 port map( A1 => n53581, A2 => n52066, B1 => n53571, B2 => 
                           n51695, ZN => n59802);
   U2769 : AOI22_X1 port map( A1 => n53584, A2 => n52063, B1 => n53583, B2 => 
                           n52065, ZN => n59801);
   U2770 : AOI22_X1 port map( A1 => n53582, A2 => n52382, B1 => n53577, B2 => 
                           n52062, ZN => n59800);
   U2771 : NAND4_X1 port map( A1 => n59803, A2 => n59802, A3 => n59801, A4 => 
                           n59800, ZN => n59809);
   U2772 : AOI22_X1 port map( A1 => n53581, A2 => n52157, B1 => n53579, B2 => 
                           n52355, ZN => n59807);
   U2773 : AOI22_X1 port map( A1 => n53513, A2 => n52275, B1 => n53578, B2 => 
                           n52278, ZN => n59806);
   U2774 : AOI22_X1 port map( A1 => n53583, A2 => n52352, B1 => n53560, B2 => 
                           n51779, ZN => n59805);
   U2775 : AOI22_X1 port map( A1 => n53516, A2 => n52339, B1 => n53520, B2 => 
                           n51789, ZN => n59804);
   U2776 : NAND4_X1 port map( A1 => n59807, A2 => n59806, A3 => n59805, A4 => 
                           n59804, ZN => n59808);
   U2777 : AOI22_X1 port map( A1 => n59810, A2 => n59809, B1 => n60054, B2 => 
                           n59808, ZN => n59811);
   U2778 : OAI21_X1 port map( B1 => n59857, B2 => n59812, A => n59811, ZN => 
                           OUT2(11));
   U2779 : AOI22_X1 port map( A1 => n52428, A2 => n51752, B1 => n52421, B2 => 
                           n52112, ZN => n59816);
   U2780 : AOI22_X1 port map( A1 => n52425, A2 => n51582, B1 => n53575, B2 => 
                           n51754, ZN => n59815);
   U2781 : AOI22_X1 port map( A1 => n53585, A2 => n51562, B1 => n52419, B2 => 
                           n51578, ZN => n59814);
   U2782 : AOI22_X1 port map( A1 => n52423, A2 => n52360, B1 => n52420, B2 => 
                           n51761, ZN => n59813);
   U2783 : NAND4_X1 port map( A1 => n59816, A2 => n59815, A3 => n59814, A4 => 
                           n59813, ZN => n59822);
   U2784 : AOI22_X1 port map( A1 => n52422, A2 => n51726, B1 => n52429, B2 => 
                           n51581, ZN => n59820);
   U2785 : AOI22_X1 port map( A1 => n52431, A2 => n51998, B1 => n52426, B2 => 
                           n51744, ZN => n59819);
   U2786 : AOI22_X1 port map( A1 => n53586, A2 => n52160, B1 => n52430, B2 => 
                           n51733, ZN => n59818);
   U2787 : AOI22_X1 port map( A1 => n52432, A2 => n51579, B1 => n52433, B2 => 
                           n51997, ZN => n59817);
   U2788 : NAND4_X1 port map( A1 => n59820, A2 => n59819, A3 => n59818, A4 => 
                           n59817, ZN => n59821);
   U2789 : NOR2_X1 port map( A1 => n59822, A2 => n59821, ZN => n59834);
   U2790 : AOI22_X1 port map( A1 => n53580, A2 => n51981, B1 => n53560, B2 => 
                           n51974, ZN => n59826);
   U2791 : AOI22_X1 port map( A1 => n53513, A2 => n51969, B1 => n53571, B2 => 
                           n51833, ZN => n59825);
   U2792 : AOI22_X1 port map( A1 => n53520, A2 => n52162, B1 => n53566, B2 => 
                           n51972, ZN => n59824);
   U2793 : AOI22_X1 port map( A1 => n53583, A2 => n51976, B1 => n53516, B2 => 
                           n51978, ZN => n59823);
   U2794 : NAND4_X1 port map( A1 => n59826, A2 => n59825, A3 => n59824, A4 => 
                           n59823, ZN => n59832);
   U2795 : AOI22_X1 port map( A1 => n53571, A2 => n51626, B1 => n53566, B2 => 
                           n51601, ZN => n59830);
   U2796 : AOI22_X1 port map( A1 => n53513, A2 => n52163, B1 => n53523, B2 => 
                           n52358, ZN => n59829);
   U2797 : AOI22_X1 port map( A1 => n53516, A2 => n51608, B1 => n53520, B2 => 
                           n51792, ZN => n59828);
   U2798 : AOI22_X1 port map( A1 => n53580, A2 => n51616, B1 => n53560, B2 => 
                           n51780, ZN => n59827);
   U2799 : NAND4_X1 port map( A1 => n59830, A2 => n59829, A3 => n59828, A4 => 
                           n59827, ZN => n59831);
   U2800 : AOI22_X1 port map( A1 => n59878, A2 => n59832, B1 => n60054, B2 => 
                           n59831, ZN => n59833);
   U2801 : OAI21_X1 port map( B1 => n59857, B2 => n59834, A => n59833, ZN => 
                           OUT2(10));
   U2802 : AOI22_X1 port map( A1 => n52432, A2 => n52304, B1 => n52433, B2 => 
                           n52018, ZN => n59838);
   U2803 : AOI22_X1 port map( A1 => n53585, A2 => n52126, B1 => n52426, B2 => 
                           n51745, ZN => n59837);
   U2804 : AOI22_X1 port map( A1 => n52423, A2 => n51545, B1 => n52420, B2 => 
                           n51775, ZN => n59836);
   U2805 : AOI22_X1 port map( A1 => n53574, A2 => n52031, B1 => n53576, B2 => 
                           n52327, ZN => n59835);
   U2806 : NAND4_X1 port map( A1 => n59838, A2 => n59837, A3 => n59836, A4 => 
                           n59835, ZN => n59844);
   U2807 : AOI22_X1 port map( A1 => n52424, A2 => n51730, B1 => n52419, B2 => 
                           n52223, ZN => n59842);
   U2808 : AOI22_X1 port map( A1 => n52428, A2 => n51751, B1 => n53564, B2 => 
                           n51748, ZN => n59841);
   U2809 : AOI22_X1 port map( A1 => n53586, A2 => n51533, B1 => n52421, B2 => 
                           n51539, ZN => n59840);
   U2810 : AOI22_X1 port map( A1 => n52429, A2 => n52287, B1 => n52430, B2 => 
                           n51729, ZN => n59839);
   U2811 : NAND4_X1 port map( A1 => n59842, A2 => n59841, A3 => n59840, A4 => 
                           n59839, ZN => n59843);
   U2812 : NOR2_X1 port map( A1 => n59844, A2 => n59843, ZN => n59856);
   U2813 : AOI22_X1 port map( A1 => n53514, A2 => n51731, B1 => n53560, B2 => 
                           n52036, ZN => n59848);
   U2814 : AOI22_X1 port map( A1 => n53580, A2 => n52037, B1 => n53582, B2 => 
                           n51552, ZN => n59847);
   U2815 : AOI22_X1 port map( A1 => n53581, A2 => n52034, B1 => n53583, B2 => 
                           n52035, ZN => n59846);
   U2816 : AOI22_X1 port map( A1 => n53513, A2 => n52038, B1 => n53516, B2 => 
                           n52033, ZN => n59845);
   U2817 : NAND4_X1 port map( A1 => n59848, A2 => n59847, A3 => n59846, A4 => 
                           n59845, ZN => n59854);
   U2818 : AOI22_X1 port map( A1 => n53581, A2 => n52148, B1 => n53523, B2 => 
                           n51592, ZN => n59852);
   U2819 : AOI22_X1 port map( A1 => n53582, A2 => n51791, B1 => n53560, B2 => 
                           n51781, ZN => n59851);
   U2820 : AOI22_X1 port map( A1 => n53580, A2 => n52193, B1 => n53571, B2 => 
                           n52277, ZN => n59850);
   U2821 : AOI22_X1 port map( A1 => n53577, A2 => n52279, B1 => n53516, B2 => 
                           n52359, ZN => n59849);
   U2822 : NAND4_X1 port map( A1 => n59852, A2 => n59851, A3 => n59850, A4 => 
                           n59849, ZN => n59853);
   U2823 : AOI22_X1 port map( A1 => n59878, A2 => n59854, B1 => n60054, B2 => 
                           n59853, ZN => n59855);
   U2824 : OAI21_X1 port map( B1 => n59857, B2 => n59856, A => n59855, ZN => 
                           OUT2(9));
   U2825 : AOI22_X1 port map( A1 => n52423, A2 => n52329, B1 => n52429, B2 => 
                           n52334, ZN => n59861);
   U2826 : AOI22_X1 port map( A1 => n52430, A2 => n51719, B1 => n52433, B2 => 
                           n52017, ZN => n59860);
   U2827 : AOI22_X1 port map( A1 => n52426, A2 => n51746, B1 => n52419, B2 => 
                           n52222, ZN => n59859);
   U2828 : AOI22_X1 port map( A1 => n52422, A2 => n51749, B1 => n52428, B2 => 
                           n51727, ZN => n59858);
   U2829 : NAND4_X1 port map( A1 => n59861, A2 => n59860, A3 => n59859, A4 => 
                           n59858, ZN => n59867);
   U2830 : AOI22_X1 port map( A1 => n52424, A2 => n51728, B1 => n52434, B2 => 
                           n52134, ZN => n59865);
   U2831 : AOI22_X1 port map( A1 => n53576, A2 => n52325, B1 => n52420, B2 => 
                           n51776, ZN => n59864);
   U2832 : AOI22_X1 port map( A1 => n52421, A2 => n52132, B1 => n52427, B2 => 
                           n52130, ZN => n59863);
   U2833 : AOI22_X1 port map( A1 => n52432, A2 => n52305, B1 => n52431, B2 => 
                           n52032, ZN => n59862);
   U2834 : NAND4_X1 port map( A1 => n59865, A2 => n59864, A3 => n59863, A4 => 
                           n59862, ZN => n59866);
   U2835 : NOR2_X1 port map( A1 => n59867, A2 => n59866, ZN => n59880);
   U2836 : AOI22_X1 port map( A1 => n53580, A2 => n52043, B1 => n53513, B2 => 
                           n52039, ZN => n59871);
   U2837 : AOI22_X1 port map( A1 => n53516, A2 => n52042, B1 => n53560, B2 => 
                           n52040, ZN => n59870);
   U2838 : AOI22_X1 port map( A1 => n53520, A2 => n52307, B1 => n53523, B2 => 
                           n52041, ZN => n59869);
   U2839 : AOI22_X1 port map( A1 => n53581, A2 => n52044, B1 => n53571, B2 => 
                           n51724, ZN => n59868);
   U2840 : NAND4_X1 port map( A1 => n59871, A2 => n59870, A3 => n59869, A4 => 
                           n59868, ZN => n59877);
   U2841 : AOI22_X1 port map( A1 => n53582, A2 => n51790, B1 => n53560, B2 => 
                           n51782, ZN => n59875);
   U2842 : AOI22_X1 port map( A1 => n53580, A2 => n52191, B1 => n52400, B2 => 
                           n52356, ZN => n59874);
   U2843 : AOI22_X1 port map( A1 => n53571, A2 => n52276, B1 => n53562, B2 => 
                           n52280, ZN => n59873);
   U2844 : AOI22_X1 port map( A1 => n53581, A2 => n52150, B1 => n53516, B2 => 
                           n52194, ZN => n59872);
   U2845 : NAND4_X1 port map( A1 => n59875, A2 => n59874, A3 => n59873, A4 => 
                           n59872, ZN => n59876);
   U2846 : AOI22_X1 port map( A1 => n59878, A2 => n59877, B1 => n60054, B2 => 
                           n59876, ZN => n59879);
   U2847 : OAI21_X1 port map( B1 => n60059, B2 => n59880, A => n59879, ZN => 
                           OUT2(8));
   U2848 : AOI22_X1 port map( A1 => n52429, A2 => n52183, B1 => n52433, B2 => 
                           n51968, ZN => n59884);
   U2849 : AOI22_X1 port map( A1 => n52425, A2 => n52187, B1 => n52428, B2 => 
                           n51888, ZN => n59883);
   U2850 : AOI22_X1 port map( A1 => n52431, A2 => n51967, B1 => n53568, B2 => 
                           n52184, ZN => n59882);
   U2851 : AOI22_X1 port map( A1 => n52421, A2 => n52117, B1 => n52419, B2 => 
                           n52083, ZN => n59881);
   U2852 : NAND4_X1 port map( A1 => n59884, A2 => n59883, A3 => n59882, A4 => 
                           n59881, ZN => n59890);
   U2853 : AOI22_X1 port map( A1 => n52426, A2 => n51874, B1 => n53564, B2 => 
                           n51891, ZN => n59888);
   U2854 : AOI22_X1 port map( A1 => n53585, A2 => n52091, B1 => n52420, B2 => 
                           n51881, ZN => n59887);
   U2855 : AOI22_X1 port map( A1 => n52424, A2 => n51887, B1 => n52434, B2 => 
                           n52123, ZN => n59886);
   U2856 : AOI22_X1 port map( A1 => n52432, A2 => n52186, B1 => n52430, B2 => 
                           n51863, ZN => n59885);
   U2857 : NAND4_X1 port map( A1 => n59888, A2 => n59887, A3 => n59886, A4 => 
                           n59885, ZN => n59889);
   U2858 : NOR2_X1 port map( A1 => n59890, A2 => n59889, ZN => n59902);
   U2859 : AOI22_X1 port map( A1 => n53581, A2 => n52004, B1 => n52400, B2 => 
                           n52003, ZN => n59894);
   U2860 : AOI22_X1 port map( A1 => n53582, A2 => n52156, B1 => n53513, B2 => 
                           n51994, ZN => n59893);
   U2861 : AOI22_X1 port map( A1 => n53571, A2 => n51851, B1 => n53560, B2 => 
                           n51983, ZN => n59892);
   U2862 : AOI22_X1 port map( A1 => n53580, A2 => n51996, B1 => n53516, B2 => 
                           n52008, ZN => n59891);
   U2863 : NAND4_X1 port map( A1 => n59894, A2 => n59893, A3 => n59892, A4 => 
                           n59891, ZN => n59900);
   U2864 : AOI22_X1 port map( A1 => n53578, A2 => n52208, B1 => n53566, B2 => 
                           n52219, ZN => n59898);
   U2865 : AOI22_X1 port map( A1 => n53580, A2 => n52249, B1 => n53513, B2 => 
                           n51674, ZN => n59897);
   U2866 : AOI22_X1 port map( A1 => n53523, A2 => n52245, B1 => n53560, B2 => 
                           n51890, ZN => n59896);
   U2867 : AOI22_X1 port map( A1 => n53584, A2 => n52247, B1 => n53582, B2 => 
                           n51830, ZN => n59895);
   U2868 : NAND4_X1 port map( A1 => n59898, A2 => n59897, A3 => n59896, A4 => 
                           n59895, ZN => n59899);
   U2869 : AOI22_X1 port map( A1 => n60056, A2 => n59900, B1 => n60054, B2 => 
                           n59899, ZN => n59901);
   U2870 : OAI21_X1 port map( B1 => n60059, B2 => n59902, A => n59901, ZN => 
                           OUT2(7));
   U2871 : AOI22_X1 port map( A1 => n52426, A2 => n51877, B1 => n53576, B2 => 
                           n52336, ZN => n59906);
   U2872 : AOI22_X1 port map( A1 => n52421, A2 => n52084, B1 => n53568, B2 => 
                           n52385, ZN => n59905);
   U2873 : AOI22_X1 port map( A1 => n52429, A2 => n52370, B1 => n52419, B2 => 
                           n52074, ZN => n59904);
   U2874 : AOI22_X1 port map( A1 => n52432, A2 => n52373, B1 => n52424, B2 => 
                           n51873, ZN => n59903);
   U2875 : NAND4_X1 port map( A1 => n59906, A2 => n59905, A3 => n59904, A4 => 
                           n59903, ZN => n59912);
   U2876 : AOI22_X1 port map( A1 => n52428, A2 => n51884, B1 => n53585, B2 => 
                           n52122, ZN => n59910);
   U2877 : AOI22_X1 port map( A1 => n52430, A2 => n51889, B1 => n52433, B2 => 
                           n51995, ZN => n59909);
   U2878 : AOI22_X1 port map( A1 => n52422, A2 => n51872, B1 => n52431, B2 => 
                           n51982, ZN => n59908);
   U2879 : AOI22_X1 port map( A1 => n52434, A2 => n52087, B1 => n52420, B2 => 
                           n51868, ZN => n59907);
   U2880 : NAND4_X1 port map( A1 => n59910, A2 => n59909, A3 => n59908, A4 => 
                           n59907, ZN => n59911);
   U2881 : NOR2_X1 port map( A1 => n59912, A2 => n59911, ZN => n59924);
   U2882 : AOI22_X1 port map( A1 => n53579, A2 => n51935, B1 => n53560, B2 => 
                           n51912, ZN => n59916);
   U2883 : AOI22_X1 port map( A1 => n53581, A2 => n51911, B1 => n53571, B2 => 
                           n51721, ZN => n59915);
   U2884 : AOI22_X1 port map( A1 => n53516, A2 => n51950, B1 => n53520, B2 => 
                           n52342, ZN => n59914);
   U2885 : AOI22_X1 port map( A1 => n53513, A2 => n51901, B1 => n53523, B2 => 
                           n51910, ZN => n59913);
   U2886 : NAND4_X1 port map( A1 => n59916, A2 => n59915, A3 => n59914, A4 => 
                           n59913, ZN => n59922);
   U2887 : AOI22_X1 port map( A1 => n53580, A2 => n52236, B1 => n53582, B2 => 
                           n51828, ZN => n59920);
   U2888 : AOI22_X1 port map( A1 => n53562, A2 => n52078, B1 => n53560, B2 => 
                           n51878, ZN => n59919);
   U2889 : AOI22_X1 port map( A1 => n53581, A2 => n52215, B1 => n53516, B2 => 
                           n52232, ZN => n59918);
   U2890 : AOI22_X1 port map( A1 => n52400, A2 => n52235, B1 => n53571, B2 => 
                           n52204, ZN => n59917);
   U2891 : NAND4_X1 port map( A1 => n59920, A2 => n59919, A3 => n59918, A4 => 
                           n59917, ZN => n59921);
   U2892 : AOI22_X1 port map( A1 => n60056, A2 => n59922, B1 => n60054, B2 => 
                           n59921, ZN => n59923);
   U2893 : OAI21_X1 port map( B1 => n60059, B2 => n59924, A => n59923, ZN => 
                           OUT2(6));
   U2894 : AOI22_X1 port map( A1 => n52422, A2 => n51870, B1 => n53585, B2 => 
                           n52105, ZN => n59928);
   U2895 : AOI22_X1 port map( A1 => n52428, A2 => n51861, B1 => n52421, B2 => 
                           n52089, ZN => n59927);
   U2896 : AOI22_X1 port map( A1 => n52430, A2 => n51860, B1 => n52433, B2 => 
                           n51993, ZN => n59926);
   U2897 : AOI22_X1 port map( A1 => n52424, A2 => n51865, B1 => n52426, B2 => 
                           n51875, ZN => n59925);
   U2898 : NAND4_X1 port map( A1 => n59928, A2 => n59927, A3 => n59926, A4 => 
                           n59925, ZN => n59934);
   U2899 : AOI22_X1 port map( A1 => n52429, A2 => n52366, B1 => n52420, B2 => 
                           n51850, ZN => n59932);
   U2900 : AOI22_X1 port map( A1 => n52432, A2 => n52341, B1 => n52431, B2 => 
                           n51985, ZN => n59931);
   U2901 : AOI22_X1 port map( A1 => n53588, A2 => n52110, B1 => n53576, B2 => 
                           n52379, ZN => n59930);
   U2902 : AOI22_X1 port map( A1 => n52434, A2 => n52093, B1 => n53568, B2 => 
                           n52377, ZN => n59929);
   U2903 : NAND4_X1 port map( A1 => n59932, A2 => n59931, A3 => n59930, A4 => 
                           n59929, ZN => n59933);
   U2904 : NOR2_X1 port map( A1 => n59934, A2 => n59933, ZN => n59946);
   U2905 : AOI22_X1 port map( A1 => n52400, A2 => n51907, B1 => n53566, B2 => 
                           n51929, ZN => n59938);
   U2906 : AOI22_X1 port map( A1 => n53580, A2 => n51934, B1 => n53578, B2 => 
                           n51708, ZN => n59937);
   U2907 : AOI22_X1 port map( A1 => n53584, A2 => n51917, B1 => n53560, B2 => 
                           n51902, ZN => n59936);
   U2908 : AOI22_X1 port map( A1 => n53577, A2 => n51908, B1 => n53520, B2 => 
                           n52354, ZN => n59935);
   U2909 : NAND4_X1 port map( A1 => n59938, A2 => n59937, A3 => n59936, A4 => 
                           n59935, ZN => n59944);
   U2910 : AOI22_X1 port map( A1 => n53580, A2 => n52246, B1 => n53583, B2 => 
                           n52230, ZN => n59942);
   U2911 : AOI22_X1 port map( A1 => n53584, A2 => n52233, B1 => n53520, B2 => 
                           n51832, ZN => n59941);
   U2912 : AOI22_X1 port map( A1 => n53513, A2 => n52086, B1 => n53566, B2 => 
                           n52216, ZN => n59940);
   U2913 : AOI22_X1 port map( A1 => n53571, A2 => n52207, B1 => n53560, B2 => 
                           n51857, ZN => n59939);
   U2914 : NAND4_X1 port map( A1 => n59942, A2 => n59941, A3 => n59940, A4 => 
                           n59939, ZN => n59943);
   U2915 : AOI22_X1 port map( A1 => n60056, A2 => n59944, B1 => n60054, B2 => 
                           n59943, ZN => n59945);
   U2916 : OAI21_X1 port map( B1 => n60059, B2 => n59946, A => n59945, ZN => 
                           OUT2(5));
   U2917 : AOI22_X1 port map( A1 => n52421, A2 => n52119, B1 => n53568, B2 => 
                           n52374, ZN => n59950);
   U2918 : AOI22_X1 port map( A1 => n52428, A2 => n51849, B1 => n53575, B2 => 
                           n51846, ZN => n59949);
   U2919 : AOI22_X1 port map( A1 => n52431, A2 => n51986, B1 => n53588, B2 => 
                           n52077, ZN => n59948);
   U2920 : AOI22_X1 port map( A1 => n52425, A2 => n52380, B1 => n52426, B2 => 
                           n51886, ZN => n59947);
   U2921 : NAND4_X1 port map( A1 => n59950, A2 => n59949, A3 => n59948, A4 => 
                           n59947, ZN => n59956);
   U2922 : AOI22_X1 port map( A1 => n52430, A2 => n51848, B1 => n52433, B2 => 
                           n51992, ZN => n59954);
   U2923 : AOI22_X1 port map( A1 => n52432, A2 => n52375, B1 => n52429, B2 => 
                           n52378, ZN => n59953);
   U2924 : AOI22_X1 port map( A1 => n53589, A2 => n51847, B1 => n53585, B2 => 
                           n52081, ZN => n59952);
   U2925 : AOI22_X1 port map( A1 => n53586, A2 => n52114, B1 => n53564, B2 => 
                           n51869, ZN => n59951);
   U2926 : NAND4_X1 port map( A1 => n59954, A2 => n59953, A3 => n59952, A4 => 
                           n59951, ZN => n59955);
   U2927 : NOR2_X1 port map( A1 => n59956, A2 => n59955, ZN => n59968);
   U2928 : AOI22_X1 port map( A1 => n53584, A2 => n51939, B1 => n53523, B2 => 
                           n51944, ZN => n59960);
   U2929 : AOI22_X1 port map( A1 => n53582, A2 => n52308, B1 => n53560, B2 => 
                           n51949, ZN => n59959);
   U2930 : AOI22_X1 port map( A1 => n53580, A2 => n51945, B1 => n53581, B2 => 
                           n51963, ZN => n59958);
   U2931 : AOI22_X1 port map( A1 => n53514, A2 => n51732, B1 => n53577, B2 => 
                           n51959, ZN => n59957);
   U2932 : NAND4_X1 port map( A1 => n59960, A2 => n59959, A3 => n59958, A4 => 
                           n59957, ZN => n59966);
   U2933 : AOI22_X1 port map( A1 => n53579, A2 => n52250, B1 => n53523, B2 => 
                           n52239, ZN => n59964);
   U2934 : AOI22_X1 port map( A1 => n53581, A2 => n52212, B1 => n53584, B2 => 
                           n52237, ZN => n59963);
   U2935 : AOI22_X1 port map( A1 => n53577, A2 => n52102, B1 => n53571, B2 => 
                           n52202, ZN => n59962);
   U2936 : AOI22_X1 port map( A1 => n53582, A2 => n51831, B1 => n53560, B2 => 
                           n51856, ZN => n59961);
   U2937 : NAND4_X1 port map( A1 => n59964, A2 => n59963, A3 => n59962, A4 => 
                           n59961, ZN => n59965);
   U2938 : AOI22_X1 port map( A1 => n60056, A2 => n59966, B1 => n60054, B2 => 
                           n59965, ZN => n59967);
   U2939 : OAI21_X1 port map( B1 => n60059, B2 => n59968, A => n59967, ZN => 
                           OUT2(4));
   U2940 : AOI22_X1 port map( A1 => n52429, A2 => n52372, B1 => n52433, B2 => 
                           n51991, ZN => n59972);
   U2941 : AOI22_X1 port map( A1 => n52421, A2 => n52107, B1 => n53576, B2 => 
                           n52364, ZN => n59971);
   U2942 : AOI22_X1 port map( A1 => n52422, A2 => n51862, B1 => n52420, B2 => 
                           n51845, ZN => n59970);
   U2943 : AOI22_X1 port map( A1 => n52430, A2 => n51839, B1 => n52419, B2 => 
                           n52108, ZN => n59969);
   U2944 : NAND4_X1 port map( A1 => n59972, A2 => n59971, A3 => n59970, A4 => 
                           n59969, ZN => n59978);
   U2945 : AOI22_X1 port map( A1 => n53586, A2 => n52106, B1 => n52432, B2 => 
                           n52368, ZN => n59976);
   U2946 : AOI22_X1 port map( A1 => n52431, A2 => n51987, B1 => n52427, B2 => 
                           n52079, ZN => n59975);
   U2947 : AOI22_X1 port map( A1 => n52428, A2 => n51840, B1 => n52426, B2 => 
                           n51885, ZN => n59974);
   U2948 : AOI22_X1 port map( A1 => n52423, A2 => n52338, B1 => n53575, B2 => 
                           n51844, ZN => n59973);
   U2949 : NAND4_X1 port map( A1 => n59976, A2 => n59975, A3 => n59974, A4 => 
                           n59973, ZN => n59977);
   U2950 : NOR2_X1 port map( A1 => n59978, A2 => n59977, ZN => n59990);
   U2951 : AOI22_X1 port map( A1 => n53581, A2 => n51930, B1 => n53584, B2 => 
                           n51948, ZN => n59982);
   U2952 : AOI22_X1 port map( A1 => n53580, A2 => n51936, B1 => n53560, B2 => 
                           n51943, ZN => n59981);
   U2953 : AOI22_X1 port map( A1 => n53520, A2 => n52315, B1 => n53562, B2 => 
                           n51942, ZN => n59980);
   U2954 : AOI22_X1 port map( A1 => n53514, A2 => n51693, B1 => n52400, B2 => 
                           n51933, ZN => n59979);
   U2955 : NAND4_X1 port map( A1 => n59982, A2 => n59981, A3 => n59980, A4 => 
                           n59979, ZN => n59988);
   U2956 : AOI22_X1 port map( A1 => n53577, A2 => n52100, B1 => n53523, B2 => 
                           n52242, ZN => n59986);
   U2957 : AOI22_X1 port map( A1 => n53584, A2 => n52248, B1 => n53560, B2 => 
                           n51855, ZN => n59985);
   U2958 : AOI22_X1 port map( A1 => n53580, A2 => n52231, B1 => n53582, B2 => 
                           n51836, ZN => n59984);
   U2959 : AOI22_X1 port map( A1 => n53581, A2 => n52220, B1 => n53571, B2 => 
                           n52205, ZN => n59983);
   U2960 : NAND4_X1 port map( A1 => n59986, A2 => n59985, A3 => n59984, A4 => 
                           n59983, ZN => n59987);
   U2961 : AOI22_X1 port map( A1 => n60056, A2 => n59988, B1 => n60054, B2 => 
                           n59987, ZN => n59989);
   U2962 : OAI21_X1 port map( B1 => n60059, B2 => n59990, A => n59989, ZN => 
                           OUT2(3));
   U2963 : AOI22_X1 port map( A1 => n52431, A2 => n51988, B1 => n52426, B2 => 
                           n51838, ZN => n59994);
   U2964 : AOI22_X1 port map( A1 => n53575, A2 => n51883, B1 => n53576, B2 => 
                           n52363, ZN => n59993);
   U2965 : AOI22_X1 port map( A1 => n52432, A2 => n52369, B1 => n52434, B2 => 
                           n52082, ZN => n59992);
   U2966 : AOI22_X1 port map( A1 => n52421, A2 => n52075, B1 => n52419, B2 => 
                           n52103, ZN => n59991);
   U2967 : NAND4_X1 port map( A1 => n59994, A2 => n59993, A3 => n59992, A4 => 
                           n59991, ZN => n60000);
   U2968 : AOI22_X1 port map( A1 => n52428, A2 => n51879, B1 => n52427, B2 => 
                           n52116, ZN => n59998);
   U2969 : AOI22_X1 port map( A1 => n52430, A2 => n51876, B1 => n52433, B2 => 
                           n51990, ZN => n59997);
   U2970 : AOI22_X1 port map( A1 => n52429, A2 => n52376, B1 => n52420, B2 => 
                           n51882, ZN => n59996);
   U2971 : AOI22_X1 port map( A1 => n52422, A2 => n51880, B1 => n52423, B2 => 
                           n52384, ZN => n59995);
   U2972 : NAND4_X1 port map( A1 => n59998, A2 => n59997, A3 => n59996, A4 => 
                           n59995, ZN => n59999);
   U2973 : NOR2_X1 port map( A1 => n60000, A2 => n59999, ZN => n60012);
   U2974 : AOI22_X1 port map( A1 => n53579, A2 => n51941, B1 => n53516, B2 => 
                           n51947, ZN => n60004);
   U2975 : AOI22_X1 port map( A1 => n52400, A2 => n51946, B1 => n53570, B2 => 
                           n52310, ZN => n60003);
   U2976 : AOI22_X1 port map( A1 => n53514, A2 => n51762, B1 => n53581, B2 => 
                           n51955, ZN => n60002);
   U2977 : AOI22_X1 port map( A1 => n53577, A2 => n51937, B1 => n53560, B2 => 
                           n51957, ZN => n60001);
   U2978 : NAND4_X1 port map( A1 => n60004, A2 => n60003, A3 => n60002, A4 => 
                           n60001, ZN => n60010);
   U2979 : AOI22_X1 port map( A1 => n53584, A2 => n52228, B1 => n53577, B2 => 
                           n52099, ZN => n60008);
   U2980 : AOI22_X1 port map( A1 => n53571, A2 => n52210, B1 => n53570, B2 => 
                           n51835, ZN => n60007);
   U2981 : AOI22_X1 port map( A1 => n53583, A2 => n52198, B1 => n53560, B2 => 
                           n51854, ZN => n60006);
   U2982 : AOI22_X1 port map( A1 => n53580, A2 => n52199, B1 => n53581, B2 => 
                           n52218, ZN => n60005);
   U2983 : NAND4_X1 port map( A1 => n60008, A2 => n60007, A3 => n60006, A4 => 
                           n60005, ZN => n60009);
   U2984 : AOI22_X1 port map( A1 => n60056, A2 => n60010, B1 => n60054, B2 => 
                           n60009, ZN => n60011);
   U2985 : OAI21_X1 port map( B1 => n60059, B2 => n60012, A => n60011, ZN => 
                           OUT2(2));
   U2986 : AOI22_X1 port map( A1 => n52420, A2 => n51843, B1 => n53564, B2 => 
                           n51858, ZN => n60016);
   U2987 : AOI22_X1 port map( A1 => n52431, A2 => n51989, B1 => n53585, B2 => 
                           n52096, ZN => n60015);
   U2988 : AOI22_X1 port map( A1 => n52421, A2 => n52115, B1 => n52419, B2 => 
                           n52118, ZN => n60014);
   U2989 : AOI22_X1 port map( A1 => n52430, A2 => n51859, B1 => n52426, B2 => 
                           n51837, ZN => n60013);
   U2990 : NAND4_X1 port map( A1 => n60016, A2 => n60015, A3 => n60014, A4 => 
                           n60013, ZN => n60022);
   U2991 : AOI22_X1 port map( A1 => n52432, A2 => n52381, B1 => n53576, B2 => 
                           n52383, ZN => n60020);
   U2992 : AOI22_X1 port map( A1 => n52429, A2 => n52365, B1 => n52434, B2 => 
                           n52113, ZN => n60019);
   U2993 : AOI22_X1 port map( A1 => n52428, A2 => n51841, B1 => n52433, B2 => 
                           n51984, ZN => n60018);
   U2994 : AOI22_X1 port map( A1 => n52423, A2 => n52386, B1 => n52424, B2 => 
                           n51842, ZN => n60017);
   U2995 : NAND4_X1 port map( A1 => n60020, A2 => n60019, A3 => n60018, A4 => 
                           n60017, ZN => n60021);
   U2996 : NOR2_X1 port map( A1 => n60022, A2 => n60021, ZN => n60034);
   U2997 : AOI22_X1 port map( A1 => n53581, A2 => n51952, B1 => n53516, B2 => 
                           n51966, ZN => n60026);
   U2998 : AOI22_X1 port map( A1 => n53520, A2 => n52317, B1 => n53571, B2 => 
                           n51743, ZN => n60025);
   U2999 : AOI22_X1 port map( A1 => n53577, A2 => n51961, B1 => n52400, B2 => 
                           n51953, ZN => n60024);
   U3000 : AOI22_X1 port map( A1 => n53580, A2 => n51954, B1 => n53519, B2 => 
                           n51951, ZN => n60023);
   U3001 : NAND4_X1 port map( A1 => n60026, A2 => n60025, A3 => n60024, A4 => 
                           n60023, ZN => n60032);
   U3002 : AOI22_X1 port map( A1 => n53584, A2 => n52244, B1 => n53513, B2 => 
                           n52094, ZN => n60030);
   U3003 : AOI22_X1 port map( A1 => n53580, A2 => n52238, B1 => n53519, B2 => 
                           n51853, ZN => n60029);
   U3004 : AOI22_X1 port map( A1 => n53514, A2 => n52203, B1 => n53570, B2 => 
                           n51834, ZN => n60028);
   U3005 : AOI22_X1 port map( A1 => n53581, A2 => n52211, B1 => n53583, B2 => 
                           n52234, ZN => n60027);
   U3006 : NAND4_X1 port map( A1 => n60030, A2 => n60029, A3 => n60028, A4 => 
                           n60027, ZN => n60031);
   U3007 : AOI22_X1 port map( A1 => n60056, A2 => n60032, B1 => n60054, B2 => 
                           n60031, ZN => n60033);
   U3008 : OAI21_X1 port map( B1 => n60059, B2 => n60034, A => n60033, ZN => 
                           OUT2(1));
   U3009 : AOI22_X1 port map( A1 => n52430, A2 => n51688, B1 => n52426, B2 => 
                           n51684, ZN => n60038);
   U3010 : AOI22_X1 port map( A1 => n52432, A2 => n52367, B1 => n52428, B2 => 
                           n51686, ZN => n60037);
   U3011 : AOI22_X1 port map( A1 => n52422, A2 => n51689, B1 => n52425, B2 => 
                           n51681, ZN => n60036);
   U3012 : AOI22_X1 port map( A1 => n53589, A2 => n51827, B1 => n52433, B2 => 
                           n51931, ZN => n60035);
   U3013 : NAND4_X1 port map( A1 => n60038, A2 => n60037, A3 => n60036, A4 => 
                           n60035, ZN => n60044);
   U3014 : AOI22_X1 port map( A1 => n52429, A2 => n52361, B1 => n52424, B2 => 
                           n51682, ZN => n60042);
   U3015 : AOI22_X1 port map( A1 => n53585, A2 => n52227, B1 => n52419, B2 => 
                           n52120, ZN => n60041);
   U3016 : AOI22_X1 port map( A1 => n52431, A2 => n51685, B1 => n52434, B2 => 
                           n52101, ZN => n60040);
   U3017 : AOI22_X1 port map( A1 => n52421, A2 => n52229, B1 => n53568, B2 => 
                           n52285, ZN => n60039);
   U3018 : NAND4_X1 port map( A1 => n60042, A2 => n60041, A3 => n60040, A4 => 
                           n60039, ZN => n60043);
   U3019 : NOR2_X1 port map( A1 => n60044, A2 => n60043, ZN => n60058);
   U3020 : AOI22_X1 port map( A1 => n53583, A2 => n51973, B1 => n53578, B2 => 
                           n51683, ZN => n60048);
   U3021 : AOI22_X1 port map( A1 => n53580, A2 => n51977, B1 => n53581, B2 => 
                           n51932, ZN => n60047);
   U3022 : AOI22_X1 port map( A1 => n53582, A2 => n52335, B1 => n53577, B2 => 
                           n51980, ZN => n60046);
   U3023 : AOI22_X1 port map( A1 => n53519, A2 => n51979, B1 => n53584, B2 => 
                           n51975, ZN => n60045);
   U3024 : NAND4_X1 port map( A1 => n60048, A2 => n60047, A3 => n60046, A4 => 
                           n60045, ZN => n60055);
   U3025 : AOI22_X1 port map( A1 => n53515, A2 => n52158, B1 => n53523, B2 => 
                           n52166, ZN => n60052);
   U3026 : AOI22_X1 port map( A1 => n53519, A2 => n51690, B1 => n53578, B2 => 
                           n52226, ZN => n60051);
   U3027 : AOI22_X1 port map( A1 => n53512, A2 => n52167, B1 => n53565, B2 => 
                           n52165, ZN => n60050);
   U3028 : AOI22_X1 port map( A1 => n53582, A2 => n51687, B1 => n53513, B2 => 
                           n52097, ZN => n60049);
   U3029 : NAND4_X1 port map( A1 => n60052, A2 => n60051, A3 => n60050, A4 => 
                           n60049, ZN => n60053);
   U3030 : AOI22_X1 port map( A1 => n60056, A2 => n60055, B1 => n60054, B2 => 
                           n60053, ZN => n60057);
   U3031 : OAI21_X1 port map( B1 => n60059, B2 => n60058, A => n60057, ZN => 
                           OUT2(0));
   U3032 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n60063)
                           ;
   U3033 : NOR2_X1 port map( A1 => n3562, A2 => n60063, ZN => n40587);
   U3034 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n3558, ZN => n60062);
   U3035 : INV_X1 port map( A => n3566, ZN => n60060);
   U3036 : NOR2_X1 port map( A1 => n60062, A2 => n60060, ZN => n40586);
   U3037 : NOR2_X1 port map( A1 => n3562, A2 => n60062, ZN => n40585);
   U3038 : NOR2_X1 port map( A1 => n60063, A2 => n3564, ZN => n40584);
   U3039 : NOR2_X1 port map( A1 => n60062, A2 => n3559, ZN => n40583);
   U3040 : NOR2_X1 port map( A1 => n60062, A2 => n3561, ZN => n40582);
   U3041 : NOR2_X1 port map( A1 => n60062, A2 => n3563, ZN => n40581);
   U3042 : NOR2_X1 port map( A1 => n60062, A2 => n3564, ZN => n40580);
   U3043 : NOR2_X1 port map( A1 => n60063, A2 => n60060, ZN => n49095);
   U3044 : NOR2_X1 port map( A1 => n60063, A2 => n3561, ZN => n47430);
   U3045 : INV_X1 port map( A => n3560, ZN => n60061);
   U3046 : NOR2_X1 port map( A1 => n60062, A2 => n60061, ZN => n40577);
   U3047 : NOR2_X1 port map( A1 => n60063, A2 => n60061, ZN => n40576);
   U3048 : NOR2_X1 port map( A1 => n60062, A2 => n3565, ZN => n49096);
   U3049 : NOR2_X1 port map( A1 => n60063, A2 => n3563, ZN => n40574);
   U3050 : NOR2_X1 port map( A1 => n60063, A2 => n3559, ZN => n49097);
   U3051 : NOR2_X1 port map( A1 => n60063, A2 => n3565, ZN => n47431);
   U3052 : AOI22_X1 port map( A1 => n51390, A2 => n52418, B1 => n51371, B2 => 
                           n53555, ZN => n60067);
   U3053 : AOI22_X1 port map( A1 => n51555, A2 => n52417, B1 => n51409, B2 => 
                           n53553, ZN => n60066);
   U3054 : AOI22_X1 port map( A1 => n51548, A2 => n53557, B1 => n51370, B2 => 
                           n52411, ZN => n60065);
   U3055 : AOI22_X1 port map( A1 => n51645, A2 => n52404, B1 => n51511, B2 => 
                           n52409, ZN => n60064);
   U3056 : NAND4_X1 port map( A1 => n60067, A2 => n60066, A3 => n60065, A4 => 
                           n60064, ZN => n60073);
   U3057 : AOI22_X1 port map( A1 => n51580, A2 => n52415, B1 => n51627, B2 => 
                           n53554, ZN => n60071);
   U3058 : AOI22_X1 port map( A1 => n51493, A2 => n53556, B1 => n51604, B2 => 
                           n52410, ZN => n60070);
   U3059 : AOI22_X1 port map( A1 => n51387, A2 => n52414, B1 => n51557, B2 => 
                           n52406, ZN => n60069);
   U3060 : AOI22_X1 port map( A1 => n51389, A2 => n53552, B1 => n51556, B2 => 
                           n53558, ZN => n60068);
   U3061 : NAND4_X1 port map( A1 => n60071, A2 => n60070, A3 => n60069, A4 => 
                           n60068, ZN => n60072);
   U3062 : NOR2_X1 port map( A1 => n60073, A2 => n60072, ZN => n60085);
   U3063 : NOR3_X1 port map( A1 => n53624, A2 => n53625, A3 => n60727, ZN => 
                           n60525);
   U3064 : CLKBUF_X1 port map( A => n60525, Z => n60570);
   U3065 : AOI22_X1 port map( A1 => n51470, A2 => n53549, B1 => n51455, B2 => 
                           n53526, ZN => n60077);
   U3066 : AOI22_X1 port map( A1 => n51465, A2 => n53527, B1 => n51405, B2 => 
                           n53551, ZN => n60076);
   U3067 : AOI22_X1 port map( A1 => n51478, A2 => n52402, B1 => n51668, B2 => 
                           n53550, ZN => n60075);
   U3068 : AOI22_X1 port map( A1 => n51452, A2 => n53517, B1 => n51464, B2 => 
                           n52401, ZN => n60074);
   U3069 : NAND4_X1 port map( A1 => n60077, A2 => n60076, A3 => n60075, A4 => 
                           n60074, ZN => n60083);
   U3070 : NOR3_X1 port map( A1 => n53625, A2 => n52483, A3 => n60727, ZN => 
                           n60303);
   U3071 : AOI22_X1 port map( A1 => n51394, A2 => n53547, B1 => n51570, B2 => 
                           n53551, ZN => n60081);
   U3072 : AOI22_X1 port map( A1 => n51617, A2 => n53546, B1 => n51583, B2 => 
                           n53525, ZN => n60080);
   U3073 : AOI22_X1 port map( A1 => n51566, A2 => n52482, B1 => n51395, B2 => 
                           n53550, ZN => n60079);
   U3074 : AOI22_X1 port map( A1 => n51565, A2 => n52481, B1 => n51596, B2 => 
                           n53527, ZN => n60078);
   U3075 : NAND4_X1 port map( A1 => n60081, A2 => n60080, A3 => n60079, A4 => 
                           n60078, ZN => n60082);
   U3076 : AOI22_X1 port map( A1 => n60570, A2 => n60083, B1 => n60303, B2 => 
                           n60082, ZN => n60084);
   U3077 : OAI21_X1 port map( B1 => n60727, B2 => n60085, A => n60084, ZN => 
                           OUT1(31));
   U3078 : AOI22_X1 port map( A1 => n51372, A2 => n52411, B1 => n51519, B2 => 
                           n52412, ZN => n60089);
   U3079 : AOI22_X1 port map( A1 => n51382, A2 => n52418, B1 => n51624, B2 => 
                           n53544, ZN => n60088);
   U3080 : AOI22_X1 port map( A1 => n51538, A2 => n53543, B1 => n51420, B2 => 
                           n52403, ZN => n60087);
   U3081 : AOI22_X1 port map( A1 => n51421, A2 => n52416, B1 => n51680, B2 => 
                           n53542, ZN => n60086);
   U3082 : NAND4_X1 port map( A1 => n60089, A2 => n60088, A3 => n60087, A4 => 
                           n60086, ZN => n60095);
   U3083 : AOI22_X1 port map( A1 => n51644, A2 => n52405, B1 => n51522, B2 => 
                           n52413, ZN => n60093);
   U3084 : AOI22_X1 port map( A1 => n51446, A2 => n52409, B1 => n51414, B2 => 
                           n52414, ZN => n60092);
   U3085 : AOI22_X1 port map( A1 => n51535, A2 => n52406, B1 => n51462, B2 => 
                           n52407, ZN => n60091);
   U3086 : AOI22_X1 port map( A1 => n51650, A2 => n53545, B1 => n51413, B2 => 
                           n53552, ZN => n60090);
   U3087 : NAND4_X1 port map( A1 => n60093, A2 => n60092, A3 => n60091, A4 => 
                           n60090, ZN => n60094);
   U3088 : NOR2_X1 port map( A1 => n60095, A2 => n60094, ZN => n60107);
   U3089 : AOI22_X1 port map( A1 => n51463, A2 => n52401, B1 => n51461, B2 => 
                           n52479, ZN => n60099);
   U3090 : AOI22_X1 port map( A1 => n51444, A2 => n53524, B1 => n51381, B2 => 
                           n53522, ZN => n60098);
   U3091 : AOI22_X1 port map( A1 => n51441, A2 => n53547, B1 => n51436, B2 => 
                           n53525, ZN => n60097);
   U3092 : AOI22_X1 port map( A1 => n51496, A2 => n53526, B1 => n51540, B2 => 
                           n53518, ZN => n60096);
   U3093 : NAND4_X1 port map( A1 => n60099, A2 => n60098, A3 => n60097, A4 => 
                           n60096, ZN => n60105);
   U3094 : CLKBUF_X1 port map( A => n60303, Z => n60769);
   U3095 : AOI22_X1 port map( A1 => n51629, A2 => n53525, B1 => n51677, B2 => 
                           n53522, ZN => n60103);
   U3096 : AOI22_X1 port map( A1 => n51407, A2 => n53518, B1 => n51564, B2 => 
                           n53540, ZN => n60102);
   U3097 : AOI22_X1 port map( A1 => n51633, A2 => n53541, B1 => n51614, B2 => 
                           n53524, ZN => n60101);
   U3098 : AOI22_X1 port map( A1 => n51411, A2 => n53517, B1 => n51639, B2 => 
                           n53546, ZN => n60100);
   U3099 : NAND4_X1 port map( A1 => n60103, A2 => n60102, A3 => n60101, A4 => 
                           n60100, ZN => n60104);
   U3100 : AOI22_X1 port map( A1 => n60570, A2 => n60105, B1 => n60769, B2 => 
                           n60104, ZN => n60106);
   U3101 : OAI21_X1 port map( B1 => n60727, B2 => n60107, A => n60106, ZN => 
                           OUT1(30));
   U3102 : AOI22_X1 port map( A1 => n51658, A2 => n52410, B1 => n51472, B2 => 
                           n53556, ZN => n60111);
   U3103 : AOI22_X1 port map( A1 => n51431, A2 => n52414, B1 => n51432, B2 => 
                           n53555, ZN => n60110);
   U3104 : AOI22_X1 port map( A1 => n51424, A2 => n53552, B1 => n51523, B2 => 
                           n52412, ZN => n60109);
   U3105 : AOI22_X1 port map( A1 => n51518, A2 => n53557, B1 => n51648, B2 => 
                           n52415, ZN => n60108);
   U3106 : NAND4_X1 port map( A1 => n60111, A2 => n60110, A3 => n60109, A4 => 
                           n60108, ZN => n60117);
   U3107 : AOI22_X1 port map( A1 => n51434, A2 => n52418, B1 => n51657, B2 => 
                           n52405, ZN => n60115);
   U3108 : AOI22_X1 port map( A1 => n51486, A2 => n52409, B1 => n51517, B2 => 
                           n52417, ZN => n60114);
   U3109 : AOI22_X1 port map( A1 => n51366, A2 => n52411, B1 => n51433, B2 => 
                           n53553, ZN => n60113);
   U3110 : AOI22_X1 port map( A1 => n51524, A2 => n52406, B1 => n51568, B2 => 
                           n52404, ZN => n60112);
   U3111 : NAND4_X1 port map( A1 => n60115, A2 => n60114, A3 => n60113, A4 => 
                           n60112, ZN => n60116);
   U3112 : NOR2_X1 port map( A1 => n60117, A2 => n60116, ZN => n60129);
   U3113 : AOI22_X1 port map( A1 => n51577, A2 => n53518, B1 => n51497, B2 => 
                           n52481, ZN => n60121);
   U3114 : AOI22_X1 port map( A1 => n51492, A2 => n53517, B1 => n51490, B2 => 
                           n53549, ZN => n60120);
   U3115 : AOI22_X1 port map( A1 => n51392, A2 => n53551, B1 => n51460, B2 => 
                           n52402, ZN => n60119);
   U3116 : AOI22_X1 port map( A1 => n51489, A2 => n52401, B1 => n51459, B2 => 
                           n53527, ZN => n60118);
   U3117 : NAND4_X1 port map( A1 => n60121, A2 => n60120, A3 => n60119, A4 => 
                           n60118, ZN => n60127);
   U3118 : AOI22_X1 port map( A1 => n51587, A2 => n53539, B1 => n51594, B2 => 
                           n53541, ZN => n60125);
   U3119 : AOI22_X1 port map( A1 => n51406, A2 => n53518, B1 => n51606, B2 => 
                           n52482, ZN => n60124);
   U3120 : AOI22_X1 port map( A1 => n51563, A2 => n53540, B1 => n51400, B2 => 
                           n53548, ZN => n60123);
   U3121 : AOI22_X1 port map( A1 => n51588, A2 => n53528, B1 => n51534, B2 => 
                           n53522, ZN => n60122);
   U3122 : NAND4_X1 port map( A1 => n60125, A2 => n60124, A3 => n60123, A4 => 
                           n60122, ZN => n60126);
   U3123 : AOI22_X1 port map( A1 => n60570, A2 => n60127, B1 => n60303, B2 => 
                           n60126, ZN => n60128);
   U3124 : OAI21_X1 port map( B1 => n60727, B2 => n60129, A => n60128, ZN => 
                           OUT1(29));
   U3125 : AOI22_X1 port map( A1 => n51426, A2 => n52403, B1 => n51643, B2 => 
                           n52405, ZN => n60133);
   U3126 : AOI22_X1 port map( A1 => n51672, A2 => n52415, B1 => n51628, B2 => 
                           n53544, ZN => n60132);
   U3127 : AOI22_X1 port map( A1 => n51448, A2 => n53556, B1 => n51368, B2 => 
                           n52411, ZN => n60131);
   U3128 : AOI22_X1 port map( A1 => n51419, A2 => n52414, B1 => n51549, B2 => 
                           n52406, ZN => n60130);
   U3129 : NAND4_X1 port map( A1 => n60133, A2 => n60132, A3 => n60131, A4 => 
                           n60130, ZN => n60139);
   U3130 : AOI22_X1 port map( A1 => n51418, A2 => n52416, B1 => n51373, B2 => 
                           n52418, ZN => n60137);
   U3131 : AOI22_X1 port map( A1 => n51454, A2 => n52409, B1 => n51415, B2 => 
                           n52408, ZN => n60136);
   U3132 : AOI22_X1 port map( A1 => n51651, A2 => n53545, B1 => n51675, B2 => 
                           n52417, ZN => n60135);
   U3133 : AOI22_X1 port map( A1 => n51550, A2 => n52412, B1 => n51571, B2 => 
                           n52413, ZN => n60134);
   U3134 : NAND4_X1 port map( A1 => n60137, A2 => n60136, A3 => n60135, A4 => 
                           n60134, ZN => n60138);
   U3135 : NOR2_X1 port map( A1 => n60139, A2 => n60138, ZN => n60151);
   U3136 : AOI22_X1 port map( A1 => n51450, A2 => n53541, B1 => n51379, B2 => 
                           n52480, ZN => n60143);
   U3137 : AOI22_X1 port map( A1 => n51505, A2 => n52401, B1 => n51671, B2 => 
                           n53538, ZN => n60142);
   U3138 : AOI22_X1 port map( A1 => n51442, A2 => n53525, B1 => n51506, B2 => 
                           n53549, ZN => n60141);
   U3139 : AOI22_X1 port map( A1 => n51503, A2 => n53548, B1 => n51447, B2 => 
                           n52481, ZN => n60140);
   U3140 : NAND4_X1 port map( A1 => n60143, A2 => n60142, A3 => n60141, A4 => 
                           n60140, ZN => n60149);
   U3141 : AOI22_X1 port map( A1 => n51634, A2 => n52479, B1 => n51647, B2 => 
                           n53525, ZN => n60147);
   U3142 : AOI22_X1 port map( A1 => n51640, A2 => n53546, B1 => n51404, B2 => 
                           n53518, ZN => n60146);
   U3143 : AOI22_X1 port map( A1 => n51428, A2 => n53548, B1 => n51673, B2 => 
                           n53522, ZN => n60145);
   U3144 : AOI22_X1 port map( A1 => n51597, A2 => n53524, B1 => n51561, B2 => 
                           n53540, ZN => n60144);
   U3145 : NAND4_X1 port map( A1 => n60147, A2 => n60146, A3 => n60145, A4 => 
                           n60144, ZN => n60148);
   U3146 : AOI22_X1 port map( A1 => n60570, A2 => n60149, B1 => n60769, B2 => 
                           n60148, ZN => n60150);
   U3147 : OAI21_X1 port map( B1 => n60727, B2 => n60151, A => n60150, ZN => 
                           OUT1(28));
   U3148 : AOI22_X1 port map( A1 => n51642, A2 => n52405, B1 => n51410, B2 => 
                           n52408, ZN => n60155);
   U3149 : AOI22_X1 port map( A1 => n51416, A2 => n52403, B1 => n51529, B2 => 
                           n52404, ZN => n60154);
   U3150 : AOI22_X1 port map( A1 => n51653, A2 => n52410, B1 => n51423, B2 => 
                           n52414, ZN => n60153);
   U3151 : AOI22_X1 port map( A1 => n51422, A2 => n52416, B1 => n51679, B2 => 
                           n53542, ZN => n60152);
   U3152 : NAND4_X1 port map( A1 => n60155, A2 => n60154, A3 => n60153, A4 => 
                           n60152, ZN => n60161);
   U3153 : AOI22_X1 port map( A1 => n51676, A2 => n52415, B1 => n51377, B2 => 
                           n53536, ZN => n60159);
   U3154 : AOI22_X1 port map( A1 => n51536, A2 => n53558, B1 => n51525, B2 => 
                           n53557, ZN => n60158);
   U3155 : AOI22_X1 port map( A1 => n51528, A2 => n53535, B1 => n51453, B2 => 
                           n52407, ZN => n60157);
   U3156 : AOI22_X1 port map( A1 => n51438, A2 => n53534, B1 => n51385, B2 => 
                           n53537, ZN => n60156);
   U3157 : NAND4_X1 port map( A1 => n60159, A2 => n60158, A3 => n60157, A4 => 
                           n60156, ZN => n60160);
   U3158 : NOR2_X1 port map( A1 => n60161, A2 => n60160, ZN => n60173);
   U3159 : AOI22_X1 port map( A1 => n51479, A2 => n53548, B1 => n51439, B2 => 
                           n53541, ZN => n60165);
   U3160 : AOI22_X1 port map( A1 => n51451, A2 => n53539, B1 => n51365, B2 => 
                           n53522, ZN => n60164);
   U3161 : AOI22_X1 port map( A1 => n51469, A2 => n53549, B1 => n51474, B2 => 
                           n52401, ZN => n60163);
   U3162 : AOI22_X1 port map( A1 => n51494, A2 => n52481, B1 => n51663, B2 => 
                           n53518, ZN => n60162);
   U3163 : NAND4_X1 port map( A1 => n60165, A2 => n60164, A3 => n60163, A4 => 
                           n60162, ZN => n60171);
   U3164 : AOI22_X1 port map( A1 => n51641, A2 => n53546, B1 => n51635, B2 => 
                           n53541, ZN => n60169);
   U3165 : AOI22_X1 port map( A1 => n51402, A2 => n53538, B1 => n51661, B2 => 
                           n53551, ZN => n60168);
   U3166 : AOI22_X1 port map( A1 => n51559, A2 => n53526, B1 => n51630, B2 => 
                           n52402, ZN => n60167);
   U3167 : AOI22_X1 port map( A1 => n51417, A2 => n53547, B1 => n51613, B2 => 
                           n53549, ZN => n60166);
   U3168 : NAND4_X1 port map( A1 => n60169, A2 => n60168, A3 => n60167, A4 => 
                           n60166, ZN => n60170);
   U3169 : AOI22_X1 port map( A1 => n60570, A2 => n60171, B1 => n60303, B2 => 
                           n60170, ZN => n60172);
   U3170 : OAI21_X1 port map( B1 => n60727, B2 => n60173, A => n60172, ZN => 
                           OUT1(27));
   U3171 : AOI22_X1 port map( A1 => n51542, A2 => n52413, B1 => n51388, B2 => 
                           n52416, ZN => n60177);
   U3172 : AOI22_X1 port map( A1 => n51430, A2 => n52403, B1 => n51399, B2 => 
                           n53536, ZN => n60176);
   U3173 : AOI22_X1 port map( A1 => n51567, A2 => n53535, B1 => n51429, B2 => 
                           n52418, ZN => n60175);
   U3174 : AOI22_X1 port map( A1 => n51649, A2 => n52415, B1 => n51425, B2 => 
                           n52414, ZN => n60174);
   U3175 : NAND4_X1 port map( A1 => n60177, A2 => n60176, A3 => n60175, A4 => 
                           n60174, ZN => n60183);
   U3176 : AOI22_X1 port map( A1 => n51485, A2 => n52409, B1 => n51491, B2 => 
                           n52407, ZN => n60181);
   U3177 : AOI22_X1 port map( A1 => n51551, A2 => n53558, B1 => n51531, B2 => 
                           n52404, ZN => n60180);
   U3178 : AOI22_X1 port map( A1 => n51427, A2 => n52408, B1 => n51660, B2 => 
                           n52405, ZN => n60179);
   U3179 : AOI22_X1 port map( A1 => n51655, A2 => n53544, B1 => n51547, B2 => 
                           n52417, ZN => n60178);
   U3180 : NAND4_X1 port map( A1 => n60181, A2 => n60180, A3 => n60179, A4 => 
                           n60178, ZN => n60182);
   U3181 : NOR2_X1 port map( A1 => n60183, A2 => n60182, ZN => n60195);
   U3182 : AOI22_X1 port map( A1 => n51458, A2 => n53525, B1 => n51467, B2 => 
                           n53528, ZN => n60187);
   U3183 : AOI22_X1 port map( A1 => n51475, A2 => n53527, B1 => n51488, B2 => 
                           n53526, ZN => n60186);
   U3184 : AOI22_X1 port map( A1 => n51466, A2 => n53549, B1 => n51589, B2 => 
                           n53538, ZN => n60185);
   U3185 : AOI22_X1 port map( A1 => n51383, A2 => n53551, B1 => n51457, B2 => 
                           n53548, ZN => n60184);
   U3186 : NAND4_X1 port map( A1 => n60187, A2 => n60186, A3 => n60185, A4 => 
                           n60184, ZN => n60193);
   U3187 : AOI22_X1 port map( A1 => n51403, A2 => n53548, B1 => n51572, B2 => 
                           n52480, ZN => n60191);
   U3188 : AOI22_X1 port map( A1 => n51546, A2 => n53526, B1 => n51610, B2 => 
                           n52401, ZN => n60190);
   U3189 : AOI22_X1 port map( A1 => n51612, A2 => n53527, B1 => n51401, B2 => 
                           n53538, ZN => n60189);
   U3190 : AOI22_X1 port map( A1 => n51591, A2 => n53539, B1 => n51598, B2 => 
                           n52482, ZN => n60188);
   U3191 : NAND4_X1 port map( A1 => n60191, A2 => n60190, A3 => n60189, A4 => 
                           n60188, ZN => n60192);
   U3192 : AOI22_X1 port map( A1 => n60570, A2 => n60193, B1 => n60769, B2 => 
                           n60192, ZN => n60194);
   U3193 : OAI21_X1 port map( B1 => n60727, B2 => n60195, A => n60194, ZN => 
                           OUT1(26));
   U3194 : AOI22_X1 port map( A1 => n51437, A2 => n53556, B1 => n51374, B2 => 
                           n53537, ZN => n60199);
   U3195 : AOI22_X1 port map( A1 => n51397, A2 => n53552, B1 => n51375, B2 => 
                           n53555, ZN => n60198);
   U3196 : AOI22_X1 port map( A1 => n51665, A2 => n52417, B1 => n51393, B2 => 
                           n52403, ZN => n60197);
   U3197 : AOI22_X1 port map( A1 => n51574, A2 => n52412, B1 => n51468, B2 => 
                           n53534, ZN => n60196);
   U3198 : NAND4_X1 port map( A1 => n60199, A2 => n60198, A3 => n60197, A4 => 
                           n60196, ZN => n60205);
   U3199 : AOI22_X1 port map( A1 => n51569, A2 => n53557, B1 => n51618, B2 => 
                           n52410, ZN => n60203);
   U3200 : AOI22_X1 port map( A1 => n51664, A2 => n53543, B1 => n51376, B2 => 
                           n53536, ZN => n60202);
   U3201 : AOI22_X1 port map( A1 => n51652, A2 => n53545, B1 => n51637, B2 => 
                           n53554, ZN => n60201);
   U3202 : AOI22_X1 port map( A1 => n51398, A2 => n53533, B1 => n51573, B2 => 
                           n52406, ZN => n60200);
   U3203 : NAND4_X1 port map( A1 => n60203, A2 => n60202, A3 => n60201, A4 => 
                           n60200, ZN => n60204);
   U3204 : NOR2_X1 port map( A1 => n60205, A2 => n60204, ZN => n60217);
   U3205 : AOI22_X1 port map( A1 => n51440, A2 => n53527, B1 => n51502, B2 => 
                           n53546, ZN => n60209);
   U3206 : AOI22_X1 port map( A1 => n51666, A2 => n53550, B1 => n51471, B2 => 
                           n52481, ZN => n60208);
   U3207 : AOI22_X1 port map( A1 => n51456, A2 => n53525, B1 => n51487, B2 => 
                           n52482, ZN => n60207);
   U3208 : AOI22_X1 port map( A1 => n51477, A2 => n53547, B1 => n51364, B2 => 
                           n53522, ZN => n60206);
   U3209 : NAND4_X1 port map( A1 => n60209, A2 => n60208, A3 => n60207, A4 => 
                           n60206, ZN => n60215);
   U3210 : AOI22_X1 port map( A1 => n51631, A2 => n52402, B1 => n51646, B2 => 
                           n52401, ZN => n60213);
   U3211 : AOI22_X1 port map( A1 => n51636, A2 => n52479, B1 => n51412, B2 => 
                           n53547, ZN => n60212);
   U3212 : AOI22_X1 port map( A1 => n51386, A2 => n53550, B1 => n51678, B2 => 
                           n53522, ZN => n60211);
   U3213 : AOI22_X1 port map( A1 => n51576, A2 => n53540, B1 => n51605, B2 => 
                           n53524, ZN => n60210);
   U3214 : NAND4_X1 port map( A1 => n60213, A2 => n60212, A3 => n60211, A4 => 
                           n60210, ZN => n60214);
   U3215 : AOI22_X1 port map( A1 => n60570, A2 => n60215, B1 => n60769, B2 => 
                           n60214, ZN => n60216);
   U3216 : OAI21_X1 port map( B1 => n60727, B2 => n60217, A => n60216, ZN => 
                           OUT1(25));
   U3217 : AOI22_X1 port map( A1 => n51530, A2 => n52417, B1 => n51367, B2 => 
                           n53537, ZN => n60221);
   U3218 : AOI22_X1 port map( A1 => n51558, A2 => n53543, B1 => n51369, B2 => 
                           n52414, ZN => n60220);
   U3219 : AOI22_X1 port map( A1 => n51396, A2 => n52416, B1 => n51408, B2 => 
                           n53536, ZN => n60219);
   U3220 : AOI22_X1 port map( A1 => n51662, A2 => n52405, B1 => n51593, B2 => 
                           n52412, ZN => n60218);
   U3221 : NAND4_X1 port map( A1 => n60221, A2 => n60220, A3 => n60219, A4 => 
                           n60218, ZN => n60227);
   U3222 : AOI22_X1 port map( A1 => n51595, A2 => n52413, B1 => n51378, B2 => 
                           n53553, ZN => n60225);
   U3223 : AOI22_X1 port map( A1 => n51625, A2 => n52406, B1 => n51443, B2 => 
                           n52407, ZN => n60224);
   U3224 : AOI22_X1 port map( A1 => n51543, A2 => n52404, B1 => n51391, B2 => 
                           n53552, ZN => n60223);
   U3225 : AOI22_X1 port map( A1 => n51484, A2 => n53534, B1 => n51654, B2 => 
                           n53544, ZN => n60222);
   U3226 : NAND4_X1 port map( A1 => n60225, A2 => n60224, A3 => n60223, A4 => 
                           n60222, ZN => n60226);
   U3227 : NOR2_X1 port map( A1 => n60227, A2 => n60226, ZN => n60239);
   U3228 : AOI22_X1 port map( A1 => n51435, A2 => n53551, B1 => n51507, B2 => 
                           n53524, ZN => n60231);
   U3229 : AOI22_X1 port map( A1 => n51473, A2 => n53539, B1 => n51501, B2 => 
                           n53540, ZN => n60230);
   U3230 : AOI22_X1 port map( A1 => n51554, A2 => n53550, B1 => n51504, B2 => 
                           n53528, ZN => n60229);
   U3231 : AOI22_X1 port map( A1 => n51499, A2 => n53547, B1 => n51515, B2 => 
                           n52479, ZN => n60228);
   U3232 : NAND4_X1 port map( A1 => n60231, A2 => n60230, A3 => n60229, A4 => 
                           n60228, ZN => n60237);
   U3233 : AOI22_X1 port map( A1 => n51584, A2 => n53541, B1 => n51620, B2 => 
                           n53522, ZN => n60235);
   U3234 : AOI22_X1 port map( A1 => n51600, A2 => n52482, B1 => n51609, B2 => 
                           n53546, ZN => n60234);
   U3235 : AOI22_X1 port map( A1 => n51603, A2 => n53525, B1 => n51380, B2 => 
                           n53547, ZN => n60233);
   U3236 : AOI22_X1 port map( A1 => n51622, A2 => n53526, B1 => n51384, B2 => 
                           n53550, ZN => n60232);
   U3237 : NAND4_X1 port map( A1 => n60235, A2 => n60234, A3 => n60233, A4 => 
                           n60232, ZN => n60236);
   U3238 : AOI22_X1 port map( A1 => n60570, A2 => n60237, B1 => n60303, B2 => 
                           n60236, ZN => n60238);
   U3239 : OAI21_X1 port map( B1 => n60727, B2 => n60239, A => n60238, ZN => 
                           OUT1(24));
   U3240 : AOI22_X1 port map( A1 => n52161, A2 => n52404, B1 => n51906, B2 => 
                           n52407, ZN => n60243);
   U3241 : AOI22_X1 port map( A1 => n52141, A2 => n52412, B1 => n51723, B2 => 
                           n53537, ZN => n60242);
   U3242 : AOI22_X1 port map( A1 => n52265, A2 => n53535, B1 => n51709, B2 => 
                           n52403, ZN => n60241);
   U3243 : AOI22_X1 port map( A1 => n51699, A2 => n53533, B1 => n51623, B2 => 
                           n53544, ZN => n60240);
   U3244 : NAND4_X1 port map( A1 => n60243, A2 => n60242, A3 => n60241, A4 => 
                           n60240, ZN => n60249);
   U3245 : AOI22_X1 port map( A1 => n51756, A2 => n53552, B1 => n52142, B2 => 
                           n53542, ZN => n60247);
   U3246 : AOI22_X1 port map( A1 => n51777, A2 => n52416, B1 => n51923, B2 => 
                           n53534, ZN => n60246);
   U3247 : AOI22_X1 port map( A1 => n51521, A2 => n52413, B1 => n52182, B2 => 
                           n53554, ZN => n60245);
   U3248 : AOI22_X1 port map( A1 => n51638, A2 => n52415, B1 => n51817, B2 => 
                           n52411, ZN => n60244);
   U3249 : NAND4_X1 port map( A1 => n60247, A2 => n60246, A3 => n60245, A4 => 
                           n60244, ZN => n60248);
   U3250 : NOR2_X1 port map( A1 => n60249, A2 => n60248, ZN => n60261);
   U3251 : AOI22_X1 port map( A1 => n51900, A2 => n53549, B1 => n52011, B2 => 
                           n53547, ZN => n60253);
   U3252 : AOI22_X1 port map( A1 => n51481, A2 => n52402, B1 => n51940, B2 => 
                           n52401, ZN => n60252);
   U3253 : AOI22_X1 port map( A1 => n51864, A2 => n52480, B1 => n52138, B2 => 
                           n53550, ZN => n60251);
   U3254 : AOI22_X1 port map( A1 => n51498, A2 => n52481, B1 => n51480, B2 => 
                           n52479, ZN => n60250);
   U3255 : NAND4_X1 port map( A1 => n60253, A2 => n60252, A3 => n60251, A4 => 
                           n60250, ZN => n60259);
   U3256 : AOI22_X1 port map( A1 => n51867, A2 => n53550, B1 => n52176, B2 => 
                           n53546, ZN => n60257);
   U3257 : AOI22_X1 port map( A1 => n52178, A2 => n52479, B1 => n52267, B2 => 
                           n53526, ZN => n60256);
   U3258 : AOI22_X1 port map( A1 => n51692, A2 => n53548, B1 => n52149, B2 => 
                           n52482, ZN => n60255);
   U3259 : AOI22_X1 port map( A1 => n52140, A2 => n53522, B1 => n52180, B2 => 
                           n52402, ZN => n60254);
   U3260 : NAND4_X1 port map( A1 => n60257, A2 => n60256, A3 => n60255, A4 => 
                           n60254, ZN => n60258);
   U3261 : AOI22_X1 port map( A1 => n60570, A2 => n60259, B1 => n60303, B2 => 
                           n60258, ZN => n60260);
   U3262 : OAI21_X1 port map( B1 => n60774, B2 => n60261, A => n60260, ZN => 
                           OUT1(23));
   U3263 : AOI22_X1 port map( A1 => n52127, A2 => n52413, B1 => n52172, B2 => 
                           n53543, ZN => n60265);
   U3264 : AOI22_X1 port map( A1 => n51704, A2 => n53533, B1 => n52139, B2 => 
                           n52417, ZN => n60264);
   U3265 : AOI22_X1 port map( A1 => n51445, A2 => n52407, B1 => n51694, B2 => 
                           n53555, ZN => n60263);
   U3266 : AOI22_X1 port map( A1 => n52181, A2 => n53554, B1 => n51818, B2 => 
                           n53536, ZN => n60262);
   U3267 : NAND4_X1 port map( A1 => n60265, A2 => n60264, A3 => n60263, A4 => 
                           n60262, ZN => n60271);
   U3268 : AOI22_X1 port map( A1 => n52136, A2 => n53558, B1 => n51707, B2 => 
                           n53553, ZN => n60269);
   U3269 : AOI22_X1 port map( A1 => n51760, A2 => n53552, B1 => n51903, B2 => 
                           n53534, ZN => n60268);
   U3270 : AOI22_X1 port map( A1 => n52174, A2 => n53544, B1 => n52264, B2 => 
                           n53535, ZN => n60267);
   U3271 : AOI22_X1 port map( A1 => n52171, A2 => n52404, B1 => n51722, B2 => 
                           n52418, ZN => n60266);
   U3272 : NAND4_X1 port map( A1 => n60269, A2 => n60268, A3 => n60267, A4 => 
                           n60266, ZN => n60270);
   U3273 : NOR2_X1 port map( A1 => n60271, A2 => n60270, ZN => n60283);
   U3274 : AOI22_X1 port map( A1 => n52137, A2 => n53550, B1 => n51958, B2 => 
                           n53539, ZN => n60275);
   U3275 : AOI22_X1 port map( A1 => n51495, A2 => n52401, B1 => n52010, B2 => 
                           n53540, ZN => n60274);
   U3276 : AOI22_X1 port map( A1 => n52002, A2 => n53541, B1 => n51500, B2 => 
                           n53547, ZN => n60273);
   U3277 : AOI22_X1 port map( A1 => n51866, A2 => n53551, B1 => n52007, B2 => 
                           n53549, ZN => n60272);
   U3278 : NAND4_X1 port map( A1 => n60275, A2 => n60274, A3 => n60273, A4 => 
                           n60272, ZN => n60281);
   U3279 : AOI22_X1 port map( A1 => n51892, A2 => n53547, B1 => n52268, B2 => 
                           n53526, ZN => n60279);
   U3280 : AOI22_X1 port map( A1 => n52179, A2 => n52402, B1 => n51871, B2 => 
                           n53518, ZN => n60278);
   U3281 : AOI22_X1 port map( A1 => n52124, A2 => n53551, B1 => n52177, B2 => 
                           n52479, ZN => n60277);
   U3282 : AOI22_X1 port map( A1 => n52175, A2 => n52401, B1 => n52155, B2 => 
                           n53524, ZN => n60276);
   U3283 : NAND4_X1 port map( A1 => n60279, A2 => n60278, A3 => n60277, A4 => 
                           n60276, ZN => n60280);
   U3284 : AOI22_X1 port map( A1 => n60570, A2 => n60281, B1 => n60303, B2 => 
                           n60280, ZN => n60282);
   U3285 : OAI21_X1 port map( B1 => n60774, B2 => n60283, A => n60282, ZN => 
                           OUT1(22));
   U3286 : AOI22_X1 port map( A1 => n51575, A2 => n52417, B1 => n51793, B2 => 
                           n53533, ZN => n60287);
   U3287 : AOI22_X1 port map( A1 => n52333, A2 => n52410, B1 => n52028, B2 => 
                           n52407, ZN => n60286);
   U3288 : AOI22_X1 port map( A1 => n51795, A2 => n52418, B1 => n52266, B2 => 
                           n52413, ZN => n60285);
   U3289 : AOI22_X1 port map( A1 => n51670, A2 => n52415, B1 => n51794, B2 => 
                           n52408, ZN => n60284);
   U3290 : NAND4_X1 port map( A1 => n60287, A2 => n60286, A3 => n60285, A4 => 
                           n60284, ZN => n60293);
   U3291 : AOI22_X1 port map( A1 => n52286, A2 => n53554, B1 => n52259, B2 => 
                           n52406, ZN => n60291);
   U3292 : AOI22_X1 port map( A1 => n52314, A2 => n52404, B1 => n52016, B2 => 
                           n52409, ZN => n60290);
   U3293 : AOI22_X1 port map( A1 => n52258, A2 => n53558, B1 => n51796, B2 => 
                           n53553, ZN => n60289);
   U3294 : AOI22_X1 port map( A1 => n51819, A2 => n52411, B1 => n51799, B2 => 
                           n52416, ZN => n60288);
   U3295 : NAND4_X1 port map( A1 => n60291, A2 => n60290, A3 => n60289, A4 => 
                           n60288, ZN => n60292);
   U3296 : NOR2_X1 port map( A1 => n60293, A2 => n60292, ZN => n60306);
   U3297 : AOI22_X1 port map( A1 => n51909, A2 => n53547, B1 => n51918, B2 => 
                           n53546, ZN => n60297);
   U3298 : AOI22_X1 port map( A1 => n51913, A2 => n52482, B1 => n51919, B2 => 
                           n53527, ZN => n60296);
   U3299 : AOI22_X1 port map( A1 => n51702, A2 => n53551, B1 => n51509, B2 => 
                           n53525, ZN => n60295);
   U3300 : AOI22_X1 port map( A1 => n51526, A2 => n53518, B1 => n51927, B2 => 
                           n52481, ZN => n60294);
   U3301 : NAND4_X1 port map( A1 => n60297, A2 => n60296, A3 => n60295, A4 => 
                           n60294, ZN => n60304);
   U3302 : AOI22_X1 port map( A1 => n52261, A2 => n53551, B1 => n51607, B2 => 
                           n52401, ZN => n60301);
   U3303 : AOI22_X1 port map( A1 => n51621, A2 => n53527, B1 => n51798, B2 => 
                           n53550, ZN => n60300);
   U3304 : AOI22_X1 port map( A1 => n52260, A2 => n52481, B1 => n52350, B2 => 
                           n52402, ZN => n60299);
   U3305 : AOI22_X1 port map( A1 => n51797, A2 => n53547, B1 => n51602, B2 => 
                           n52482, ZN => n60298);
   U3306 : NAND4_X1 port map( A1 => n60301, A2 => n60300, A3 => n60299, A4 => 
                           n60298, ZN => n60302);
   U3307 : AOI22_X1 port map( A1 => n60570, A2 => n60304, B1 => n60303, B2 => 
                           n60302, ZN => n60305);
   U3308 : OAI21_X1 port map( B1 => n60774, B2 => n60306, A => n60305, ZN => 
                           OUT1(21));
   U3309 : AOI22_X1 port map( A1 => n52263, A2 => n52406, B1 => n52168, B2 => 
                           n52415, ZN => n60310);
   U3310 : AOI22_X1 port map( A1 => n51615, A2 => n52404, B1 => n52128, B2 => 
                           n52413, ZN => n60309);
   U3311 : AOI22_X1 port map( A1 => n51820, A2 => n52411, B1 => n51714, B2 => 
                           n52418, ZN => n60308);
   U3312 : AOI22_X1 port map( A1 => n52164, A2 => n52405, B1 => n52145, B2 => 
                           n53542, ZN => n60307);
   U3313 : NAND4_X1 port map( A1 => n60310, A2 => n60309, A3 => n60308, A4 => 
                           n60307, ZN => n60316);
   U3314 : AOI22_X1 port map( A1 => n52143, A2 => n52412, B1 => n51716, B2 => 
                           n52416, ZN => n60314);
   U3315 : AOI22_X1 port map( A1 => n51715, A2 => n53533, B1 => n52173, B2 => 
                           n52410, ZN => n60313);
   U3316 : AOI22_X1 port map( A1 => n51920, A2 => n52407, B1 => n51763, B2 => 
                           n52408, ZN => n60312);
   U3317 : AOI22_X1 port map( A1 => n51921, A2 => n52409, B1 => n51706, B2 => 
                           n53553, ZN => n60311);
   U3318 : NAND4_X1 port map( A1 => n60314, A2 => n60313, A3 => n60312, A4 => 
                           n60311, ZN => n60315);
   U3319 : NOR2_X1 port map( A1 => n60316, A2 => n60315, ZN => n60328);
   U3320 : AOI22_X1 port map( A1 => n51852, A2 => n53522, B1 => n52152, B2 => 
                           n53518, ZN => n60320);
   U3321 : AOI22_X1 port map( A1 => n52006, A2 => n53525, B1 => n52005, B2 => 
                           n53524, ZN => n60319);
   U3322 : AOI22_X1 port map( A1 => n51999, A2 => n53517, B1 => n52001, B2 => 
                           n53527, ZN => n60318);
   U3323 : AOI22_X1 port map( A1 => n52000, A2 => n53540, B1 => n52009, B2 => 
                           n53528, ZN => n60317);
   U3324 : NAND4_X1 port map( A1 => n60320, A2 => n60319, A3 => n60318, A4 => 
                           n60317, ZN => n60326);
   U3325 : AOI22_X1 port map( A1 => n52104, A2 => n53551, B1 => n52206, B2 => 
                           n53528, ZN => n60324);
   U3326 : AOI22_X1 port map( A1 => n51667, A2 => n53541, B1 => n51800, B2 => 
                           n53538, ZN => n60323);
   U3327 : AOI22_X1 port map( A1 => n52269, A2 => n53526, B1 => n52214, B2 => 
                           n53549, ZN => n60322);
   U3328 : AOI22_X1 port map( A1 => n51656, A2 => n53525, B1 => n51893, B2 => 
                           n53548, ZN => n60321);
   U3329 : NAND4_X1 port map( A1 => n60324, A2 => n60323, A3 => n60322, A4 => 
                           n60321, ZN => n60325);
   U3330 : AOI22_X1 port map( A1 => n60570, A2 => n60326, B1 => n60769, B2 => 
                           n60325, ZN => n60327);
   U3331 : OAI21_X1 port map( B1 => n60774, B2 => n60328, A => n60327, ZN => 
                           OUT1(20));
   U3332 : AOI22_X1 port map( A1 => n51713, A2 => n53537, B1 => n51718, B2 => 
                           n53555, ZN => n60332);
   U3333 : AOI22_X1 port map( A1 => n52318, A2 => n52404, B1 => n51711, B2 => 
                           n52403, ZN => n60331);
   U3334 : AOI22_X1 port map( A1 => n52294, A2 => n53543, B1 => n51659, B2 => 
                           n52405, ZN => n60330);
   U3335 : AOI22_X1 port map( A1 => n51560, A2 => n52417, B1 => n51821, B2 => 
                           n52411, ZN => n60329);
   U3336 : NAND4_X1 port map( A1 => n60332, A2 => n60331, A3 => n60330, A4 => 
                           n60329, ZN => n60338);
   U3337 : AOI22_X1 port map( A1 => n52027, A2 => n53556, B1 => n52015, B2 => 
                           n52409, ZN => n60336);
   U3338 : AOI22_X1 port map( A1 => n51537, A2 => n52413, B1 => n51553, B2 => 
                           n52412, ZN => n60335);
   U3339 : AOI22_X1 port map( A1 => n51691, A2 => n53533, B1 => n51764, B2 => 
                           n52408, ZN => n60334);
   U3340 : AOI22_X1 port map( A1 => n52332, A2 => n52410, B1 => n52262, B2 => 
                           n53535, ZN => n60333);
   U3341 : NAND4_X1 port map( A1 => n60336, A2 => n60335, A3 => n60334, A4 => 
                           n60333, ZN => n60337);
   U3342 : NOR2_X1 port map( A1 => n60338, A2 => n60337, ZN => n60350);
   U3343 : AOI22_X1 port map( A1 => n51926, A2 => n53541, B1 => n51512, B2 => 
                           n52482, ZN => n60342);
   U3344 : AOI22_X1 port map( A1 => n51514, A2 => n53528, B1 => n52371, B2 => 
                           n53518, ZN => n60341);
   U3345 : AOI22_X1 port map( A1 => n51700, A2 => n53522, B1 => n51916, B2 => 
                           n53526, ZN => n60340);
   U3346 : AOI22_X1 port map( A1 => n52067, A2 => n53539, B1 => n51508, B2 => 
                           n53547, ZN => n60339);
   U3347 : NAND4_X1 port map( A1 => n60342, A2 => n60341, A3 => n60340, A4 => 
                           n60339, ZN => n60348);
   U3348 : AOI22_X1 port map( A1 => n51611, A2 => n53549, B1 => n52270, B2 => 
                           n53540, ZN => n60346);
   U3349 : AOI22_X1 port map( A1 => n51783, A2 => n53518, B1 => n52343, B2 => 
                           n53546, ZN => n60345);
   U3350 : AOI22_X1 port map( A1 => n51894, A2 => n53548, B1 => n52340, B2 => 
                           n53541, ZN => n60344);
   U3351 : AOI22_X1 port map( A1 => n52345, A2 => n52402, B1 => n51516, B2 => 
                           n53522, ZN => n60343);
   U3352 : NAND4_X1 port map( A1 => n60346, A2 => n60345, A3 => n60344, A4 => 
                           n60343, ZN => n60347);
   U3353 : AOI22_X1 port map( A1 => n60570, A2 => n60348, B1 => n60769, B2 => 
                           n60347, ZN => n60349);
   U3354 : OAI21_X1 port map( B1 => n60774, B2 => n60350, A => n60349, ZN => 
                           OUT1(19));
   U3355 : AOI22_X1 port map( A1 => n51701, A2 => n52414, B1 => n51735, B2 => 
                           n53555, ZN => n60354);
   U3356 : AOI22_X1 port map( A1 => n51765, A2 => n52408, B1 => n51717, B2 => 
                           n52418, ZN => n60353);
   U3357 : AOI22_X1 port map( A1 => n52295, A2 => n53543, B1 => n52135, B2 => 
                           n53542, ZN => n60352);
   U3358 : AOI22_X1 port map( A1 => n52331, A2 => n52410, B1 => n52129, B2 => 
                           n53557, ZN => n60351);
   U3359 : NAND4_X1 port map( A1 => n60354, A2 => n60353, A3 => n60352, A4 => 
                           n60351, ZN => n60360);
   U3360 : AOI22_X1 port map( A1 => n52257, A2 => n52406, B1 => n51544, B2 => 
                           n53558, ZN => n60358);
   U3361 : AOI22_X1 port map( A1 => n51698, A2 => n52403, B1 => n52026, B2 => 
                           n52407, ZN => n60357);
   U3362 : AOI22_X1 port map( A1 => n52014, A2 => n52409, B1 => n51822, B2 => 
                           n52411, ZN => n60356);
   U3363 : AOI22_X1 port map( A1 => n52288, A2 => n52405, B1 => n52320, B2 => 
                           n52404, ZN => n60355);
   U3364 : NAND4_X1 port map( A1 => n60358, A2 => n60357, A3 => n60356, A4 => 
                           n60355, ZN => n60359);
   U3365 : NOR2_X1 port map( A1 => n60360, A2 => n60359, ZN => n60372);
   U3366 : AOI22_X1 port map( A1 => n51904, A2 => n53540, B1 => n51925, B2 => 
                           n53546, ZN => n60364);
   U3367 : AOI22_X1 port map( A1 => n51922, A2 => n53517, B1 => n52362, B2 => 
                           n53518, ZN => n60363);
   U3368 : AOI22_X1 port map( A1 => n51905, A2 => n52479, B1 => n51924, B2 => 
                           n52482, ZN => n60362);
   U3369 : AOI22_X1 port map( A1 => n52056, A2 => n53525, B1 => n51697, B2 => 
                           n52480, ZN => n60361);
   U3370 : NAND4_X1 port map( A1 => n60364, A2 => n60363, A3 => n60362, A4 => 
                           n60361, ZN => n60370);
   U3371 : AOI22_X1 port map( A1 => n52196, A2 => n53527, B1 => n52151, B2 => 
                           n53549, ZN => n60368);
   U3372 : AOI22_X1 port map( A1 => n51784, A2 => n53550, B1 => n51895, B2 => 
                           n53517, ZN => n60367);
   U3373 : AOI22_X1 port map( A1 => n51586, A2 => n53539, B1 => n52271, B2 => 
                           n52481, ZN => n60366);
   U3374 : AOI22_X1 port map( A1 => n51520, A2 => n53522, B1 => n52344, B2 => 
                           n52401, ZN => n60365);
   U3375 : NAND4_X1 port map( A1 => n60368, A2 => n60367, A3 => n60366, A4 => 
                           n60365, ZN => n60369);
   U3376 : AOI22_X1 port map( A1 => n60570, A2 => n60370, B1 => n60769, B2 => 
                           n60369, ZN => n60371);
   U3377 : OAI21_X1 port map( B1 => n60774, B2 => n60372, A => n60371, ZN => 
                           OUT1(18));
   U3378 : AOI22_X1 port map( A1 => n52013, A2 => n52409, B1 => n52024, B2 => 
                           n53556, ZN => n60376);
   U3379 : AOI22_X1 port map( A1 => n52326, A2 => n53544, B1 => n52296, B2 => 
                           n52415, ZN => n60375);
   U3380 : AOI22_X1 port map( A1 => n51805, A2 => n53553, B1 => n51802, B2 => 
                           n52414, ZN => n60374);
   U3381 : AOI22_X1 port map( A1 => n52225, A2 => n52417, B1 => n51814, B2 => 
                           n53536, ZN => n60373);
   U3382 : NAND4_X1 port map( A1 => n60376, A2 => n60375, A3 => n60374, A4 => 
                           n60373, ZN => n60382);
   U3383 : AOI22_X1 port map( A1 => n51808, A2 => n52416, B1 => n52224, B2 => 
                           n53557, ZN => n60380);
   U3384 : AOI22_X1 port map( A1 => n51804, A2 => n52418, B1 => n51803, B2 => 
                           n53552, ZN => n60379);
   U3385 : AOI22_X1 port map( A1 => n52292, A2 => n52405, B1 => n52299, B2 => 
                           n52404, ZN => n60378);
   U3386 : AOI22_X1 port map( A1 => n51590, A2 => n52406, B1 => n52251, B2 => 
                           n52412, ZN => n60377);
   U3387 : NAND4_X1 port map( A1 => n60380, A2 => n60379, A3 => n60378, A4 => 
                           n60377, ZN => n60381);
   U3388 : NOR2_X1 port map( A1 => n60382, A2 => n60381, ZN => n60394);
   U3389 : AOI22_X1 port map( A1 => n52330, A2 => n53518, B1 => n51971, B2 => 
                           n53546, ZN => n60386);
   U3390 : AOI22_X1 port map( A1 => n51962, A2 => n53547, B1 => n51970, B2 => 
                           n52479, ZN => n60385);
   U3391 : AOI22_X1 port map( A1 => n51965, A2 => n52481, B1 => n52061, B2 => 
                           n53525, ZN => n60384);
   U3392 : AOI22_X1 port map( A1 => n51960, A2 => n53524, B1 => n51766, B2 => 
                           n53522, ZN => n60383);
   U3393 : NAND4_X1 port map( A1 => n60386, A2 => n60385, A3 => n60384, A4 => 
                           n60383, ZN => n60392);
   U3394 : AOI22_X1 port map( A1 => n52213, A2 => n53524, B1 => n52200, B2 => 
                           n52479, ZN => n60390);
   U3395 : AOI22_X1 port map( A1 => n52209, A2 => n52401, B1 => n51807, B2 => 
                           n53550, ZN => n60389);
   U3396 : AOI22_X1 port map( A1 => n51806, A2 => n53517, B1 => n52221, B2 => 
                           n52480, ZN => n60388);
   U3397 : AOI22_X1 port map( A1 => n51585, A2 => n53526, B1 => n52240, B2 => 
                           n53525, ZN => n60387);
   U3398 : NAND4_X1 port map( A1 => n60390, A2 => n60389, A3 => n60388, A4 => 
                           n60387, ZN => n60391);
   U3399 : AOI22_X1 port map( A1 => n60570, A2 => n60392, B1 => n60769, B2 => 
                           n60391, ZN => n60393);
   U3400 : OAI21_X1 port map( B1 => n60774, B2 => n60394, A => n60393, ZN => 
                           OUT1(17));
   U3401 : AOI22_X1 port map( A1 => n51811, A2 => n52408, B1 => n52025, B2 => 
                           n52409, ZN => n60398);
   U3402 : AOI22_X1 port map( A1 => n52170, A2 => n53542, B1 => n51813, B2 => 
                           n52414, ZN => n60397);
   U3403 : AOI22_X1 port map( A1 => n52023, A2 => n52407, B1 => n51824, B2 => 
                           n52411, ZN => n60396);
   U3404 : AOI22_X1 port map( A1 => n52133, A2 => n53554, B1 => n52169, B2 => 
                           n53558, ZN => n60395);
   U3405 : NAND4_X1 port map( A1 => n60398, A2 => n60397, A3 => n60396, A4 => 
                           n60395, ZN => n60404);
   U3406 : AOI22_X1 port map( A1 => n51812, A2 => n53555, B1 => n51619, B2 => 
                           n52406, ZN => n60402);
   U3407 : AOI22_X1 port map( A1 => n51815, A2 => n53537, B1 => n52297, B2 => 
                           n52415, ZN => n60401);
   U3408 : AOI22_X1 port map( A1 => n52185, A2 => n52413, B1 => n52324, B2 => 
                           n52410, ZN => n60400);
   U3409 : AOI22_X1 port map( A1 => n51816, A2 => n52403, B1 => n51527, B2 => 
                           n52404, ZN => n60399);
   U3410 : NAND4_X1 port map( A1 => n60402, A2 => n60401, A3 => n60400, A4 => 
                           n60399, ZN => n60403);
   U3411 : NOR2_X1 port map( A1 => n60404, A2 => n60403, ZN => n60416);
   U3412 : CLKBUF_X1 port map( A => n60525, Z => n60771);
   U3413 : AOI22_X1 port map( A1 => n51964, A2 => n52402, B1 => n52071, B2 => 
                           n52482, ZN => n60408);
   U3414 : AOI22_X1 port map( A1 => n52070, A2 => n52401, B1 => n52072, B2 => 
                           n53517, ZN => n60407);
   U3415 : AOI22_X1 port map( A1 => n52069, A2 => n53527, B1 => n51696, B2 => 
                           n52480, ZN => n60406);
   U3416 : AOI22_X1 port map( A1 => n52309, A2 => n53550, B1 => n52073, B2 => 
                           n53526, ZN => n60405);
   U3417 : NAND4_X1 port map( A1 => n60408, A2 => n60407, A3 => n60406, A4 => 
                           n60405, ZN => n60414);
   U3418 : AOI22_X1 port map( A1 => n51599, A2 => n53528, B1 => n51810, B2 => 
                           n53550, ZN => n60412);
   U3419 : AOI22_X1 port map( A1 => n52197, A2 => n53522, B1 => n52154, B2 => 
                           n53524, ZN => n60411);
   U3420 : AOI22_X1 port map( A1 => n52195, A2 => n53526, B1 => n52337, B2 => 
                           n52479, ZN => n60410);
   U3421 : AOI22_X1 port map( A1 => n51809, A2 => n53547, B1 => n52349, B2 => 
                           n53525, ZN => n60409);
   U3422 : NAND4_X1 port map( A1 => n60412, A2 => n60411, A3 => n60410, A4 => 
                           n60409, ZN => n60413);
   U3423 : AOI22_X1 port map( A1 => n60771, A2 => n60414, B1 => n60769, B2 => 
                           n60413, ZN => n60415);
   U3424 : OAI21_X1 port map( B1 => n60774, B2 => n60416, A => n60415, ZN => 
                           OUT1(16));
   U3425 : AOI22_X1 port map( A1 => n51541, A2 => n52410, B1 => n52293, B2 => 
                           n52405, ZN => n60420);
   U3426 : AOI22_X1 port map( A1 => n51737, A2 => n52403, B1 => n52319, B2 => 
                           n52404, ZN => n60419);
   U3427 : AOI22_X1 port map( A1 => n51767, A2 => n52408, B1 => n52012, B2 => 
                           n52409, ZN => n60418);
   U3428 : AOI22_X1 port map( A1 => n52256, A2 => n53535, B1 => n51738, B2 => 
                           n52414, ZN => n60417);
   U3429 : NAND4_X1 port map( A1 => n60420, A2 => n60419, A3 => n60418, A4 => 
                           n60417, ZN => n60426);
   U3430 : AOI22_X1 port map( A1 => n51736, A2 => n52416, B1 => n52298, B2 => 
                           n52415, ZN => n60424);
   U3431 : AOI22_X1 port map( A1 => n51823, A2 => n52411, B1 => n52111, B2 => 
                           n52413, ZN => n60423);
   U3432 : AOI22_X1 port map( A1 => n52125, A2 => n52412, B1 => n51734, B2 => 
                           n52418, ZN => n60422);
   U3433 : AOI22_X1 port map( A1 => n52121, A2 => n53542, B1 => n52022, B2 => 
                           n53556, ZN => n60421);
   U3434 : NAND4_X1 port map( A1 => n60424, A2 => n60423, A3 => n60422, A4 => 
                           n60421, ZN => n60425);
   U3435 : NOR2_X1 port map( A1 => n60426, A2 => n60425, ZN => n60438);
   U3436 : AOI22_X1 port map( A1 => n51928, A2 => n53526, B1 => n51914, B2 => 
                           n53517, ZN => n60430);
   U3437 : AOI22_X1 port map( A1 => n52047, A2 => n53525, B1 => n51725, B2 => 
                           n53551, ZN => n60429);
   U3438 : AOI22_X1 port map( A1 => n51938, A2 => n53527, B1 => n52306, B2 => 
                           n53550, ZN => n60428);
   U3439 : AOI22_X1 port map( A1 => n51899, A2 => n53524, B1 => n51915, B2 => 
                           n53546, ZN => n60427);
   U3440 : NAND4_X1 port map( A1 => n60430, A2 => n60429, A3 => n60428, A4 => 
                           n60427, ZN => n60436);
   U3441 : AOI22_X1 port map( A1 => n51896, A2 => n53517, B1 => n52241, B2 => 
                           n52401, ZN => n60434);
   U3442 : AOI22_X1 port map( A1 => n52243, A2 => n53539, B1 => n52201, B2 => 
                           n53541, ZN => n60433);
   U3443 : AOI22_X1 port map( A1 => n52217, A2 => n52482, B1 => n52284, B2 => 
                           n53551, ZN => n60432);
   U3444 : AOI22_X1 port map( A1 => n51532, A2 => n53540, B1 => n51785, B2 => 
                           n53550, ZN => n60431);
   U3445 : NAND4_X1 port map( A1 => n60434, A2 => n60433, A3 => n60432, A4 => 
                           n60431, ZN => n60435);
   U3446 : AOI22_X1 port map( A1 => n60525, A2 => n60436, B1 => n60769, B2 => 
                           n60435, ZN => n60437);
   U3447 : OAI21_X1 port map( B1 => n60774, B2 => n60438, A => n60437, ZN => 
                           OUT1(15));
   U3448 : AOI22_X1 port map( A1 => n51703, A2 => n52403, B1 => n52144, B2 => 
                           n52412, ZN => n60442);
   U3449 : AOI22_X1 port map( A1 => n52131, A2 => n52413, B1 => n52146, B2 => 
                           n53542, ZN => n60441);
   U3450 : AOI22_X1 port map( A1 => n51768, A2 => n52408, B1 => n51747, B2 => 
                           n52414, ZN => n60440);
   U3451 : AOI22_X1 port map( A1 => n51482, A2 => n52409, B1 => n52300, B2 => 
                           n53543, ZN => n60439);
   U3452 : NAND4_X1 port map( A1 => n60442, A2 => n60441, A3 => n60440, A4 => 
                           n60439, ZN => n60448);
   U3453 : AOI22_X1 port map( A1 => n51739, A2 => n52416, B1 => n52255, B2 => 
                           n52406, ZN => n60446);
   U3454 : AOI22_X1 port map( A1 => n52021, A2 => n53556, B1 => n52312, B2 => 
                           n52404, ZN => n60445);
   U3455 : AOI22_X1 port map( A1 => n51826, A2 => n53536, B1 => n52291, B2 => 
                           n53554, ZN => n60444);
   U3456 : AOI22_X1 port map( A1 => n51710, A2 => n52418, B1 => n52323, B2 => 
                           n52410, ZN => n60443);
   U3457 : NAND4_X1 port map( A1 => n60446, A2 => n60445, A3 => n60444, A4 => 
                           n60443, ZN => n60447);
   U3458 : NOR2_X1 port map( A1 => n60448, A2 => n60447, ZN => n60460);
   U3459 : AOI22_X1 port map( A1 => n51483, A2 => n53540, B1 => n52048, B2 => 
                           n53517, ZN => n60452);
   U3460 : AOI22_X1 port map( A1 => n51956, A2 => n53539, B1 => n51720, B2 => 
                           n53522, ZN => n60451);
   U3461 : AOI22_X1 port map( A1 => n52046, A2 => n53541, B1 => n52045, B2 => 
                           n53528, ZN => n60450);
   U3462 : AOI22_X1 port map( A1 => n52049, A2 => n53549, B1 => n52387, B2 => 
                           n53550, ZN => n60449);
   U3463 : NAND4_X1 port map( A1 => n60452, A2 => n60451, A3 => n60450, A4 => 
                           n60449, ZN => n60458);
   U3464 : AOI22_X1 port map( A1 => n51897, A2 => n53517, B1 => n52283, B2 => 
                           n53551, ZN => n60456);
   U3465 : AOI22_X1 port map( A1 => n51786, A2 => n53550, B1 => n52192, B2 => 
                           n53539, ZN => n60455);
   U3466 : AOI22_X1 port map( A1 => n52348, A2 => n53528, B1 => n52147, B2 => 
                           n53549, ZN => n60454);
   U3467 : AOI22_X1 port map( A1 => n52190, A2 => n53541, B1 => n52272, B2 => 
                           n53526, ZN => n60453);
   U3468 : NAND4_X1 port map( A1 => n60456, A2 => n60455, A3 => n60454, A4 => 
                           n60453, ZN => n60457);
   U3469 : AOI22_X1 port map( A1 => n60570, A2 => n60458, B1 => n60769, B2 => 
                           n60457, ZN => n60459);
   U3470 : OAI21_X1 port map( B1 => n60774, B2 => n60460, A => n60459, ZN => 
                           OUT1(14));
   U3471 : AOI22_X1 port map( A1 => n51755, A2 => n52403, B1 => n52088, B2 => 
                           n52413, ZN => n60464);
   U3472 : AOI22_X1 port map( A1 => n52322, A2 => n52410, B1 => n52254, B2 => 
                           n53535, ZN => n60463);
   U3473 : AOI22_X1 port map( A1 => n51753, A2 => n52418, B1 => n52290, B2 => 
                           n53554, ZN => n60462);
   U3474 : AOI22_X1 port map( A1 => n52020, A2 => n52407, B1 => n51825, B2 => 
                           n52411, ZN => n60461);
   U3475 : NAND4_X1 port map( A1 => n60464, A2 => n60463, A3 => n60462, A4 => 
                           n60461, ZN => n60470);
   U3476 : AOI22_X1 port map( A1 => n51769, A2 => n52408, B1 => n51740, B2 => 
                           n53555, ZN => n60468);
   U3477 : AOI22_X1 port map( A1 => n52311, A2 => n52404, B1 => n52029, B2 => 
                           n53534, ZN => n60467);
   U3478 : AOI22_X1 port map( A1 => n52301, A2 => n53543, B1 => n52080, B2 => 
                           n52412, ZN => n60466);
   U3479 : AOI22_X1 port map( A1 => n52076, A2 => n52417, B1 => n51750, B2 => 
                           n52414, ZN => n60465);
   U3480 : NAND4_X1 port map( A1 => n60468, A2 => n60467, A3 => n60466, A4 => 
                           n60465, ZN => n60469);
   U3481 : NOR2_X1 port map( A1 => n60470, A2 => n60469, ZN => n60482);
   U3482 : AOI22_X1 port map( A1 => n52050, A2 => n52481, B1 => n52052, B2 => 
                           n53527, ZN => n60474);
   U3483 : AOI22_X1 port map( A1 => n52053, A2 => n52401, B1 => n52347, B2 => 
                           n53550, ZN => n60473);
   U3484 : AOI22_X1 port map( A1 => n52051, A2 => n52402, B1 => n52054, B2 => 
                           n53517, ZN => n60472);
   U3485 : AOI22_X1 port map( A1 => n51510, A2 => n53549, B1 => n51712, B2 => 
                           n53522, ZN => n60471);
   U3486 : NAND4_X1 port map( A1 => n60474, A2 => n60473, A3 => n60472, A4 => 
                           n60471, ZN => n60480);
   U3487 : AOI22_X1 port map( A1 => n51898, A2 => n53517, B1 => n52357, B2 => 
                           n53546, ZN => n60478);
   U3488 : AOI22_X1 port map( A1 => n51787, A2 => n53550, B1 => n52346, B2 => 
                           n53525, ZN => n60477);
   U3489 : AOI22_X1 port map( A1 => n52282, A2 => n52480, B1 => n52153, B2 => 
                           n53524, ZN => n60476);
   U3490 : AOI22_X1 port map( A1 => n52273, A2 => n52481, B1 => n52353, B2 => 
                           n53527, ZN => n60475);
   U3491 : NAND4_X1 port map( A1 => n60478, A2 => n60477, A3 => n60476, A4 => 
                           n60475, ZN => n60479);
   U3492 : AOI22_X1 port map( A1 => n60771, A2 => n60480, B1 => n60769, B2 => 
                           n60479, ZN => n60481);
   U3493 : OAI21_X1 port map( B1 => n60774, B2 => n60482, A => n60481, ZN => 
                           OUT1(13));
   U3494 : AOI22_X1 port map( A1 => n52316, A2 => n52410, B1 => n52321, B2 => 
                           n52404, ZN => n60486);
   U3495 : AOI22_X1 port map( A1 => n52085, A2 => n52412, B1 => n51757, B2 => 
                           n53533, ZN => n60485);
   U3496 : AOI22_X1 port map( A1 => n51741, A2 => n53555, B1 => n51770, B2 => 
                           n53552, ZN => n60484);
   U3497 : AOI22_X1 port map( A1 => n52253, A2 => n53535, B1 => n51759, B2 => 
                           n52403, ZN => n60483);
   U3498 : NAND4_X1 port map( A1 => n60486, A2 => n60485, A3 => n60484, A4 => 
                           n60483, ZN => n60492);
   U3499 : AOI22_X1 port map( A1 => n51476, A2 => n52409, B1 => n51669, B2 => 
                           n52405, ZN => n60490);
   U3500 : AOI22_X1 port map( A1 => n51758, A2 => n52418, B1 => n51829, B2 => 
                           n52411, ZN => n60489);
   U3501 : AOI22_X1 port map( A1 => n52090, A2 => n52417, B1 => n51449, B2 => 
                           n52407, ZN => n60488);
   U3502 : AOI22_X1 port map( A1 => n52092, A2 => n53557, B1 => n52302, B2 => 
                           n52415, ZN => n60487);
   U3503 : NAND4_X1 port map( A1 => n60490, A2 => n60489, A3 => n60488, A4 => 
                           n60487, ZN => n60491);
   U3504 : NOR2_X1 port map( A1 => n60492, A2 => n60491, ZN => n60504);
   U3505 : AOI22_X1 port map( A1 => n52060, A2 => n53517, B1 => n52058, B2 => 
                           n53528, ZN => n60496);
   U3506 : AOI22_X1 port map( A1 => n51513, A2 => n53541, B1 => n51632, B2 => 
                           n53550, ZN => n60495);
   U3507 : AOI22_X1 port map( A1 => n52059, A2 => n52482, B1 => n52057, B2 => 
                           n53539, ZN => n60494);
   U3508 : AOI22_X1 port map( A1 => n52055, A2 => n53526, B1 => n51705, B2 => 
                           n53551, ZN => n60493);
   U3509 : NAND4_X1 port map( A1 => n60496, A2 => n60495, A3 => n60494, A4 => 
                           n60493, ZN => n60502);
   U3510 : AOI22_X1 port map( A1 => n52189, A2 => n52402, B1 => n52159, B2 => 
                           n53524, ZN => n60500);
   U3511 : AOI22_X1 port map( A1 => n51788, A2 => n53550, B1 => n51778, B2 => 
                           n53547, ZN => n60499);
   U3512 : AOI22_X1 port map( A1 => n52188, A2 => n53527, B1 => n52274, B2 => 
                           n52481, ZN => n60498);
   U3513 : AOI22_X1 port map( A1 => n52281, A2 => n53551, B1 => n52351, B2 => 
                           n53528, ZN => n60497);
   U3514 : NAND4_X1 port map( A1 => n60500, A2 => n60499, A3 => n60498, A4 => 
                           n60497, ZN => n60501);
   U3515 : AOI22_X1 port map( A1 => n60570, A2 => n60502, B1 => n60769, B2 => 
                           n60501, ZN => n60503);
   U3516 : OAI21_X1 port map( B1 => n60774, B2 => n60504, A => n60503, ZN => 
                           OUT1(12));
   U3517 : AOI22_X1 port map( A1 => n52328, A2 => n53544, B1 => n52303, B2 => 
                           n52415, ZN => n60508);
   U3518 : AOI22_X1 port map( A1 => n51771, A2 => n52414, B1 => n52098, B2 => 
                           n52417, ZN => n60507);
   U3519 : AOI22_X1 port map( A1 => n52109, A2 => n53557, B1 => n52030, B2 => 
                           n53534, ZN => n60506);
   U3520 : AOI22_X1 port map( A1 => n52019, A2 => n53556, B1 => n52095, B2 => 
                           n52412, ZN => n60505);
   U3521 : NAND4_X1 port map( A1 => n60508, A2 => n60507, A3 => n60506, A4 => 
                           n60505, ZN => n60514);
   U3522 : AOI22_X1 port map( A1 => n51773, A2 => n53537, B1 => n51772, B2 => 
                           n53552, ZN => n60512);
   U3523 : AOI22_X1 port map( A1 => n52289, A2 => n52405, B1 => n52313, B2 => 
                           n52404, ZN => n60511);
   U3524 : AOI22_X1 port map( A1 => n51774, A2 => n53553, B1 => n51742, B2 => 
                           n52416, ZN => n60510);
   U3525 : AOI22_X1 port map( A1 => n52252, A2 => n52406, B1 => n51801, B2 => 
                           n53536, ZN => n60509);
   U3526 : NAND4_X1 port map( A1 => n60512, A2 => n60511, A3 => n60510, A4 => 
                           n60509, ZN => n60513);
   U3527 : NOR2_X1 port map( A1 => n60514, A2 => n60513, ZN => n60527);
   U3528 : AOI22_X1 port map( A1 => n52068, A2 => n53547, B1 => n52064, B2 => 
                           n52479, ZN => n60518);
   U3529 : AOI22_X1 port map( A1 => n52065, A2 => n53546, B1 => n52382, B2 => 
                           n53518, ZN => n60517);
   U3530 : AOI22_X1 port map( A1 => n51695, A2 => n53551, B1 => n52063, B2 => 
                           n53539, ZN => n60516);
   U3531 : AOI22_X1 port map( A1 => n52066, A2 => n53549, B1 => n52062, B2 => 
                           n53540, ZN => n60515);
   U3532 : NAND4_X1 port map( A1 => n60518, A2 => n60517, A3 => n60516, A4 => 
                           n60515, ZN => n60524);
   U3533 : AOI22_X1 port map( A1 => n52278, A2 => n52480, B1 => n52352, B2 => 
                           n53546, ZN => n60522);
   U3534 : AOI22_X1 port map( A1 => n52157, A2 => n52482, B1 => n52275, B2 => 
                           n53540, ZN => n60521);
   U3535 : AOI22_X1 port map( A1 => n52355, A2 => n52479, B1 => n51789, B2 => 
                           n53550, ZN => n60520);
   U3536 : AOI22_X1 port map( A1 => n51779, A2 => n53517, B1 => n52339, B2 => 
                           n53525, ZN => n60519);
   U3537 : NAND4_X1 port map( A1 => n60522, A2 => n60521, A3 => n60520, A4 => 
                           n60519, ZN => n60523);
   U3538 : AOI22_X1 port map( A1 => n60525, A2 => n60524, B1 => n60769, B2 => 
                           n60523, ZN => n60526);
   U3539 : OAI21_X1 port map( B1 => n60774, B2 => n60527, A => n60526, ZN => 
                           OUT1(11));
   U3540 : AOI22_X1 port map( A1 => n51744, A2 => n52416, B1 => n51998, B2 => 
                           n53534, ZN => n60531);
   U3541 : AOI22_X1 port map( A1 => n51581, A2 => n52405, B1 => n51997, B2 => 
                           n52407, ZN => n60530);
   U3542 : AOI22_X1 port map( A1 => n51562, A2 => n53557, B1 => n51578, B2 => 
                           n52406, ZN => n60529);
   U3543 : AOI22_X1 port map( A1 => n51754, A2 => n52418, B1 => n52360, B2 => 
                           n52404, ZN => n60528);
   U3544 : NAND4_X1 port map( A1 => n60531, A2 => n60530, A3 => n60529, A4 => 
                           n60528, ZN => n60537);
   U3545 : AOI22_X1 port map( A1 => n51579, A2 => n52415, B1 => n51582, B2 => 
                           n52410, ZN => n60535);
   U3546 : AOI22_X1 port map( A1 => n52160, A2 => n53542, B1 => n51761, B2 => 
                           n53552, ZN => n60534);
   U3547 : AOI22_X1 port map( A1 => n51733, A2 => n53536, B1 => n52112, B2 => 
                           n52412, ZN => n60533);
   U3548 : AOI22_X1 port map( A1 => n51726, A2 => n53533, B1 => n51752, B2 => 
                           n53553, ZN => n60532);
   U3549 : NAND4_X1 port map( A1 => n60535, A2 => n60534, A3 => n60533, A4 => 
                           n60532, ZN => n60536);
   U3550 : NOR2_X1 port map( A1 => n60537, A2 => n60536, ZN => n60549);
   U3551 : AOI22_X1 port map( A1 => n51972, A2 => n53524, B1 => n51976, B2 => 
                           n53528, ZN => n60541);
   U3552 : AOI22_X1 port map( A1 => n51981, A2 => n53527, B1 => n52162, B2 => 
                           n53538, ZN => n60540);
   U3553 : AOI22_X1 port map( A1 => n51974, A2 => n53517, B1 => n51833, B2 => 
                           n52480, ZN => n60539);
   U3554 : AOI22_X1 port map( A1 => n51969, A2 => n53526, B1 => n51978, B2 => 
                           n53525, ZN => n60538);
   U3555 : NAND4_X1 port map( A1 => n60541, A2 => n60540, A3 => n60539, A4 => 
                           n60538, ZN => n60547);
   U3556 : AOI22_X1 port map( A1 => n51601, A2 => n53524, B1 => n51792, B2 => 
                           n53518, ZN => n60545);
   U3557 : AOI22_X1 port map( A1 => n51608, A2 => n53539, B1 => n51780, B2 => 
                           n53517, ZN => n60544);
   U3558 : AOI22_X1 port map( A1 => n52358, A2 => n53546, B1 => n52163, B2 => 
                           n53526, ZN => n60543);
   U3559 : AOI22_X1 port map( A1 => n51626, A2 => n53551, B1 => n51616, B2 => 
                           n53541, ZN => n60542);
   U3560 : NAND4_X1 port map( A1 => n60545, A2 => n60544, A3 => n60543, A4 => 
                           n60542, ZN => n60546);
   U3561 : AOI22_X1 port map( A1 => n60570, A2 => n60547, B1 => n60769, B2 => 
                           n60546, ZN => n60548);
   U3562 : OAI21_X1 port map( B1 => n60727, B2 => n60549, A => n60548, ZN => 
                           OUT1(10));
   U3563 : AOI22_X1 port map( A1 => n52287, A2 => n53554, B1 => n52018, B2 => 
                           n52407, ZN => n60553);
   U3564 : AOI22_X1 port map( A1 => n52031, A2 => n53534, B1 => n51775, B2 => 
                           n52408, ZN => n60552);
   U3565 : AOI22_X1 port map( A1 => n51729, A2 => n52411, B1 => n52304, B2 => 
                           n52415, ZN => n60551);
   U3566 : AOI22_X1 port map( A1 => n51751, A2 => n53553, B1 => n51545, B2 => 
                           n52404, ZN => n60550);
   U3567 : NAND4_X1 port map( A1 => n60553, A2 => n60552, A3 => n60551, A4 => 
                           n60550, ZN => n60559);
   U3568 : AOI22_X1 port map( A1 => n52223, A2 => n52406, B1 => n51745, B2 => 
                           n52416, ZN => n60557);
   U3569 : AOI22_X1 port map( A1 => n52126, A2 => n53557, B1 => n52327, B2 => 
                           n52410, ZN => n60556);
   U3570 : AOI22_X1 port map( A1 => n51539, A2 => n53558, B1 => n51533, B2 => 
                           n53542, ZN => n60555);
   U3571 : AOI22_X1 port map( A1 => n51748, A2 => n52414, B1 => n51730, B2 => 
                           n53537, ZN => n60554);
   U3572 : NAND4_X1 port map( A1 => n60557, A2 => n60556, A3 => n60555, A4 => 
                           n60554, ZN => n60558);
   U3573 : NOR2_X1 port map( A1 => n60559, A2 => n60558, ZN => n60572);
   U3574 : AOI22_X1 port map( A1 => n52037, A2 => n52479, B1 => n52033, B2 => 
                           n53539, ZN => n60563);
   U3575 : AOI22_X1 port map( A1 => n51552, A2 => n53518, B1 => n52034, B2 => 
                           n52482, ZN => n60562);
   U3576 : AOI22_X1 port map( A1 => n52035, A2 => n53528, B1 => n52038, B2 => 
                           n53540, ZN => n60561);
   U3577 : AOI22_X1 port map( A1 => n51731, A2 => n53551, B1 => n52036, B2 => 
                           n53548, ZN => n60560);
   U3578 : NAND4_X1 port map( A1 => n60563, A2 => n60562, A3 => n60561, A4 => 
                           n60560, ZN => n60569);
   U3579 : AOI22_X1 port map( A1 => n52148, A2 => n53524, B1 => n52359, B2 => 
                           n53525, ZN => n60567);
   U3580 : AOI22_X1 port map( A1 => n52277, A2 => n53522, B1 => n52279, B2 => 
                           n52481, ZN => n60566);
   U3581 : AOI22_X1 port map( A1 => n51592, A2 => n53528, B1 => n51791, B2 => 
                           n53518, ZN => n60565);
   U3582 : AOI22_X1 port map( A1 => n51781, A2 => n53517, B1 => n52193, B2 => 
                           n53527, ZN => n60564);
   U3583 : NAND4_X1 port map( A1 => n60567, A2 => n60566, A3 => n60565, A4 => 
                           n60564, ZN => n60568);
   U3584 : AOI22_X1 port map( A1 => n60570, A2 => n60569, B1 => n60769, B2 => 
                           n60568, ZN => n60571);
   U3585 : OAI21_X1 port map( B1 => n60774, B2 => n60572, A => n60571, ZN => 
                           OUT1(9));
   U3586 : AOI22_X1 port map( A1 => n52134, A2 => n52417, B1 => n51746, B2 => 
                           n52416, ZN => n60576);
   U3587 : AOI22_X1 port map( A1 => n51776, A2 => n52408, B1 => n51728, B2 => 
                           n53537, ZN => n60575);
   U3588 : AOI22_X1 port map( A1 => n52130, A2 => n53557, B1 => n52329, B2 => 
                           n52404, ZN => n60574);
   U3589 : AOI22_X1 port map( A1 => n52032, A2 => n52409, B1 => n51719, B2 => 
                           n53536, ZN => n60573);
   U3590 : NAND4_X1 port map( A1 => n60576, A2 => n60575, A3 => n60574, A4 => 
                           n60573, ZN => n60582);
   U3591 : AOI22_X1 port map( A1 => n52132, A2 => n53558, B1 => n52017, B2 => 
                           n53556, ZN => n60580);
   U3592 : AOI22_X1 port map( A1 => n52325, A2 => n52410, B1 => n52305, B2 => 
                           n52415, ZN => n60579);
   U3593 : AOI22_X1 port map( A1 => n51727, A2 => n52403, B1 => n51749, B2 => 
                           n52414, ZN => n60578);
   U3594 : AOI22_X1 port map( A1 => n52334, A2 => n52405, B1 => n52222, B2 => 
                           n52406, ZN => n60577);
   U3595 : NAND4_X1 port map( A1 => n60580, A2 => n60579, A3 => n60578, A4 => 
                           n60577, ZN => n60581);
   U3596 : NOR2_X1 port map( A1 => n60582, A2 => n60581, ZN => n60594);
   U3597 : AOI22_X1 port map( A1 => n52039, A2 => n53540, B1 => n52041, B2 => 
                           n53528, ZN => n60586);
   U3598 : AOI22_X1 port map( A1 => n52040, A2 => n53548, B1 => n51724, B2 => 
                           n53522, ZN => n60585);
   U3599 : AOI22_X1 port map( A1 => n52043, A2 => n52479, B1 => n52307, B2 => 
                           n53518, ZN => n60584);
   U3600 : AOI22_X1 port map( A1 => n52042, A2 => n53525, B1 => n52044, B2 => 
                           n53549, ZN => n60583);
   U3601 : NAND4_X1 port map( A1 => n60586, A2 => n60585, A3 => n60584, A4 => 
                           n60583, ZN => n60592);
   U3602 : AOI22_X1 port map( A1 => n51782, A2 => n53548, B1 => n52194, B2 => 
                           n53539, ZN => n60590);
   U3603 : AOI22_X1 port map( A1 => n52356, A2 => n53528, B1 => n52276, B2 => 
                           n52480, ZN => n60589);
   U3604 : AOI22_X1 port map( A1 => n52280, A2 => n53526, B1 => n52150, B2 => 
                           n53524, ZN => n60588);
   U3605 : AOI22_X1 port map( A1 => n51790, A2 => n53538, B1 => n52191, B2 => 
                           n53541, ZN => n60587);
   U3606 : NAND4_X1 port map( A1 => n60590, A2 => n60589, A3 => n60588, A4 => 
                           n60587, ZN => n60591);
   U3607 : AOI22_X1 port map( A1 => n60771, A2 => n60592, B1 => n60769, B2 => 
                           n60591, ZN => n60593);
   U3608 : OAI21_X1 port map( B1 => n60774, B2 => n60594, A => n60593, ZN => 
                           OUT1(8));
   U3609 : AOI22_X1 port map( A1 => n52186, A2 => n53543, B1 => n52187, B2 => 
                           n52410, ZN => n60598);
   U3610 : AOI22_X1 port map( A1 => n51888, A2 => n53553, B1 => n51967, B2 => 
                           n52409, ZN => n60597);
   U3611 : AOI22_X1 port map( A1 => n51881, A2 => n52408, B1 => n52184, B2 => 
                           n53545, ZN => n60596);
   U3612 : AOI22_X1 port map( A1 => n52091, A2 => n52413, B1 => n51887, B2 => 
                           n52418, ZN => n60595);
   U3613 : NAND4_X1 port map( A1 => n60598, A2 => n60597, A3 => n60596, A4 => 
                           n60595, ZN => n60604);
   U3614 : AOI22_X1 port map( A1 => n52117, A2 => n52412, B1 => n52083, B2 => 
                           n52406, ZN => n60602);
   U3615 : AOI22_X1 port map( A1 => n51874, A2 => n52416, B1 => n51863, B2 => 
                           n53536, ZN => n60601);
   U3616 : AOI22_X1 port map( A1 => n52183, A2 => n52405, B1 => n51968, B2 => 
                           n53556, ZN => n60600);
   U3617 : AOI22_X1 port map( A1 => n51891, A2 => n52414, B1 => n52123, B2 => 
                           n52417, ZN => n60599);
   U3618 : NAND4_X1 port map( A1 => n60602, A2 => n60601, A3 => n60600, A4 => 
                           n60599, ZN => n60603);
   U3619 : NOR2_X1 port map( A1 => n60604, A2 => n60603, ZN => n60616);
   U3620 : AOI22_X1 port map( A1 => n51994, A2 => n52481, B1 => n51983, B2 => 
                           n53548, ZN => n60608);
   U3621 : AOI22_X1 port map( A1 => n52156, A2 => n53518, B1 => n52008, B2 => 
                           n53525, ZN => n60607);
   U3622 : AOI22_X1 port map( A1 => n52003, A2 => n53546, B1 => n52004, B2 => 
                           n52482, ZN => n60606);
   U3623 : AOI22_X1 port map( A1 => n51851, A2 => n53551, B1 => n51996, B2 => 
                           n53527, ZN => n60605);
   U3624 : NAND4_X1 port map( A1 => n60608, A2 => n60607, A3 => n60606, A4 => 
                           n60605, ZN => n60614);
   U3625 : AOI22_X1 port map( A1 => n52208, A2 => n52480, B1 => n52247, B2 => 
                           n53539, ZN => n60612);
   U3626 : AOI22_X1 port map( A1 => n51890, A2 => n53548, B1 => n51830, B2 => 
                           n53538, ZN => n60611);
   U3627 : AOI22_X1 port map( A1 => n51674, A2 => n52481, B1 => n52245, B2 => 
                           n53546, ZN => n60610);
   U3628 : AOI22_X1 port map( A1 => n52219, A2 => n53549, B1 => n52249, B2 => 
                           n52479, ZN => n60609);
   U3629 : NAND4_X1 port map( A1 => n60612, A2 => n60611, A3 => n60610, A4 => 
                           n60609, ZN => n60613);
   U3630 : AOI22_X1 port map( A1 => n60771, A2 => n60614, B1 => n60769, B2 => 
                           n60613, ZN => n60615);
   U3631 : OAI21_X1 port map( B1 => n60774, B2 => n60616, A => n60615, ZN => 
                           OUT1(7));
   U3632 : AOI22_X1 port map( A1 => n51868, A2 => n52408, B1 => n52370, B2 => 
                           n52405, ZN => n60620);
   U3633 : AOI22_X1 port map( A1 => n51995, A2 => n52407, B1 => n51873, B2 => 
                           n53537, ZN => n60619);
   U3634 : AOI22_X1 port map( A1 => n52122, A2 => n52413, B1 => n51982, B2 => 
                           n53534, ZN => n60618);
   U3635 : AOI22_X1 port map( A1 => n52084, A2 => n52412, B1 => n52074, B2 => 
                           n52406, ZN => n60617);
   U3636 : NAND4_X1 port map( A1 => n60620, A2 => n60619, A3 => n60618, A4 => 
                           n60617, ZN => n60626);
   U3637 : AOI22_X1 port map( A1 => n52385, A2 => n53545, B1 => n51877, B2 => 
                           n53555, ZN => n60624);
   U3638 : AOI22_X1 port map( A1 => n51872, A2 => n52414, B1 => n52336, B2 => 
                           n52410, ZN => n60623);
   U3639 : AOI22_X1 port map( A1 => n51889, A2 => n52411, B1 => n52373, B2 => 
                           n52415, ZN => n60622);
   U3640 : AOI22_X1 port map( A1 => n51884, A2 => n52403, B1 => n52087, B2 => 
                           n52417, ZN => n60621);
   U3641 : NAND4_X1 port map( A1 => n60624, A2 => n60623, A3 => n60622, A4 => 
                           n60621, ZN => n60625);
   U3642 : NOR2_X1 port map( A1 => n60626, A2 => n60625, ZN => n60638);
   U3643 : AOI22_X1 port map( A1 => n52342, A2 => n53518, B1 => n51910, B2 => 
                           n52401, ZN => n60630);
   U3644 : AOI22_X1 port map( A1 => n51721, A2 => n52480, B1 => n51950, B2 => 
                           n53539, ZN => n60629);
   U3645 : AOI22_X1 port map( A1 => n51912, A2 => n53548, B1 => n51911, B2 => 
                           n53524, ZN => n60628);
   U3646 : AOI22_X1 port map( A1 => n51935, A2 => n53541, B1 => n51901, B2 => 
                           n53526, ZN => n60627);
   U3647 : NAND4_X1 port map( A1 => n60630, A2 => n60629, A3 => n60628, A4 => 
                           n60627, ZN => n60636);
   U3648 : AOI22_X1 port map( A1 => n52236, A2 => n53527, B1 => n52078, B2 => 
                           n53540, ZN => n60634);
   U3649 : AOI22_X1 port map( A1 => n51828, A2 => n53538, B1 => n52232, B2 => 
                           n53525, ZN => n60633);
   U3650 : AOI22_X1 port map( A1 => n52215, A2 => n53524, B1 => n52204, B2 => 
                           n53522, ZN => n60632);
   U3651 : AOI22_X1 port map( A1 => n51878, A2 => n53548, B1 => n52235, B2 => 
                           n53546, ZN => n60631);
   U3652 : NAND4_X1 port map( A1 => n60634, A2 => n60633, A3 => n60632, A4 => 
                           n60631, ZN => n60635);
   U3653 : AOI22_X1 port map( A1 => n60771, A2 => n60636, B1 => n60769, B2 => 
                           n60635, ZN => n60637);
   U3654 : OAI21_X1 port map( B1 => n60774, B2 => n60638, A => n60637, ZN => 
                           OUT1(6));
   U3655 : AOI22_X1 port map( A1 => n52093, A2 => n53542, B1 => n52379, B2 => 
                           n52410, ZN => n60642);
   U3656 : AOI22_X1 port map( A1 => n51993, A2 => n52407, B1 => n51860, B2 => 
                           n52411, ZN => n60641);
   U3657 : AOI22_X1 port map( A1 => n51850, A2 => n52408, B1 => n52089, B2 => 
                           n52412, ZN => n60640);
   U3658 : AOI22_X1 port map( A1 => n51861, A2 => n52403, B1 => n51870, B2 => 
                           n53533, ZN => n60639);
   U3659 : NAND4_X1 port map( A1 => n60642, A2 => n60641, A3 => n60640, A4 => 
                           n60639, ZN => n60648);
   U3660 : AOI22_X1 port map( A1 => n52110, A2 => n52406, B1 => n51865, B2 => 
                           n52418, ZN => n60646);
   U3661 : AOI22_X1 port map( A1 => n52377, A2 => n52404, B1 => n51875, B2 => 
                           n52416, ZN => n60645);
   U3662 : AOI22_X1 port map( A1 => n52366, A2 => n52405, B1 => n52105, B2 => 
                           n52413, ZN => n60644);
   U3663 : AOI22_X1 port map( A1 => n51985, A2 => n52409, B1 => n52341, B2 => 
                           n53543, ZN => n60643);
   U3664 : NAND4_X1 port map( A1 => n60646, A2 => n60645, A3 => n60644, A4 => 
                           n60643, ZN => n60647);
   U3665 : NOR2_X1 port map( A1 => n60648, A2 => n60647, ZN => n60660);
   U3666 : AOI22_X1 port map( A1 => n51917, A2 => n53525, B1 => n52354, B2 => 
                           n53538, ZN => n60652);
   U3667 : AOI22_X1 port map( A1 => n51708, A2 => n53522, B1 => n51934, B2 => 
                           n52479, ZN => n60651);
   U3668 : AOI22_X1 port map( A1 => n51929, A2 => n53524, B1 => n51908, B2 => 
                           n52481, ZN => n60650);
   U3669 : AOI22_X1 port map( A1 => n51907, A2 => n53528, B1 => n51902, B2 => 
                           n53517, ZN => n60649);
   U3670 : NAND4_X1 port map( A1 => n60652, A2 => n60651, A3 => n60650, A4 => 
                           n60649, ZN => n60658);
   U3671 : AOI22_X1 port map( A1 => n52246, A2 => n53527, B1 => n51832, B2 => 
                           n53518, ZN => n60656);
   U3672 : AOI22_X1 port map( A1 => n52233, A2 => n52402, B1 => n51857, B2 => 
                           n53548, ZN => n60655);
   U3673 : AOI22_X1 port map( A1 => n52086, A2 => n53526, B1 => n52216, B2 => 
                           n53549, ZN => n60654);
   U3674 : AOI22_X1 port map( A1 => n52230, A2 => n53528, B1 => n52207, B2 => 
                           n52480, ZN => n60653);
   U3675 : NAND4_X1 port map( A1 => n60656, A2 => n60655, A3 => n60654, A4 => 
                           n60653, ZN => n60657);
   U3676 : AOI22_X1 port map( A1 => n60771, A2 => n60658, B1 => n60769, B2 => 
                           n60657, ZN => n60659);
   U3677 : OAI21_X1 port map( B1 => n60727, B2 => n60660, A => n60659, ZN => 
                           OUT1(5));
   U3678 : AOI22_X1 port map( A1 => n52374, A2 => n52404, B1 => n51886, B2 => 
                           n53555, ZN => n60664);
   U3679 : AOI22_X1 port map( A1 => n52081, A2 => n52413, B1 => n52380, B2 => 
                           n52410, ZN => n60663);
   U3680 : AOI22_X1 port map( A1 => n51848, A2 => n52411, B1 => n51847, B2 => 
                           n52408, ZN => n60662);
   U3681 : AOI22_X1 port map( A1 => n51869, A2 => n53533, B1 => n51846, B2 => 
                           n53537, ZN => n60661);
   U3682 : NAND4_X1 port map( A1 => n60664, A2 => n60663, A3 => n60662, A4 => 
                           n60661, ZN => n60670);
   U3683 : AOI22_X1 port map( A1 => n52378, A2 => n53554, B1 => n52077, B2 => 
                           n52406, ZN => n60668);
   U3684 : AOI22_X1 port map( A1 => n52375, A2 => n53543, B1 => n51992, B2 => 
                           n52407, ZN => n60667);
   U3685 : AOI22_X1 port map( A1 => n52114, A2 => n52417, B1 => n51849, B2 => 
                           n52403, ZN => n60666);
   U3686 : AOI22_X1 port map( A1 => n52119, A2 => n52412, B1 => n51986, B2 => 
                           n53534, ZN => n60665);
   U3687 : NAND4_X1 port map( A1 => n60668, A2 => n60667, A3 => n60666, A4 => 
                           n60665, ZN => n60669);
   U3688 : NOR2_X1 port map( A1 => n60670, A2 => n60669, ZN => n60682);
   U3689 : AOI22_X1 port map( A1 => n51944, A2 => n53528, B1 => n51959, B2 => 
                           n53540, ZN => n60674);
   U3690 : AOI22_X1 port map( A1 => n52308, A2 => n53538, B1 => n51963, B2 => 
                           n53549, ZN => n60673);
   U3691 : AOI22_X1 port map( A1 => n51939, A2 => n52402, B1 => n51945, B2 => 
                           n53541, ZN => n60672);
   U3692 : AOI22_X1 port map( A1 => n51949, A2 => n53517, B1 => n51732, B2 => 
                           n53522, ZN => n60671);
   U3693 : NAND4_X1 port map( A1 => n60674, A2 => n60673, A3 => n60672, A4 => 
                           n60671, ZN => n60680);
   U3694 : AOI22_X1 port map( A1 => n52202, A2 => n52480, B1 => n51856, B2 => 
                           n53517, ZN => n60678);
   U3695 : AOI22_X1 port map( A1 => n52239, A2 => n53546, B1 => n52212, B2 => 
                           n53524, ZN => n60677);
   U3696 : AOI22_X1 port map( A1 => n52237, A2 => n52402, B1 => n52102, B2 => 
                           n52481, ZN => n60676);
   U3697 : AOI22_X1 port map( A1 => n52250, A2 => n52479, B1 => n51831, B2 => 
                           n53538, ZN => n60675);
   U3698 : NAND4_X1 port map( A1 => n60678, A2 => n60677, A3 => n60676, A4 => 
                           n60675, ZN => n60679);
   U3699 : AOI22_X1 port map( A1 => n60771, A2 => n60680, B1 => n60769, B2 => 
                           n60679, ZN => n60681);
   U3700 : OAI21_X1 port map( B1 => n60774, B2 => n60682, A => n60681, ZN => 
                           OUT1(4));
   U3701 : AOI22_X1 port map( A1 => n52106, A2 => n53542, B1 => n51840, B2 => 
                           n53553, ZN => n60686);
   U3702 : AOI22_X1 port map( A1 => n51987, A2 => n52409, B1 => n51862, B2 => 
                           n52414, ZN => n60685);
   U3703 : AOI22_X1 port map( A1 => n51885, A2 => n52416, B1 => n52364, B2 => 
                           n52410, ZN => n60684);
   U3704 : AOI22_X1 port map( A1 => n52107, A2 => n53558, B1 => n51845, B2 => 
                           n52408, ZN => n60683);
   U3705 : NAND4_X1 port map( A1 => n60686, A2 => n60685, A3 => n60684, A4 => 
                           n60683, ZN => n60692);
   U3706 : AOI22_X1 port map( A1 => n52368, A2 => n53543, B1 => n52338, B2 => 
                           n53545, ZN => n60690);
   U3707 : AOI22_X1 port map( A1 => n51844, A2 => n52418, B1 => n52372, B2 => 
                           n53554, ZN => n60689);
   U3708 : AOI22_X1 port map( A1 => n52079, A2 => n52413, B1 => n52108, B2 => 
                           n52406, ZN => n60688);
   U3709 : AOI22_X1 port map( A1 => n51991, A2 => n52407, B1 => n51839, B2 => 
                           n52411, ZN => n60687);
   U3710 : NAND4_X1 port map( A1 => n60690, A2 => n60689, A3 => n60688, A4 => 
                           n60687, ZN => n60691);
   U3711 : NOR2_X1 port map( A1 => n60692, A2 => n60691, ZN => n60704);
   U3712 : AOI22_X1 port map( A1 => n51936, A2 => n53527, B1 => n52315, B2 => 
                           n53518, ZN => n60696);
   U3713 : AOI22_X1 port map( A1 => n51942, A2 => n53526, B1 => n51933, B2 => 
                           n52401, ZN => n60695);
   U3714 : AOI22_X1 port map( A1 => n51930, A2 => n52482, B1 => n51693, B2 => 
                           n52480, ZN => n60694);
   U3715 : AOI22_X1 port map( A1 => n51948, A2 => n52402, B1 => n51943, B2 => 
                           n53548, ZN => n60693);
   U3716 : NAND4_X1 port map( A1 => n60696, A2 => n60695, A3 => n60694, A4 => 
                           n60693, ZN => n60702);
   U3717 : AOI22_X1 port map( A1 => n52231, A2 => n53541, B1 => n52220, B2 => 
                           n53524, ZN => n60700);
   U3718 : AOI22_X1 port map( A1 => n52242, A2 => n53546, B1 => n51836, B2 => 
                           n53518, ZN => n60699);
   U3719 : AOI22_X1 port map( A1 => n52248, A2 => n52402, B1 => n52205, B2 => 
                           n53522, ZN => n60698);
   U3720 : AOI22_X1 port map( A1 => n52100, A2 => n53526, B1 => n51855, B2 => 
                           n53548, ZN => n60697);
   U3721 : NAND4_X1 port map( A1 => n60700, A2 => n60699, A3 => n60698, A4 => 
                           n60697, ZN => n60701);
   U3722 : AOI22_X1 port map( A1 => n60771, A2 => n60702, B1 => n60769, B2 => 
                           n60701, ZN => n60703);
   U3723 : OAI21_X1 port map( B1 => n60774, B2 => n60704, A => n60703, ZN => 
                           OUT1(3));
   U3724 : AOI22_X1 port map( A1 => n52384, A2 => n53545, B1 => n51838, B2 => 
                           n52416, ZN => n60708);
   U3725 : AOI22_X1 port map( A1 => n51990, A2 => n52407, B1 => n52363, B2 => 
                           n52410, ZN => n60707);
   U3726 : AOI22_X1 port map( A1 => n52075, A2 => n53558, B1 => n52103, B2 => 
                           n52406, ZN => n60706);
   U3727 : AOI22_X1 port map( A1 => n51882, A2 => n53552, B1 => n51883, B2 => 
                           n52418, ZN => n60705);
   U3728 : NAND4_X1 port map( A1 => n60708, A2 => n60707, A3 => n60706, A4 => 
                           n60705, ZN => n60714);
   U3729 : AOI22_X1 port map( A1 => n51876, A2 => n52411, B1 => n51988, B2 => 
                           n52409, ZN => n60712);
   U3730 : AOI22_X1 port map( A1 => n51880, A2 => n53533, B1 => n52082, B2 => 
                           n52417, ZN => n60711);
   U3731 : AOI22_X1 port map( A1 => n51879, A2 => n52403, B1 => n52369, B2 => 
                           n52415, ZN => n60710);
   U3732 : AOI22_X1 port map( A1 => n52116, A2 => n52413, B1 => n52376, B2 => 
                           n52405, ZN => n60709);
   U3733 : NAND4_X1 port map( A1 => n60712, A2 => n60711, A3 => n60710, A4 => 
                           n60709, ZN => n60713);
   U3734 : NOR2_X1 port map( A1 => n60714, A2 => n60713, ZN => n60726);
   U3735 : AOI22_X1 port map( A1 => n51941, A2 => n53527, B1 => n51762, B2 => 
                           n53522, ZN => n60718);
   U3736 : AOI22_X1 port map( A1 => n52310, A2 => n53538, B1 => n51957, B2 => 
                           n53548, ZN => n60717);
   U3737 : AOI22_X1 port map( A1 => n51946, A2 => n53528, B1 => n51937, B2 => 
                           n53540, ZN => n60716);
   U3738 : AOI22_X1 port map( A1 => n51947, A2 => n53539, B1 => n51955, B2 => 
                           n53549, ZN => n60715);
   U3739 : NAND4_X1 port map( A1 => n60718, A2 => n60717, A3 => n60716, A4 => 
                           n60715, ZN => n60724);
   U3740 : AOI22_X1 port map( A1 => n52228, A2 => n52402, B1 => n51854, B2 => 
                           n53517, ZN => n60722);
   U3741 : AOI22_X1 port map( A1 => n51835, A2 => n53538, B1 => n52218, B2 => 
                           n53524, ZN => n60721);
   U3742 : AOI22_X1 port map( A1 => n52099, A2 => n53540, B1 => n52210, B2 => 
                           n52480, ZN => n60720);
   U3743 : AOI22_X1 port map( A1 => n52198, A2 => n53528, B1 => n52199, B2 => 
                           n53527, ZN => n60719);
   U3744 : NAND4_X1 port map( A1 => n60722, A2 => n60721, A3 => n60720, A4 => 
                           n60719, ZN => n60723);
   U3745 : AOI22_X1 port map( A1 => n60771, A2 => n60724, B1 => n60769, B2 => 
                           n60723, ZN => n60725);
   U3746 : OAI21_X1 port map( B1 => n60727, B2 => n60726, A => n60725, ZN => 
                           OUT1(2));
   U3747 : AOI22_X1 port map( A1 => n52383, A2 => n52410, B1 => n51859, B2 => 
                           n53536, ZN => n60731);
   U3748 : AOI22_X1 port map( A1 => n51842, A2 => n53537, B1 => n51989, B2 => 
                           n53534, ZN => n60730);
   U3749 : AOI22_X1 port map( A1 => n52381, A2 => n52415, B1 => n51837, B2 => 
                           n53555, ZN => n60729);
   U3750 : AOI22_X1 port map( A1 => n52365, A2 => n53554, B1 => n52118, B2 => 
                           n52406, ZN => n60728);
   U3751 : NAND4_X1 port map( A1 => n60731, A2 => n60730, A3 => n60729, A4 => 
                           n60728, ZN => n60737);
   U3752 : AOI22_X1 port map( A1 => n51841, A2 => n52403, B1 => n51858, B2 => 
                           n53533, ZN => n60735);
   U3753 : AOI22_X1 port map( A1 => n52096, A2 => n53557, B1 => n52115, B2 => 
                           n53558, ZN => n60734);
   U3754 : AOI22_X1 port map( A1 => n52113, A2 => n52417, B1 => n51984, B2 => 
                           n53556, ZN => n60733);
   U3755 : AOI22_X1 port map( A1 => n52386, A2 => n53545, B1 => n51843, B2 => 
                           n52408, ZN => n60732);
   U3756 : NAND4_X1 port map( A1 => n60735, A2 => n60734, A3 => n60733, A4 => 
                           n60732, ZN => n60736);
   U3757 : NOR2_X1 port map( A1 => n60737, A2 => n60736, ZN => n60749);
   U3758 : AOI22_X1 port map( A1 => n51966, A2 => n53525, B1 => n52317, B2 => 
                           n53518, ZN => n60741);
   U3759 : AOI22_X1 port map( A1 => n51952, A2 => n52482, B1 => n51953, B2 => 
                           n52401, ZN => n60740);
   U3760 : AOI22_X1 port map( A1 => n51743, A2 => n52480, B1 => n51954, B2 => 
                           n53541, ZN => n60739);
   U3761 : AOI22_X1 port map( A1 => n51961, A2 => n53526, B1 => n51951, B2 => 
                           n53517, ZN => n60738);
   U3762 : NAND4_X1 port map( A1 => n60741, A2 => n60740, A3 => n60739, A4 => 
                           n60738, ZN => n60747);
   U3763 : AOI22_X1 port map( A1 => n52244, A2 => n53539, B1 => n51834, B2 => 
                           n53518, ZN => n60745);
   U3764 : AOI22_X1 port map( A1 => n52238, A2 => n52479, B1 => n51853, B2 => 
                           n53517, ZN => n60744);
   U3765 : AOI22_X1 port map( A1 => n52094, A2 => n53540, B1 => n52203, B2 => 
                           n52480, ZN => n60743);
   U3766 : AOI22_X1 port map( A1 => n52234, A2 => n53528, B1 => n52211, B2 => 
                           n53524, ZN => n60742);
   U3767 : NAND4_X1 port map( A1 => n60745, A2 => n60744, A3 => n60743, A4 => 
                           n60742, ZN => n60746);
   U3768 : AOI22_X1 port map( A1 => n60771, A2 => n60747, B1 => n60769, B2 => 
                           n60746, ZN => n60748);
   U3769 : OAI21_X1 port map( B1 => n60774, B2 => n60749, A => n60748, ZN => 
                           OUT1(1));
   U3770 : AOI22_X1 port map( A1 => n51682, A2 => n52418, B1 => n51688, B2 => 
                           n52411, ZN => n60753);
   U3771 : AOI22_X1 port map( A1 => n52101, A2 => n52417, B1 => n52367, B2 => 
                           n52415, ZN => n60752);
   U3772 : AOI22_X1 port map( A1 => n52229, A2 => n52412, B1 => n51681, B2 => 
                           n52410, ZN => n60751);
   U3773 : AOI22_X1 port map( A1 => n51684, A2 => n52416, B1 => n51827, B2 => 
                           n52408, ZN => n60750);
   U3774 : NAND4_X1 port map( A1 => n60753, A2 => n60752, A3 => n60751, A4 => 
                           n60750, ZN => n60759);
   U3775 : AOI22_X1 port map( A1 => n51685, A2 => n52409, B1 => n51689, B2 => 
                           n52414, ZN => n60757);
   U3776 : AOI22_X1 port map( A1 => n52361, A2 => n52405, B1 => n51931, B2 => 
                           n52407, ZN => n60756);
   U3777 : AOI22_X1 port map( A1 => n52227, A2 => n52413, B1 => n51686, B2 => 
                           n52403, ZN => n60755);
   U3778 : AOI22_X1 port map( A1 => n52120, A2 => n52406, B1 => n52285, B2 => 
                           n52404, ZN => n60754);
   U3779 : NAND4_X1 port map( A1 => n60757, A2 => n60756, A3 => n60755, A4 => 
                           n60754, ZN => n60758);
   U3780 : NOR2_X1 port map( A1 => n60759, A2 => n60758, ZN => n60773);
   U3781 : AOI22_X1 port map( A1 => n51683, A2 => n52480, B1 => n51979, B2 => 
                           n53548, ZN => n60763);
   U3782 : AOI22_X1 port map( A1 => n51977, A2 => n53541, B1 => n51975, B2 => 
                           n52402, ZN => n60762);
   U3783 : AOI22_X1 port map( A1 => n51973, A2 => n53528, B1 => n51932, B2 => 
                           n53549, ZN => n60761);
   U3784 : AOI22_X1 port map( A1 => n51980, A2 => n53540, B1 => n52335, B2 => 
                           n53550, ZN => n60760);
   U3785 : NAND4_X1 port map( A1 => n60763, A2 => n60762, A3 => n60761, A4 => 
                           n60760, ZN => n60770);
   U3786 : AOI22_X1 port map( A1 => n52226, A2 => n52480, B1 => n52167, B2 => 
                           n53527, ZN => n60767);
   U3787 : AOI22_X1 port map( A1 => n52165, A2 => n53539, B1 => n51687, B2 => 
                           n53550, ZN => n60766);
   U3788 : AOI22_X1 port map( A1 => n52158, A2 => n52482, B1 => n52097, B2 => 
                           n52481, ZN => n60765);
   U3789 : AOI22_X1 port map( A1 => n52166, A2 => n53528, B1 => n51690, B2 => 
                           n53548, ZN => n60764);
   U3790 : NAND4_X1 port map( A1 => n60767, A2 => n60766, A3 => n60765, A4 => 
                           n60764, ZN => n60768);
   U3791 : AOI22_X1 port map( A1 => n60771, A2 => n60770, B1 => n60769, B2 => 
                           n60768, ZN => n60772);
   U3792 : OAI21_X1 port map( B1 => n60774, B2 => n60773, A => n60772, ZN => 
                           OUT1(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_17_port, curr_instruction_to_cu_i_16_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n151, cu_i_N279, 
      cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, 
      cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_3_port, cu_i_cmd_word_6_port, 
      cu_i_cmd_word_8_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_decode_stage_dp_n44, datapath_i_decode_stage_dp_n43, 
      datapath_i_decode_stage_dp_n42, datapath_i_decode_stage_dp_n41, 
      datapath_i_decode_stage_dp_n40, datapath_i_decode_stage_dp_n39, 
      datapath_i_decode_stage_dp_n38, datapath_i_decode_stage_dp_n37, 
      datapath_i_decode_stage_dp_n36, datapath_i_decode_stage_dp_n35, 
      datapath_i_decode_stage_dp_n34, datapath_i_decode_stage_dp_n33, 
      datapath_i_decode_stage_dp_n32, datapath_i_decode_stage_dp_n31, 
      datapath_i_decode_stage_dp_n30, datapath_i_decode_stage_dp_n29, 
      datapath_i_decode_stage_dp_n28, datapath_i_decode_stage_dp_n27, 
      datapath_i_decode_stage_dp_n26, datapath_i_decode_stage_dp_n25, 
      datapath_i_decode_stage_dp_n24, datapath_i_decode_stage_dp_n23, 
      datapath_i_decode_stage_dp_n22, datapath_i_decode_stage_dp_n21, 
      datapath_i_decode_stage_dp_n20, datapath_i_decode_stage_dp_n19, 
      datapath_i_decode_stage_dp_n18, datapath_i_decode_stage_dp_n17, 
      datapath_i_decode_stage_dp_n16, datapath_i_decode_stage_dp_n15, 
      datapath_i_decode_stage_dp_n14, datapath_i_decode_stage_dp_n13, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, n302, n474, n477, n492, n1443, 
      n1445, n1447, n1449, n1453, n1613, n1614, n1615, n1617, n1619, n1621, 
      n1623, n1625, n1627, n1629, n1631, n1633, n1635, n1637, n1639, n1641, 
      n1643, n1645, n1647, n1649, n1651, n1653, n1655, n1657, n1659, n1661, 
      n1663, n1665, n1667, n1669, n1671, n1673, n2299, n5478, n5479, n3284, 
      n4052, n4060, n4128, n4337, n4417, n4953, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5388, n6772, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6808, n6809, n6810, n6811, n6812, n6813, n6814, 
      n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6823, n6835, n6836, 
      n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, 
      n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, 
      n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, 
      n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, 
      n6877, n6878, n6879, n6881, n6887, n6889, n6890, n6892, n6894, n6896, 
      n6898, n6900, n6902, n6907, n6908, n6910, n6914, n6916, n6917, n6919, 
      n6920, n6928, n6932, n6933, n6942, n6946, n6949, n6952, n6955, n6958, 
      n6961, n6964, n6967, n6970, n6973, n6976, n6979, n6982, n6985, n6988, 
      n6991, n6994, n6997, n7000, n7003, n7006, n7009, n7012, n7015, n7018, 
      n7021, n7024, n7027, n7030, n7033, n7036, n7039, n7193, n7215, n7737, 
      n7739, n7789, n7839, n7852, n7861, n7912, n8000, n8001, n8055, n9209, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_8_port, n8608, n8609, n8610, n8611, 
      n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, 
      n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, 
      n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, 
      n8642, n8643, n8645, n8646, n8647, n8648, n8649, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_27_port, n8658, n8659, n8660, n8661, n8662, n8663, n8664, 
      n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, 
      n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, 
      n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, 
      n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, 
      n8705, IRAM_ADDRESS_13_port, IRAM_ADDRESS_11_port, n8709, 
      IRAM_ADDRESS_6_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, n8714, n8715, n8716, n8717, n8718, n8719, n8720, 
      n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, 
      n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, 
      n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, 
      n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8762, 
      n8763, n8766, n8767, n8769, n8770, n8771, n8773, n8775, n8776, n8777, 
      n8778, n8779, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, 
      n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, 
      n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, 
      n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, 
      n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, 
      n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, 
      n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, 
      n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, 
      n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, 
      n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, 
      n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, 
      n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, 
      n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, 
      n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, 
      n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, 
      n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, 
      n8939, n8940, n8941, n8942, n8943, n8945, n8947, n8948, n8950, n8951, 
      n8953, n8955, n8956, n8958, n8959, n8961, n8962, n8964, n8965, n8967, 
      n8968, n8970, n8971, n8973, n8974, n8976, n8977, n8979, n8980, n8982, 
      n8983, n8985, n8986, n8988, n8989, n8991, n8993, n8994, n8995, n8996, 
      n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9006, n9008, 
      n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, 
      n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, 
      n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, 
      n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, 
      n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9067, n9068, 
      n9069, n9070, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, 
      n9081, n9082, n9083, n9084, n9085, n9086, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_7_port, n9089, n9090, IRAM_ADDRESS_9_port, n9093, n9094, 
      n9095, n9096, n9097, n9098, n9099, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9110, n9111, n9112, n9113, n9114, n9115, n9116, 
      n9117, n9118, n9119, n9120, n9121, n9122, IRAM_ADDRESS_12_port, n9141, 
      n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9152, 
      n9153, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9203, n9204, n9205, n9206, n9207, n9208, 
      n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, 
      n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
      n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, 
      n9376, n9377, n9378, n9379, n9522, n9523, n9524, n9525, n9526, n9527, 
      n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, 
      n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, 
      n9548, n9549, n9550, IRAM_ADDRESS_1_port, n9552, n9553, n9554, n9555, 
      n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, 
      n9566, n9567, n9568, n9569, n9570, n9571, IRAM_ADDRESS_0_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_30_port, n9582, 
      n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, 
      n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, 
      n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, 
      IRAM_ADDRESS_31_port, n9612, n9613, n9614, n9615, n9616, n9617, n9618, 
      n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, 
      n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, 
      n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, 
      n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, 
      n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, 
      n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, 
      n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, 
      n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, 
      n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, 
      n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, 
      n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, 
      n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, 
      n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, 
      n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, 
      n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, 
      n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, 
      n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, 
      n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, 
      n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, 
      n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, 
      n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, 
      n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, 
      n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, 
      n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, 
      n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, 
      n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, 
      n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, 
      n9889, n9890, n9891, n9892, n9893, n9894, n9895, n_3819, n_3820, n_3821, 
      n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, 
      n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, 
      n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, 
      n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, 
      n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, 
      n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, 
      n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, 
      n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, 
      n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, 
      n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, 
      n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, 
      n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, 
      n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, 
      n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, 
      n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, 
      n_3957, n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, 
      n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, 
      n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, 
      n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, 
      n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, 
      n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, 
      n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, 
      n_4020, n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, 
      n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, 
      n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, 
      n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, 
      n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, 
      n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, 
      n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, 
      n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, 
      n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, 
      n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, 
      n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, 
      n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, 
      n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, 
      n_4137, n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, 
      n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, 
      n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, 
      n_4164, n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, 
      n_4173, n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, 
      n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, 
      n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, 
      n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, 
      n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, 
      n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, 
      n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, 
      n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, 
      n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, 
      n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, 
      n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, 
      n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, 
      n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, 
      n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, 
      n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, 
      n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, 
      n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, 
      n_4326, n_4327, n_4328 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_n151);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => n6942);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n9014, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n9067, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n9067, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n9067, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n9067, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n9067, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n9067, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n9067, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n9067, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n9067, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n9067, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n9067, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n8642, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n8642, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n8642, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n8642, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n8642, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n9067, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n9014, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n9014, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n9014, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n9014, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n9014, Z 
                           => DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n9014, Z 
                           => DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n9014, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n9014, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n9014, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n9014, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n9014, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n9014, Z 
                           => DRAM_ADDRESS_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n9895, D => n9106, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n7737, D => n9201, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n7737, D => n9200, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n7737, D => n8723, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n9895, D => n8724, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n9895, D => n9105, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n9895, D => n8693, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n9895, D => n8694, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n9895, D => n8695, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n9895, D => n8696, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n9895, D => n8697, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n9895, D => n8722, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n9895, D => n8721, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n7737, D => n9099, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n7737, D => n8720, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n9895, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n9895, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n9895, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n9895, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n9895, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n9895, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n7737, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n9541, D => n9106, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n9541, D => n9201, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n9892, D => n9200, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n9541, D => n8723, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n9892, D => n8724, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n9541, D => n9105, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n9892, D => n8693, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n9892, D => n8694, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n9541, D => n8695, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n9892, D => n8696, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n9541, D => n8697, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n9892, D => n8722, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n9541, D => n8721, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n9541, D => n9099, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n9541, D => n8720, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n9541, D => n8716, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n9892, D => n8715, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n9892, D => n8714, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n9541, D => n9098, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n9892, D => n8719, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n9541, D => n8717, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n9892, D => n8698, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n9541, D => n8705, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n9892, D => n8726, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n9892, D => n8699, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n9541, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n9892, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n9892, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n9892, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n9541, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n9892, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n9892, D => n8700, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => n3284);
   clk_r_REG16834_S6 : DFFR_X1 port map( D => n5388, CK => CLK, RN => RST, Q =>
                           n_3819, QN => n9121);
   clk_r_REG16746_S3 : DFFR_X1 port map( D => n7789, CK => CLK, RN => RST, Q =>
                           n_3820, QN => n9120);
   clk_r_REG16971_S7 : DFFR_X1 port map( D => n9540, CK => CLK, RN => RST, Q =>
                           n9119, QN => n_3821);
   clk_r_REG16976_S7 : DFFR_X1 port map( D => n9545, CK => CLK, RN => RST, Q =>
                           n9118, QN => n_3822);
   clk_r_REG16975_S1 : DFFR_X1 port map( D => n9539, CK => CLK, RN => RST, Q =>
                           n9117, QN => n_3823);
   clk_r_REG16794_S2 : DFFR_X1 port map( D => n9892, CK => CLK, RN => RST, Q =>
                           n9116, QN => n_3824);
   clk_r_REG16795_S3 : DFFR_X1 port map( D => n9116, CK => CLK, RN => RST, Q =>
                           n9115, QN => n_3825);
   clk_r_REG14480_S10 : DFFS_X1 port map( D => n9571, CK => CLK, SN => RST, Q 
                           => n9114, QN => n_3826);
   clk_r_REG14584_S11 : DFFS_X1 port map( D => n9114, CK => CLK, SN => RST, Q 
                           => n9113, QN => n_3827);
   clk_r_REG14486_S8 : DFFS_X1 port map( D => n9570, CK => CLK, SN => RST, Q =>
                           n9112, QN => n_3828);
   clk_r_REG14577_S9 : DFFS_X1 port map( D => n9112, CK => CLK, SN => RST, Q =>
                           n9111, QN => n_3829);
   clk_r_REG17010_S1 : DFFR_X1 port map( D => n9547, CK => CLK, RN => RST, Q =>
                           n9110, QN => n_3830);
   clk_r_REG16734_S2 : DFFR_X1 port map( D => n9534, CK => CLK, RN => RST, Q =>
                           DRAM_READNOTWRITE, QN => n_3831);
   clk_r_REG14589_S8 : DFFS_X1 port map( D => n9569, CK => CLK, SN => RST, Q =>
                           n9108, QN => n_3832);
   clk_r_REG14594_S9 : DFFS_X1 port map( D => n9108, CK => CLK, SN => RST, Q =>
                           n9107, QN => n_3833);
   clk_r_REG16984_S7 : DFFR_X1 port map( D => n9548, CK => CLK, RN => RST, Q =>
                           n9106, QN => n9174);
   clk_r_REG16990_S7 : DFFR_X1 port map( D => n9549, CK => CLK, RN => RST, Q =>
                           n9105, QN => n_3834);
   clk_r_REG16983_S7 : DFFR_X1 port map( D => n9550, CK => CLK, RN => RST, Q =>
                           n9104, QN => n_3835);
   clk_r_REG14492_S8 : DFFS_X1 port map( D => n9568, CK => CLK, SN => RST, Q =>
                           n9103, QN => n_3836);
   clk_r_REG14570_S9 : DFFS_X1 port map( D => n9103, CK => CLK, SN => RST, Q =>
                           n9102, QN => n_3837);
   clk_r_REG16688_S2 : DFFR_X1 port map( D => n9546, CK => CLK, RN => RST, Q =>
                           n9101, QN => n_3838);
   clk_r_REG16690_S2 : DFFS_X1 port map( D => n7193, CK => CLK, SN => RST, Q =>
                           n_3839, QN => DRAM_ENABLE);
   clk_r_REG16962_S7 : DFFR_X1 port map( D => n9538, CK => CLK, RN => RST, Q =>
                           n9099, QN => n_3840);
   clk_r_REG16963_S7 : DFFR_X1 port map( D => n9537, CK => CLK, RN => RST, Q =>
                           n9098, QN => n_3841);
   clk_r_REG14499_S8 : DFFS_X1 port map( D => n9567, CK => CLK, SN => RST, Q =>
                           n9097, QN => n_3842);
   clk_r_REG14562_S9 : DFFS_X1 port map( D => n9097, CK => CLK, SN => RST, Q =>
                           n9096, QN => n_3843);
   clk_r_REG16749_S2 : DFFR_X1 port map( D => n9895, CK => CLK, RN => RST, Q =>
                           n9095, QN => n_3844);
   clk_r_REG14506_S8 : DFFS_X1 port map( D => n9566, CK => CLK, SN => RST, Q =>
                           n9094, QN => n_3845);
   clk_r_REG14554_S9 : DFFS_X1 port map( D => n9094, CK => CLK, SN => RST, Q =>
                           n9093, QN => n_3846);
   clk_r_REG17008_S4 : DFFS_X1 port map( D => n9528, CK => CLK, SN => RST, Q =>
                           n_3847, QN => n9206);
   clk_r_REG14614_S11 : DFFR_X1 port map( D => n9607, CK => CLK, RN => RST, Q 
                           => IRAM_ADDRESS_9_port, QN => n_3848);
   clk_r_REG14512_S8 : DFFS_X1 port map( D => n9565, CK => CLK, SN => RST, Q =>
                           n9090, QN => n_3849);
   clk_r_REG14547_S9 : DFFS_X1 port map( D => n9090, CK => CLK, SN => RST, Q =>
                           n9089, QN => n_3850);
   clk_r_REG14617_S11 : DFFR_X1 port map( D => n9582, CK => CLK, RN => RST, Q 
                           => IRAM_ADDRESS_7_port, QN => n_3851);
   clk_r_REG16589_S5 : DFFR_X1 port map( D => n9552, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_5_port, QN => n_3852);
   clk_r_REG14518_S8 : DFFS_X1 port map( D => n9564, CK => CLK, SN => RST, Q =>
                           n9086, QN => n_3853);
   clk_r_REG14540_S9 : DFFS_X1 port map( D => n9086, CK => CLK, SN => RST, Q =>
                           n9085, QN => n_3854);
   clk_r_REG14525_S8 : DFFS_X1 port map( D => n9563, CK => CLK, SN => RST, Q =>
                           n9084, QN => n_3855);
   clk_r_REG14533_S9 : DFFS_X1 port map( D => n9084, CK => CLK, SN => RST, Q =>
                           n9083, QN => n_3856);
   clk_r_REG14527_S8 : DFFS_X1 port map( D => n9562, CK => CLK, SN => RST, Q =>
                           n9082, QN => n_3857);
   clk_r_REG14530_S9 : DFFS_X1 port map( D => n9082, CK => CLK, SN => RST, Q =>
                           n9081, QN => n_3858);
   clk_r_REG15047_S5 : DFFR_X1 port map( D => n5478, CK => CLK, RN => RST, Q =>
                           n_3859, QN => n9152);
   clk_r_REG15043_S5 : DFFS_X1 port map( D => n7839, CK => CLK, SN => RST, Q =>
                           n_3860, QN => n9079);
   clk_r_REG13653_S4 : DFFR_X1 port map( D => n9554, CK => CLK, RN => RST, Q =>
                           n9078, QN => n_3861);
   clk_r_REG14453_S6 : DFFS_X1 port map( D => n9555, CK => CLK, SN => RST, Q =>
                           n9077, QN => n_3862);
   clk_r_REG14454_S7 : DFFS_X1 port map( D => n9077, CK => CLK, SN => RST, Q =>
                           n9076, QN => n_3863);
   clk_r_REG14616_S8 : DFFS_X1 port map( D => n9076, CK => CLK, SN => RST, Q =>
                           n9075, QN => n_3864);
   clk_r_REG16742_S2 : DFFR_X1 port map( D => n9542, CK => CLK, RN => RST, Q =>
                           n9074, QN => n_3865);
   clk_r_REG16611_S5 : DFFR_X1 port map( D => n9073, CK => CLK, RN => RST, Q =>
                           n9072, QN => n_3866);
   clk_r_REG16601_S5 : DFFR_X1 port map( D => n5479, CK => CLK, RN => RST, Q =>
                           n_3867, QN => n9153);
   clk_r_REG16593_S5 : DFFS_X1 port map( D => n7852, CK => CLK, SN => RST, Q =>
                           n_3868, QN => n9070);
   clk_r_REG14471_S7 : DFFS_X1 port map( D => n9179, CK => CLK, SN => RST, Q =>
                           n9069, QN => n_3869);
   clk_r_REG14605_S8 : DFFS_X1 port map( D => n9069, CK => CLK, SN => RST, Q =>
                           n9068, QN => n_3870);
   clk_r_REG16694_S2 : DFFS_X1 port map( D => n7193, CK => CLK, SN => RST, Q =>
                           n9067, QN => n_3871);
   clk_r_REG14593_S8 : DFFR_X1 port map( D => n1443, CK => CLK, RN => RST, Q =>
                           n_3872, QN => n9145);
   clk_r_REG14583_S10 : DFFR_X1 port map( D => n5342, CK => CLK, RN => RST, Q 
                           => n_3873, QN => n9142);
   clk_r_REG14576_S8 : DFFR_X1 port map( D => n5343, CK => CLK, RN => RST, Q =>
                           n_3874, QN => n9148);
   clk_r_REG14569_S8 : DFFR_X1 port map( D => n5344, CK => CLK, RN => RST, Q =>
                           n_3875, QN => n9150);
   clk_r_REG14561_S8 : DFFR_X1 port map( D => n5345, CK => CLK, RN => RST, Q =>
                           n_3876, QN => n9147);
   clk_r_REG14553_S8 : DFFR_X1 port map( D => n5346, CK => CLK, RN => RST, Q =>
                           n_3877, QN => n9143);
   clk_r_REG14546_S8 : DFFR_X1 port map( D => n5347, CK => CLK, RN => RST, Q =>
                           n_3878, QN => n9146);
   clk_r_REG14539_S8 : DFFR_X1 port map( D => n5348, CK => CLK, RN => RST, Q =>
                           n_3879, QN => n9149);
   clk_r_REG14532_S8 : DFFR_X1 port map( D => n5349, CK => CLK, RN => RST, Q =>
                           n_3880, QN => n9144);
   clk_r_REG14450_S7 : DFFR_X1 port map( D => n9198, CK => CLK, RN => RST, Q =>
                           n9057, QN => n_3881);
   clk_r_REG14451_S8 : DFFR_X1 port map( D => n9057, CK => CLK, RN => RST, Q =>
                           n9056, QN => n_3882);
   clk_r_REG16617_S4 : DFFS_X1 port map( D => n9195, CK => CLK, SN => RST, Q =>
                           n9055, QN => n_3883);
   clk_r_REG16610_S5 : DFFS_X1 port map( D => n9052, CK => CLK, SN => RST, Q =>
                           n9051, QN => n_3884);
   clk_r_REG16793_S2 : DFFR_X1 port map( D => n9892, CK => CLK, RN => RST, Q =>
                           n9050, QN => n_3885);
   clk_r_REG14477_S8 : DFFR_X1 port map( D => n9600, CK => CLK, RN => RST, Q =>
                           n9049, QN => n_3886);
   clk_r_REG14478_S8 : DFFS_X1 port map( D => n9600, CK => CLK, SN => RST, Q =>
                           n9048, QN => n_3887);
   clk_r_REG14484_S8 : DFFR_X1 port map( D => n9594, CK => CLK, RN => RST, Q =>
                           n9047, QN => n_3888);
   clk_r_REG14485_S8 : DFFS_X1 port map( D => n9594, CK => CLK, SN => RST, Q =>
                           n9046, QN => n_3889);
   clk_r_REG14490_S8 : DFFR_X1 port map( D => n9592, CK => CLK, RN => RST, Q =>
                           n9045, QN => n_3890);
   clk_r_REG14491_S8 : DFFS_X1 port map( D => n9592, CK => CLK, SN => RST, Q =>
                           n9044, QN => n_3891);
   clk_r_REG14496_S8 : DFFR_X1 port map( D => n9586, CK => CLK, RN => RST, Q =>
                           n9043, QN => n_3892);
   clk_r_REG14497_S8 : DFFS_X1 port map( D => n9586, CK => CLK, SN => RST, Q =>
                           n9042, QN => n_3893);
   clk_r_REG14503_S8 : DFFR_X1 port map( D => n9588, CK => CLK, RN => RST, Q =>
                           n9041, QN => n_3894);
   clk_r_REG14504_S8 : DFFS_X1 port map( D => n9588, CK => CLK, SN => RST, Q =>
                           n9040, QN => n_3895);
   clk_r_REG14510_S8 : DFFR_X1 port map( D => n9590, CK => CLK, RN => RST, Q =>
                           n9039, QN => n_3896);
   clk_r_REG14511_S8 : DFFS_X1 port map( D => n9590, CK => CLK, SN => RST, Q =>
                           n9038, QN => n_3897);
   clk_r_REG14516_S8 : DFFR_X1 port map( D => n9596, CK => CLK, RN => RST, Q =>
                           n9037, QN => n_3898);
   clk_r_REG14517_S8 : DFFS_X1 port map( D => n9596, CK => CLK, SN => RST, Q =>
                           n9036, QN => n_3899);
   clk_r_REG14522_S8 : DFFR_X1 port map( D => n9598, CK => CLK, RN => RST, Q =>
                           n9035, QN => n_3900);
   clk_r_REG14523_S8 : DFFS_X1 port map( D => n9598, CK => CLK, SN => RST, Q =>
                           n9034, QN => n_3901);
   clk_r_REG14526_S8 : DFFR_X1 port map( D => n5349, CK => CLK, RN => RST, Q =>
                           n9033, QN => n_3902);
   clk_r_REG14519_S8 : DFFR_X1 port map( D => n5348, CK => CLK, RN => RST, Q =>
                           n9032, QN => n_3903);
   clk_r_REG14513_S8 : DFFR_X1 port map( D => n5347, CK => CLK, RN => RST, Q =>
                           n9031, QN => n_3904);
   clk_r_REG14507_S8 : DFFR_X1 port map( D => n5346, CK => CLK, RN => RST, Q =>
                           n9030, QN => n_3905);
   clk_r_REG14500_S8 : DFFR_X1 port map( D => n5345, CK => CLK, RN => RST, Q =>
                           n9029, QN => n_3906);
   clk_r_REG14493_S8 : DFFR_X1 port map( D => n5344, CK => CLK, RN => RST, Q =>
                           n9028, QN => n_3907);
   clk_r_REG14487_S8 : DFFR_X1 port map( D => n5343, CK => CLK, RN => RST, Q =>
                           n9027, QN => n_3908);
   clk_r_REG14481_S10 : DFFR_X1 port map( D => n5342, CK => CLK, RN => RST, Q 
                           => n9026, QN => n_3909);
   clk_r_REG14590_S8 : DFFR_X1 port map( D => n1443, CK => CLK, RN => RST, Q =>
                           n9025, QN => n_3910);
   clk_r_REG14597_S8 : DFFR_X1 port map( D => n9602, CK => CLK, RN => RST, Q =>
                           n9024, QN => n_3911);
   clk_r_REG14598_S8 : DFFS_X1 port map( D => n9602, CK => CLK, SN => RST, Q =>
                           n9023, QN => n_3912);
   clk_r_REG16699_S3 : DFFS_X1 port map( D => n9536, CK => CLK, SN => RST, Q =>
                           n9022, QN => n_3913);
   clk_r_REG16607_S3 : DFFR_X1 port map( D => n9530, CK => CLK, RN => RST, Q =>
                           n9021, QN => n_3914);
   clk_r_REG16598_S5 : DFFS_X1 port map( D => n7852, CK => CLK, SN => RST, Q =>
                           n9020, QN => n_3915);
   clk_r_REG16599_S6 : DFFS_X1 port map( D => n9020, CK => CLK, SN => RST, Q =>
                           n9019, QN => n_3916);
   clk_r_REG16600_S7 : DFFS_X1 port map( D => n9019, CK => CLK, SN => RST, Q =>
                           n9018, QN => n_3917);
   clk_r_REG15044_S5 : DFFS_X1 port map( D => n7839, CK => CLK, SN => RST, Q =>
                           n9017, QN => n_3918);
   clk_r_REG15045_S6 : DFFS_X1 port map( D => n9017, CK => CLK, SN => RST, Q =>
                           n9016, QN => n_3919);
   clk_r_REG15046_S7 : DFFS_X1 port map( D => n9016, CK => CLK, SN => RST, Q =>
                           n9015, QN => n_3920);
   clk_r_REG16693_S2 : DFFS_X1 port map( D => n7193, CK => CLK, SN => RST, Q =>
                           n9014, QN => n_3921);
   clk_r_REG16747_S3 : DFFR_X1 port map( D => n7789, CK => CLK, RN => RST, Q =>
                           n9012, QN => n_3922);
   clk_r_REG16686_S1 : DFFS_X1 port map( D => n9182, CK => CLK, SN => RST, Q =>
                           n9011, QN => n9888);
   clk_r_REG13652_S3 : DFFR_X1 port map( D => n9170, CK => CLK, RN => RST, Q =>
                           n9010, QN => n_3923);
   clk_r_REG16754_S2 : DFFR_X1 port map( D => n9168, CK => CLK, RN => RST, Q =>
                           n_3924, QN => n9199);
   clk_r_REG16602_S3 : DFFS_X1 port map( D => n9169, CK => CLK, SN => RST, Q =>
                           n9008, QN => n_3925);
   clk_r_REG14458_S6 : DFFS_X1 port map( D => n9556, CK => CLK, SN => RST, Q =>
                           n_3926, QN => n9197);
   clk_r_REG14459_S7 : DFFR_X1 port map( D => n9197, CK => CLK, RN => RST, Q =>
                           n_3927, QN => n9006);
   clk_r_REG14448_S6 : DFFS_X1 port map( D => n9557, CK => CLK, SN => RST, Q =>
                           n_3928, QN => n9198);
   clk_r_REG14449_S7 : DFFR_X1 port map( D => n9198, CK => CLK, RN => RST, Q =>
                           n_3929, QN => n9004);
   clk_r_REG16683_S1 : DFFS_X1 port map( D => n9180, CK => CLK, SN => RST, Q =>
                           n9003, QN => n_3930);
   clk_r_REG14465_S6 : DFFS_X1 port map( D => n9178, CK => CLK, SN => RST, Q =>
                           n9002, QN => n_3931);
   clk_r_REG16752_S2 : DFFR_X1 port map( D => n8055, CK => CLK, RN => RST, Q =>
                           n9001, QN => n_3932);
   clk_r_REG17006_S4 : DFFR_X1 port map( D => n9527, CK => CLK, RN => RST, Q =>
                           n9000, QN => n_3933);
   clk_r_REG16692_S2 : DFFS_X1 port map( D => n7215, CK => CLK, SN => RST, Q =>
                           n8999, QN => n_3934);
   clk_r_REG16987_S7 : DFFR_X1 port map( D => n9603, CK => CLK, RN => RST, Q =>
                           n8998, QN => n_3935);
   clk_r_REG16989_S7 : DFFR_X1 port map( D => n9604, CK => CLK, RN => RST, Q =>
                           n8997, QN => n_3936);
   clk_r_REG16978_S7 : DFFR_X1 port map( D => n9605, CK => CLK, RN => RST, Q =>
                           n8996, QN => n_3937);
   clk_r_REG16982_S7 : DFFR_X1 port map( D => n9606, CK => CLK, RN => RST, Q =>
                           n8995, QN => n_3938);
   clk_r_REG16828_S2 : DFFR_X1 port map( D => n9892, CK => CLK, RN => RST, Q =>
                           n8994, QN => n_3939);
   clk_r_REG16614_S4 : DFFS_X1 port map( D => n9193, CK => CLK, SN => RST, Q =>
                           n8993, QN => n_3940);
   clk_r_REG16612_S3 : DFFR_X1 port map( D => n9530, CK => CLK, RN => RST, Q =>
                           n_3941, QN => n9193);
   clk_r_REG16613_S4 : DFFS_X1 port map( D => n9193, CK => CLK, SN => RST, Q =>
                           n_3942, QN => n8991);
   clk_r_REG16590_S3 : DFFR_X1 port map( D => n9170, CK => CLK, RN => RST, Q =>
                           n_3943, QN => n9194);
   clk_r_REG16591_S4 : DFFS_X1 port map( D => n9194, CK => CLK, SN => RST, Q =>
                           n_3944, QN => n8989);
   clk_r_REG16588_S7 : DFFR_X1 port map( D => n9196, CK => CLK, RN => RST, Q =>
                           n8988, QN => n_3945);
   clk_r_REG16586_S6 : DFFS_X1 port map( D => n9553, CK => CLK, SN => RST, Q =>
                           n_3946, QN => n9196);
   clk_r_REG16587_S7 : DFFR_X1 port map( D => n9196, CK => CLK, RN => RST, Q =>
                           n_3947, QN => n8986);
   clk_r_REG14462_S8 : DFFS_X1 port map( D => n9172, CK => CLK, SN => RST, Q =>
                           n8985, QN => n_3948);
   clk_r_REG14460_S7 : DFFR_X1 port map( D => n9197, CK => CLK, RN => RST, Q =>
                           n_3949, QN => n9172);
   clk_r_REG14461_S8 : DFFS_X1 port map( D => n9172, CK => CLK, SN => RST, Q =>
                           n_3950, QN => n8983);
   clk_r_REG14611_S8 : DFFS_X1 port map( D => n9192, CK => CLK, SN => RST, Q =>
                           n8982, QN => n_3951);
   clk_r_REG14609_S7 : DFFR_X1 port map( D => n9171, CK => CLK, RN => RST, Q =>
                           n_3952, QN => n9192);
   clk_r_REG14610_S8 : DFFS_X1 port map( D => n9192, CK => CLK, SN => RST, Q =>
                           n_3953, QN => n8980);
   clk_r_REG14603_S9 : DFFS_X1 port map( D => n9191, CK => CLK, SN => RST, Q =>
                           n8979, QN => n_3954);
   clk_r_REG14601_S8 : DFFR_X1 port map( D => n9601, CK => CLK, RN => RST, Q =>
                           n_3955, QN => n9191);
   clk_r_REG14602_S9 : DFFS_X1 port map( D => n9191, CK => CLK, SN => RST, Q =>
                           n_3956, QN => n8977);
   clk_r_REG14588_S9 : DFFS_X1 port map( D => n9190, CK => CLK, SN => RST, Q =>
                           n8976, QN => n_3957);
   clk_r_REG14586_S8 : DFFR_X1 port map( D => n9599, CK => CLK, RN => RST, Q =>
                           n_3958, QN => n9190);
   clk_r_REG14587_S9 : DFFS_X1 port map( D => n9190, CK => CLK, SN => RST, Q =>
                           n_3959, QN => n8974);
   clk_r_REG14582_S9 : DFFS_X1 port map( D => n9189, CK => CLK, SN => RST, Q =>
                           n8973, QN => n_3960);
   clk_r_REG14580_S8 : DFFR_X1 port map( D => n9593, CK => CLK, RN => RST, Q =>
                           n_3961, QN => n9189);
   clk_r_REG14581_S9 : DFFS_X1 port map( D => n9189, CK => CLK, SN => RST, Q =>
                           n_3962, QN => n8971);
   clk_r_REG14574_S9 : DFFS_X1 port map( D => n9188, CK => CLK, SN => RST, Q =>
                           n8970, QN => n_3963);
   clk_r_REG14572_S8 : DFFR_X1 port map( D => n9591, CK => CLK, RN => RST, Q =>
                           n_3964, QN => n9188);
   clk_r_REG14573_S9 : DFFS_X1 port map( D => n9188, CK => CLK, SN => RST, Q =>
                           n_3965, QN => n8968);
   clk_r_REG14567_S9 : DFFS_X1 port map( D => n9187, CK => CLK, SN => RST, Q =>
                           n8967, QN => n_3966);
   clk_r_REG14565_S8 : DFFR_X1 port map( D => n9585, CK => CLK, RN => RST, Q =>
                           n_3967, QN => n9187);
   clk_r_REG14566_S9 : DFFS_X1 port map( D => n9187, CK => CLK, SN => RST, Q =>
                           n_3968, QN => n8965);
   clk_r_REG14559_S9 : DFFS_X1 port map( D => n9186, CK => CLK, SN => RST, Q =>
                           n8964, QN => n_3969);
   clk_r_REG14557_S8 : DFFR_X1 port map( D => n9587, CK => CLK, RN => RST, Q =>
                           n_3970, QN => n9186);
   clk_r_REG14558_S9 : DFFS_X1 port map( D => n9186, CK => CLK, SN => RST, Q =>
                           n_3971, QN => n8962);
   clk_r_REG14551_S9 : DFFS_X1 port map( D => n9185, CK => CLK, SN => RST, Q =>
                           n8961, QN => n_3972);
   clk_r_REG14549_S8 : DFFR_X1 port map( D => n9589, CK => CLK, RN => RST, Q =>
                           n_3973, QN => n9185);
   clk_r_REG14550_S9 : DFFS_X1 port map( D => n9185, CK => CLK, SN => RST, Q =>
                           n_3974, QN => n8959);
   clk_r_REG14544_S9 : DFFS_X1 port map( D => n9184, CK => CLK, SN => RST, Q =>
                           n8958, QN => n_3975);
   clk_r_REG14542_S8 : DFFR_X1 port map( D => n9595, CK => CLK, RN => RST, Q =>
                           n_3976, QN => n9184);
   clk_r_REG14543_S9 : DFFS_X1 port map( D => n9184, CK => CLK, SN => RST, Q =>
                           n_3977, QN => n8956);
   clk_r_REG14537_S9 : DFFS_X1 port map( D => n9183, CK => CLK, SN => RST, Q =>
                           n8955, QN => n_3978);
   clk_r_REG14535_S8 : DFFR_X1 port map( D => n9597, CK => CLK, RN => RST, Q =>
                           n_3979, QN => n9183);
   clk_r_REG14536_S9 : DFFS_X1 port map( D => n9183, CK => CLK, SN => RST, Q =>
                           n_3980, QN => n8953);
   clk_r_REG16615_S3 : DFFR_X1 port map( D => n9530, CK => CLK, RN => RST, Q =>
                           n_3981, QN => n9195);
   clk_r_REG16616_S4 : DFFS_X1 port map( D => n9195, CK => CLK, SN => RST, Q =>
                           n9884, QN => n8951);
   clk_r_REG16605_S4 : DFFR_X1 port map( D => n9181, CK => CLK, RN => RST, Q =>
                           n8950, QN => n_3982);
   clk_r_REG16603_S3 : DFFS_X1 port map( D => n9169, CK => CLK, SN => RST, Q =>
                           n_3983, QN => n9181);
   clk_r_REG16604_S4 : DFFR_X1 port map( D => n9181, CK => CLK, RN => RST, Q =>
                           n_3984, QN => n8948);
   clk_r_REG16757_S4 : DFFR_X1 port map( D => n9173, CK => CLK, RN => RST, Q =>
                           n8947, QN => n_3985);
   clk_r_REG16755_S3 : DFFS_X1 port map( D => n9199, CK => CLK, SN => RST, Q =>
                           n_3986, QN => n9173);
   clk_r_REG16606_S4 : DFFR_X1 port map( D => n9181, CK => CLK, RN => RST, Q =>
                           n_3987, QN => n9886);
   clk_r_REG14442_S6 : DFFS_X1 port map( D => n9558, CK => CLK, SN => RST, Q =>
                           n8943, QN => n_3988);
   clk_r_REG14443_S7 : DFFS_X1 port map( D => n8943, CK => CLK, SN => RST, Q =>
                           n8942, QN => n_3989);
   clk_r_REG14444_S8 : DFFS_X1 port map( D => n8942, CK => CLK, SN => RST, Q =>
                           n8941, QN => n_3990);
   clk_r_REG14434_S5 : DFFS_X1 port map( D => n9561, CK => CLK, SN => RST, Q =>
                           n8940, QN => n_3991);
   clk_r_REG14435_S6 : DFFS_X1 port map( D => n8940, CK => CLK, SN => RST, Q =>
                           n8939, QN => n_3992);
   clk_r_REG14436_S7 : DFFS_X1 port map( D => n8939, CK => CLK, SN => RST, Q =>
                           n8938, QN => n_3993);
   clk_r_REG14763_S5 : DFFS_X1 port map( D => n9559, CK => CLK, SN => RST, Q =>
                           n8937, QN => n_3994);
   clk_r_REG14764_S6 : DFFS_X1 port map( D => n8937, CK => CLK, SN => RST, Q =>
                           n8936, QN => n_3995);
   clk_r_REG14765_S7 : DFFS_X1 port map( D => n8936, CK => CLK, SN => RST, Q =>
                           n8935, QN => n_3996);
   clk_r_REG14903_S5 : DFFS_X1 port map( D => n9560, CK => CLK, SN => RST, Q =>
                           n8934, QN => n_3997);
   clk_r_REG14904_S6 : DFFS_X1 port map( D => n8934, CK => CLK, SN => RST, Q =>
                           n8933, QN => n_3998);
   clk_r_REG14905_S7 : DFFS_X1 port map( D => n8933, CK => CLK, SN => RST, Q =>
                           n8932, QN => n_3999);
   clk_r_REG16964_S6 : DFFS_X1 port map( D => n9535, CK => CLK, SN => RST, Q =>
                           n8931, QN => n_4000);
   clk_r_REG13716_S3 : DFFR_X1 port map( D => n8930, CK => CLK, RN => RST, Q =>
                           n8929, QN => n_4001);
   clk_r_REG16327_S2 : DFF_X1 port map( D => n1671, CK => CLK, Q => n8928, QN 
                           => n_4002);
   clk_r_REG16328_S3 : DFFR_X1 port map( D => n8928, CK => CLK, RN => RST, Q =>
                           n8927, QN => n_4003);
   clk_r_REG13789_S2 : DFF_X1 port map( D => n1669, CK => CLK, Q => n8926, QN 
                           => n_4004);
   clk_r_REG13790_S3 : DFFR_X1 port map( D => n8926, CK => CLK, RN => RST, Q =>
                           n8925, QN => n_4005);
   clk_r_REG15752_S2 : DFF_X1 port map( D => n1667, CK => CLK, Q => n8924, QN 
                           => n_4006);
   clk_r_REG15753_S3 : DFFR_X1 port map( D => n8924, CK => CLK, RN => RST, Q =>
                           n8923, QN => n_4007);
   clk_r_REG15816_S2 : DFF_X1 port map( D => n1665, CK => CLK, Q => n8922, QN 
                           => n_4008);
   clk_r_REG15817_S3 : DFFR_X1 port map( D => n8922, CK => CLK, RN => RST, Q =>
                           n8921, QN => n_4009);
   clk_r_REG15880_S2 : DFF_X1 port map( D => n1663, CK => CLK, Q => n8920, QN 
                           => n_4010);
   clk_r_REG15881_S3 : DFFR_X1 port map( D => n8920, CK => CLK, RN => RST, Q =>
                           n8919, QN => n_4011);
   clk_r_REG15944_S2 : DFF_X1 port map( D => n1661, CK => CLK, Q => n8918, QN 
                           => n_4012);
   clk_r_REG15945_S3 : DFFR_X1 port map( D => n8918, CK => CLK, RN => RST, Q =>
                           n8917, QN => n_4013);
   clk_r_REG16008_S2 : DFF_X1 port map( D => n1659, CK => CLK, Q => n8916, QN 
                           => n_4014);
   clk_r_REG16009_S3 : DFFR_X1 port map( D => n8916, CK => CLK, RN => RST, Q =>
                           n8915, QN => n_4015);
   clk_r_REG16073_S2 : DFF_X1 port map( D => n1657, CK => CLK, Q => n8914, QN 
                           => n_4016);
   clk_r_REG16074_S3 : DFFR_X1 port map( D => n8914, CK => CLK, RN => RST, Q =>
                           n8913, QN => n_4017);
   clk_r_REG16137_S2 : DFF_X1 port map( D => n1655, CK => CLK, Q => n8912, QN 
                           => n_4018);
   clk_r_REG16138_S3 : DFFR_X1 port map( D => n8912, CK => CLK, RN => RST, Q =>
                           n8911, QN => n_4019);
   clk_r_REG16201_S2 : DFF_X1 port map( D => n1653, CK => CLK, Q => n8910, QN 
                           => n_4020);
   clk_r_REG16202_S3 : DFFR_X1 port map( D => n8910, CK => CLK, RN => RST, Q =>
                           n8909, QN => n_4021);
   clk_r_REG13831_S2 : DFF_X1 port map( D => n1651, CK => CLK, Q => n8908, QN 
                           => n_4022);
   clk_r_REG13832_S3 : DFFR_X1 port map( D => n8908, CK => CLK, RN => RST, Q =>
                           n8907, QN => n_4023);
   clk_r_REG15434_S2 : DFF_X1 port map( D => n1649, CK => CLK, Q => n8906, QN 
                           => n_4024);
   clk_r_REG15435_S3 : DFFR_X1 port map( D => n8906, CK => CLK, RN => RST, Q =>
                           n8905, QN => n_4025);
   clk_r_REG15498_S2 : DFF_X1 port map( D => n1647, CK => CLK, Q => n8904, QN 
                           => n_4026);
   clk_r_REG15499_S3 : DFFR_X1 port map( D => n8904, CK => CLK, RN => RST, Q =>
                           n8903, QN => n_4027);
   clk_r_REG15562_S2 : DFF_X1 port map( D => n1645, CK => CLK, Q => n8902, QN 
                           => n_4028);
   clk_r_REG15563_S3 : DFFR_X1 port map( D => n8902, CK => CLK, RN => RST, Q =>
                           n8901, QN => n_4029);
   clk_r_REG15626_S2 : DFF_X1 port map( D => n1643, CK => CLK, Q => n8900, QN 
                           => n_4030);
   clk_r_REG15627_S3 : DFFR_X1 port map( D => n8900, CK => CLK, RN => RST, Q =>
                           n8899, QN => n_4031);
   clk_r_REG13986_S2 : DFF_X1 port map( D => n1641, CK => CLK, Q => n8898, QN 
                           => n_4032);
   clk_r_REG13987_S3 : DFFR_X1 port map( D => n8898, CK => CLK, RN => RST, Q =>
                           n8897, QN => n_4033);
   clk_r_REG16391_S2 : DFF_X1 port map( D => n1639, CK => CLK, Q => n8896, QN 
                           => n_4034);
   clk_r_REG16392_S3 : DFFR_X1 port map( D => n8896, CK => CLK, RN => RST, Q =>
                           n8895, QN => n_4035);
   clk_r_REG16456_S2 : DFF_X1 port map( D => n1637, CK => CLK, Q => n8894, QN 
                           => n_4036);
   clk_r_REG16457_S3 : DFFR_X1 port map( D => n8894, CK => CLK, RN => RST, Q =>
                           n8893, QN => n_4037);
   clk_r_REG15114_S2 : DFF_X1 port map( D => n1635, CK => CLK, Q => n8892, QN 
                           => n_4038);
   clk_r_REG15115_S3 : DFFR_X1 port map( D => n8892, CK => CLK, RN => RST, Q =>
                           n8891, QN => n_4039);
   clk_r_REG15181_S2 : DFF_X1 port map( D => n1633, CK => CLK, Q => n8890, QN 
                           => n_4040);
   clk_r_REG15182_S3 : DFFR_X1 port map( D => n8890, CK => CLK, RN => RST, Q =>
                           n8889, QN => n_4041);
   clk_r_REG16520_S2 : DFF_X1 port map( D => n1631, CK => CLK, Q => n8888, QN 
                           => n_4042);
   clk_r_REG16521_S3 : DFFR_X1 port map( D => n8888, CK => CLK, RN => RST, Q =>
                           n8887, QN => n_4043);
   clk_r_REG15246_S2 : DFF_X1 port map( D => n1629, CK => CLK, Q => n8886, QN 
                           => n_4044);
   clk_r_REG14057_S2 : DFF_X1 port map( D => n1627, CK => CLK, Q => n8885, QN 
                           => n_4045);
   clk_r_REG14093_S2 : DFF_X1 port map( D => n1625, CK => CLK, Q => n8884, QN 
                           => n_4046);
   clk_r_REG15309_S2 : DFF_X1 port map( D => n1623, CK => CLK, Q => n8883, QN 
                           => n_4047);
   clk_r_REG14622_S2 : DFF_X1 port map( D => n1621, CK => CLK, Q => n8882, QN 
                           => n_4048);
   clk_r_REG14337_S2 : DFF_X1 port map( D => n1619, CK => CLK, Q => n8881, QN 
                           => n_4049);
   clk_r_REG14696_S2 : DFF_X1 port map( D => n1617, CK => CLK, Q => n8880, QN 
                           => n_4050);
   clk_r_REG14836_S2 : DFF_X1 port map( D => n1615, CK => CLK, Q => n8879, QN 
                           => n_4051);
   clk_r_REG14977_S2 : DFF_X1 port map( D => n1614, CK => CLK, Q => n8878, QN 
                           => n_4052);
   clk_r_REG13650_S2 : DFF_X1 port map( D => n1613, CK => CLK, Q => n8877, QN 
                           => n_4053);
   clk_r_REG13710_S2 : DFF_X1 port map( D => n7039, CK => CLK, Q => n8876, QN 
                           => n_4054);
   clk_r_REG13711_S3 : DFFR_X1 port map( D => n8876, CK => CLK, RN => RST, Q =>
                           n8875, QN => n_4055);
   clk_r_REG13712_S4 : DFFR_X1 port map( D => n8875, CK => CLK, RN => RST, Q =>
                           n8874, QN => n_4056);
   clk_r_REG13703_S2 : DFF_X1 port map( D => n7036, CK => CLK, Q => n8873, QN 
                           => n_4057);
   clk_r_REG13704_S3 : DFFR_X1 port map( D => n8873, CK => CLK, RN => RST, Q =>
                           n8872, QN => n_4058);
   clk_r_REG13705_S4 : DFFR_X1 port map( D => n8872, CK => CLK, RN => RST, Q =>
                           n8871, QN => n_4059);
   clk_r_REG13780_S2 : DFF_X1 port map( D => n7033, CK => CLK, Q => n8870, QN 
                           => n_4060);
   clk_r_REG13781_S3 : DFFR_X1 port map( D => n8870, CK => CLK, RN => RST, Q =>
                           n8869, QN => n_4061);
   clk_r_REG13782_S4 : DFFR_X1 port map( D => n8869, CK => CLK, RN => RST, Q =>
                           n8868, QN => n_4062);
   clk_r_REG13773_S2 : DFF_X1 port map( D => n7030, CK => CLK, Q => n8867, QN 
                           => n_4063);
   clk_r_REG13774_S3 : DFFR_X1 port map( D => n8867, CK => CLK, RN => RST, Q =>
                           n8866, QN => n_4064);
   clk_r_REG13775_S4 : DFFR_X1 port map( D => n8866, CK => CLK, RN => RST, Q =>
                           n8865, QN => n_4065);
   clk_r_REG13766_S2 : DFF_X1 port map( D => n7027, CK => CLK, Q => n8864, QN 
                           => n_4066);
   clk_r_REG13767_S3 : DFFR_X1 port map( D => n8864, CK => CLK, RN => RST, Q =>
                           n8863, QN => n_4067);
   clk_r_REG13768_S4 : DFFR_X1 port map( D => n8863, CK => CLK, RN => RST, Q =>
                           n8862, QN => n_4068);
   clk_r_REG13759_S2 : DFF_X1 port map( D => n7024, CK => CLK, Q => n8861, QN 
                           => n_4069);
   clk_r_REG13760_S3 : DFFR_X1 port map( D => n8861, CK => CLK, RN => RST, Q =>
                           n8860, QN => n_4070);
   clk_r_REG13761_S4 : DFFR_X1 port map( D => n8860, CK => CLK, RN => RST, Q =>
                           n8859, QN => n_4071);
   clk_r_REG13752_S2 : DFF_X1 port map( D => n7021, CK => CLK, Q => n8858, QN 
                           => n_4072);
   clk_r_REG13753_S3 : DFFR_X1 port map( D => n8858, CK => CLK, RN => RST, Q =>
                           n8857, QN => n_4073);
   clk_r_REG13754_S4 : DFFR_X1 port map( D => n8857, CK => CLK, RN => RST, Q =>
                           n8856, QN => n_4074);
   clk_r_REG13743_S2 : DFF_X1 port map( D => n7018, CK => CLK, Q => n8855, QN 
                           => n_4075);
   clk_r_REG13744_S3 : DFFR_X1 port map( D => n8855, CK => CLK, RN => RST, Q =>
                           n8854, QN => n_4076);
   clk_r_REG13745_S4 : DFFR_X1 port map( D => n8854, CK => CLK, RN => RST, Q =>
                           n8853, QN => n_4077);
   clk_r_REG13736_S1 : DFF_X1 port map( D => n7015, CK => CLK, Q => n8852, QN 
                           => n_4078);
   clk_r_REG13737_S2 : DFFR_X1 port map( D => n8852, CK => CLK, RN => RST, Q =>
                           n8851, QN => n_4079);
   clk_r_REG13738_S3 : DFFR_X1 port map( D => n8851, CK => CLK, RN => RST, Q =>
                           n8850, QN => n_4080);
   clk_r_REG13729_S1 : DFF_X1 port map( D => n7012, CK => CLK, Q => n8849, QN 
                           => n_4081);
   clk_r_REG13730_S2 : DFFR_X1 port map( D => n8849, CK => CLK, RN => RST, Q =>
                           n8848, QN => n_4082);
   clk_r_REG13731_S3 : DFFR_X1 port map( D => n8848, CK => CLK, RN => RST, Q =>
                           n8847, QN => n_4083);
   clk_r_REG13722_S1 : DFF_X1 port map( D => n7009, CK => CLK, Q => n8846, QN 
                           => n_4084);
   clk_r_REG13723_S2 : DFFR_X1 port map( D => n8846, CK => CLK, RN => RST, Q =>
                           n8845, QN => n_4085);
   clk_r_REG13724_S3 : DFFR_X1 port map( D => n8845, CK => CLK, RN => RST, Q =>
                           n8844, QN => n_4086);
   clk_r_REG13826_S1 : DFF_X1 port map( D => n7006, CK => CLK, Q => n8843, QN 
                           => n_4087);
   clk_r_REG13827_S2 : DFFR_X1 port map( D => n8843, CK => CLK, RN => RST, Q =>
                           n8842, QN => n_4088);
   clk_r_REG13828_S3 : DFFR_X1 port map( D => n8842, CK => CLK, RN => RST, Q =>
                           n8841, QN => n_4089);
   clk_r_REG13819_S1 : DFF_X1 port map( D => n7003, CK => CLK, Q => n8840, QN 
                           => n_4090);
   clk_r_REG13820_S2 : DFFR_X1 port map( D => n8840, CK => CLK, RN => RST, Q =>
                           n8839, QN => n_4091);
   clk_r_REG13821_S3 : DFFR_X1 port map( D => n8839, CK => CLK, RN => RST, Q =>
                           n8838, QN => n_4092);
   clk_r_REG13812_S1 : DFF_X1 port map( D => n7000, CK => CLK, Q => n8837, QN 
                           => n_4093);
   clk_r_REG13813_S2 : DFFR_X1 port map( D => n8837, CK => CLK, RN => RST, Q =>
                           n8836, QN => n_4094);
   clk_r_REG13814_S3 : DFFR_X1 port map( D => n8836, CK => CLK, RN => RST, Q =>
                           n8835, QN => n_4095);
   clk_r_REG13805_S1 : DFF_X1 port map( D => n6997, CK => CLK, Q => n8834, QN 
                           => n_4096);
   clk_r_REG13806_S2 : DFFR_X1 port map( D => n8834, CK => CLK, RN => RST, Q =>
                           n8833, QN => n_4097);
   clk_r_REG13807_S3 : DFFR_X1 port map( D => n8833, CK => CLK, RN => RST, Q =>
                           n8832, QN => n_4098);
   clk_r_REG13796_S1 : DFF_X1 port map( D => n6994, CK => CLK, Q => n8831, QN 
                           => n_4099);
   clk_r_REG13797_S2 : DFFR_X1 port map( D => n8831, CK => CLK, RN => RST, Q =>
                           n8830, QN => n_4100);
   clk_r_REG13798_S3 : DFFR_X1 port map( D => n8830, CK => CLK, RN => RST, Q =>
                           n8829, QN => n_4101);
   clk_r_REG13919_S1 : DFF_X1 port map( D => n6991, CK => CLK, Q => n8828, QN 
                           => n_4102);
   clk_r_REG13920_S2 : DFFR_X1 port map( D => n8828, CK => CLK, RN => RST, Q =>
                           n8827, QN => n_4103);
   clk_r_REG13921_S3 : DFFR_X1 port map( D => n8827, CK => CLK, RN => RST, Q =>
                           n8826, QN => n_4104);
   clk_r_REG13689_S1 : DFF_X1 port map( D => n6988, CK => CLK, Q => n8825, QN 
                           => n_4105);
   clk_r_REG13690_S2 : DFFR_X1 port map( D => n8825, CK => CLK, RN => RST, Q =>
                           n8824, QN => n_4106);
   clk_r_REG13691_S3 : DFFR_X1 port map( D => n8824, CK => CLK, RN => RST, Q =>
                           n8823, QN => n_4107);
   clk_r_REG13675_S1 : DFF_X1 port map( D => n6985, CK => CLK, Q => n8822, QN 
                           => n_4108);
   clk_r_REG13676_S2 : DFFR_X1 port map( D => n8822, CK => CLK, RN => RST, Q =>
                           n8821, QN => n_4109);
   clk_r_REG13677_S3 : DFFR_X1 port map( D => n8821, CK => CLK, RN => RST, Q =>
                           n8820, QN => n_4110);
   clk_r_REG13906_S1 : DFF_X1 port map( D => n6982, CK => CLK, Q => n8819, QN 
                           => n_4111);
   clk_r_REG13907_S2 : DFFR_X1 port map( D => n8819, CK => CLK, RN => RST, Q =>
                           n8818, QN => n_4112);
   clk_r_REG13908_S3 : DFFR_X1 port map( D => n8818, CK => CLK, RN => RST, Q =>
                           n8817, QN => n_4113);
   clk_r_REG13870_S2 : DFF_X1 port map( D => n6979, CK => CLK, Q => n8816, QN 
                           => n_4114);
   clk_r_REG13871_S3 : DFFR_X1 port map( D => n8816, CK => CLK, RN => RST, Q =>
                           n8815, QN => n_4115);
   clk_r_REG13872_S4 : DFFR_X1 port map( D => n8815, CK => CLK, RN => RST, Q =>
                           n8814, QN => n_4116);
   clk_r_REG13661_S2 : DFF_X1 port map( D => n6976, CK => CLK, Q => n8813, QN 
                           => n_4117);
   clk_r_REG13662_S3 : DFFR_X1 port map( D => n8813, CK => CLK, RN => RST, Q =>
                           n8812, QN => n_4118);
   clk_r_REG13663_S4 : DFFR_X1 port map( D => n8812, CK => CLK, RN => RST, Q =>
                           n8811, QN => n_4119);
   clk_r_REG13851_S2 : DFF_X1 port map( D => n6973, CK => CLK, Q => n8810, QN 
                           => n_4120);
   clk_r_REG13852_S3 : DFFR_X1 port map( D => n8810, CK => CLK, RN => RST, Q =>
                           n8809, QN => n_4121);
   clk_r_REG13853_S4 : DFFR_X1 port map( D => n8809, CK => CLK, RN => RST, Q =>
                           n8808, QN => n_4122);
   clk_r_REG14033_S2 : DFF_X1 port map( D => n6970, CK => CLK, Q => n8807, QN 
                           => n_4123);
   clk_r_REG14034_S3 : DFFR_X1 port map( D => n8807, CK => CLK, RN => RST, Q =>
                           n8806, QN => n_4124);
   clk_r_REG14035_S4 : DFFR_X1 port map( D => n8806, CK => CLK, RN => RST, Q =>
                           n8805, QN => n_4125);
   clk_r_REG14080_S1 : DFF_X1 port map( D => n6967, CK => CLK, Q => n8804, QN 
                           => n_4126);
   clk_r_REG14081_S2 : DFFR_X1 port map( D => n8804, CK => CLK, RN => RST, Q =>
                           n8803, QN => n_4127);
   clk_r_REG14082_S3 : DFFR_X1 port map( D => n8803, CK => CLK, RN => RST, Q =>
                           n8802, QN => n_4128);
   clk_r_REG13838_S1 : DFF_X1 port map( D => n6964, CK => CLK, Q => n8801, QN 
                           => n_4129);
   clk_r_REG13839_S2 : DFFR_X1 port map( D => n8801, CK => CLK, RN => RST, Q =>
                           n8800, QN => n_4130);
   clk_r_REG13840_S3 : DFFR_X1 port map( D => n8800, CK => CLK, RN => RST, Q =>
                           n8799, QN => n_4131);
   clk_r_REG14142_S1 : DFF_X1 port map( D => n6961, CK => CLK, Q => n8798, QN 
                           => n_4132);
   clk_r_REG14143_S2 : DFFR_X1 port map( D => n8798, CK => CLK, RN => RST, Q =>
                           n8797, QN => n_4133);
   clk_r_REG14144_S3 : DFFR_X1 port map( D => n8797, CK => CLK, RN => RST, Q =>
                           n8796, QN => n_4134);
   clk_r_REG14161_S1 : DFF_X1 port map( D => n6958, CK => CLK, Q => n8795, QN 
                           => n_4135);
   clk_r_REG14162_S2 : DFFR_X1 port map( D => n8795, CK => CLK, RN => RST, Q =>
                           n8794, QN => n_4136);
   clk_r_REG14163_S3 : DFFR_X1 port map( D => n8794, CK => CLK, RN => RST, Q =>
                           n8793, QN => n_4137);
   clk_r_REG14121_S1 : DFF_X1 port map( D => n6955, CK => CLK, Q => n8792, QN 
                           => n_4138);
   clk_r_REG14122_S2 : DFFR_X1 port map( D => n8792, CK => CLK, RN => RST, Q =>
                           n8791, QN => n_4139);
   clk_r_REG14123_S3 : DFFR_X1 port map( D => n8791, CK => CLK, RN => RST, Q =>
                           n8790, QN => n_4140);
   clk_r_REG14067_S1 : DFF_X1 port map( D => n6952, CK => CLK, Q => n8789, QN 
                           => n_4141);
   clk_r_REG14068_S2 : DFFR_X1 port map( D => n8789, CK => CLK, RN => RST, Q =>
                           n8788, QN => n_4142);
   clk_r_REG14069_S3 : DFFR_X1 port map( D => n8788, CK => CLK, RN => RST, Q =>
                           n8787, QN => n_4143);
   clk_r_REG14012_S1 : DFF_X1 port map( D => n6949, CK => CLK, Q => n8786, QN 
                           => n_4144);
   clk_r_REG14013_S2 : DFFR_X1 port map( D => n8786, CK => CLK, RN => RST, Q =>
                           n8785, QN => n_4145);
   clk_r_REG14014_S3 : DFFR_X1 port map( D => n8785, CK => CLK, RN => RST, Q =>
                           n8784, QN => n_4146);
   clk_r_REG13637_S1 : DFF_X1 port map( D => n6946, CK => CLK, Q => n8783, QN 
                           => n_4147);
   clk_r_REG13638_S2 : DFFR_X1 port map( D => n8783, CK => CLK, RN => RST, Q =>
                           n8782, QN => n_4148);
   clk_r_REG13639_S3 : DFFR_X1 port map( D => n8782, CK => CLK, RN => RST, Q =>
                           n8781, QN => n_4149);
   clk_r_REG17007_S4 : DFFR_X1 port map( D => n4417, CK => CLK, RN => RST, Q =>
                           n_4150, QN => n9204);
   clk_r_REG16831_S4 : DFFR_X1 port map( D => n6942, CK => CLK, RN => RST, Q =>
                           n8779, QN => n9889);
   clk_r_REG16969_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port, CK 
                           => CLK, RN => RST, Q => n8778, QN => n_4151);
   clk_r_REG16967_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port, CK 
                           => CLK, RN => RST, Q => n8777, QN => n_4152);
   clk_r_REG16968_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port, CK 
                           => CLK, RN => RST, Q => n8776, QN => n_4153);
   clk_r_REG16970_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port, CK 
                           => CLK, RN => RST, Q => n8775, QN => n_4154);
   clk_r_REG17005_S4 : DFFR_X1 port map( D => n3284, CK => CLK, RN => RST, Q =>
                           n_4155, QN => n9205);
   clk_r_REG16973_S1 : DFFS_X1 port map( D => n2299, CK => CLK, SN => RST, Q =>
                           n_4156, QN => n9207);
   clk_r_REG14474_S7 : DFFS_X1 port map( D => n7861, CK => CLK, SN => RST, Q =>
                           n8771, QN => n_4157);
   clk_r_REG16696_S2 : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => CLK, 
                           RN => RST, Q => n8770, QN => n_4158);
   clk_r_REG16753_S2 : DFFR_X1 port map( D => n9892, CK => CLK, RN => RST, Q =>
                           n_4159, QN => n8769);
   clk_r_REG16980_S7 : DFFR_X1 port map( D => n7739, CK => CLK, RN => RST, Q =>
                           n_4160, QN => n9177);
   clk_r_REG16829_S2 : DFFS_X1 port map( D => n9543, CK => CLK, SN => RST, Q =>
                           n_4161, QN => n8767);
   clk_r_REG16697_S2 : DFFR_X1 port map( D => n6933, CK => CLK, RN => RST, Q =>
                           n8766, QN => n_4162);
   clk_r_REG16981_S7 : DFFS_X1 port map( D => n474, CK => CLK, SN => RST, Q => 
                           n_4163, QN => n9175);
   clk_r_REG16830_S2 : DFFS_X1 port map( D => n6928, CK => CLK, SN => RST, Q =>
                           n8763, QN => n_4164);
   clk_r_REG16966_S1 : DFFS_X1 port map( D => n477, CK => CLK, SN => RST, Q => 
                           n8762, QN => n_4165);
   clk_r_REG14470_S6 : DFFR_X1 port map( D => n7912, CK => CLK, RN => RST, Q =>
                           n9885, QN => n9179);
   clk_r_REG14607_S6 : DFFS_X1 port map( D => n4128, CK => CLK, SN => RST, Q =>
                           n_4166, QN => n9171);
   clk_r_REG14608_S7 : DFFR_X1 port map( D => n9171, CK => CLK, RN => RST, Q =>
                           n_4167, QN => n8759);
   clk_r_REG14595_S8 : DFFR_X1 port map( D => n9601, CK => CLK, RN => RST, Q =>
                           n_4168, QN => n8758);
   clk_r_REG14475_S8 : DFFR_X1 port map( D => n9599, CK => CLK, RN => RST, Q =>
                           n_4169, QN => n8757);
   clk_r_REG14520_S8 : DFFR_X1 port map( D => n9597, CK => CLK, RN => RST, Q =>
                           n_4170, QN => n8756);
   clk_r_REG14514_S8 : DFFR_X1 port map( D => n9595, CK => CLK, RN => RST, Q =>
                           n_4171, QN => n8755);
   clk_r_REG14482_S8 : DFFR_X1 port map( D => n9593, CK => CLK, RN => RST, Q =>
                           n_4172, QN => n8754);
   clk_r_REG14488_S8 : DFFR_X1 port map( D => n9591, CK => CLK, RN => RST, Q =>
                           n_4173, QN => n8753);
   clk_r_REG14508_S8 : DFFR_X1 port map( D => n9589, CK => CLK, RN => RST, Q =>
                           n_4174, QN => n8752);
   clk_r_REG14501_S8 : DFFR_X1 port map( D => n9587, CK => CLK, RN => RST, Q =>
                           n_4175, QN => n8751);
   clk_r_REG14494_S8 : DFFR_X1 port map( D => n9585, CK => CLK, RN => RST, Q =>
                           n_4176, QN => n8750);
   clk_r_REG14464_S6 : DFFR_X1 port map( D => n9178, CK => CLK, RN => RST, Q =>
                           n_4177, QN => n8749);
   clk_r_REG14466_S7 : DFFS_X1 port map( D => n8749, CK => CLK, SN => RST, Q =>
                           n8748, QN => n_4178);
   clk_r_REG14613_S8 : DFFS_X1 port map( D => n8748, CK => CLK, SN => RST, Q =>
                           n8747, QN => n_4179);
   clk_r_REG14447_S6 : DFFS_X1 port map( D => n9557, CK => CLK, SN => RST, Q =>
                           n_4180, QN => n8746);
   clk_r_REG16685_S1 : DFFS_X1 port map( D => n9182, CK => CLK, SN => RST, Q =>
                           n9882, QN => n8745);
   clk_r_REG14457_S6 : DFFS_X1 port map( D => n9556, CK => CLK, SN => RST, Q =>
                           n_4181, QN => n8744);
   clk_r_REG16744_S2 : DFFR_X1 port map( D => n6919, CK => CLK, RN => RST, Q =>
                           n8743, QN => n_4182);
   clk_r_REG16743_S2 : DFFS_X1 port map( D => n6920, CK => CLK, SN => RST, Q =>
                           n8742, QN => n_4183);
   clk_r_REG14472_S7 : DFFS_X1 port map( D => n6917, CK => CLK, SN => RST, Q =>
                           n8741, QN => n_4184);
   clk_r_REG14473_S7 : DFFR_X1 port map( D => n6916, CK => CLK, RN => RST, Q =>
                           n8740, QN => n_4185);
   clk_r_REG14438_S6 : DFFS_X1 port map( D => n9558, CK => CLK, SN => RST, Q =>
                           n_4186, QN => n8739);
   clk_r_REG14433_S5 : DFFS_X1 port map( D => n9561, CK => CLK, SN => RST, Q =>
                           n_4187, QN => n8738);
   clk_r_REG17009_S1 : DFFS_X1 port map( D => n6914, CK => CLK, SN => RST, Q =>
                           n8737, QN => n_4188);
   clk_r_REG14468_S5 : DFFS_X1 port map( D => n6910, CK => CLK, SN => RST, Q =>
                           n8736, QN => n_4189);
   clk_r_REG14599_S5 : DFFR_X1 port map( D => n8001, CK => CLK, RN => RST, Q =>
                           n8735, QN => n_4190);
   clk_r_REG14591_S8 : DFFS_X1 port map( D => n8000, CK => CLK, SN => RST, Q =>
                           n8734, QN => n_4191);
   clk_r_REG16985_S7 : DFFR_X1 port map( D => n6932, CK => CLK, RN => RST, Q =>
                           n8733, QN => n_4192);
   clk_r_REG16992_S7 : DFFS_X1 port map( D => n492, CK => CLK, SN => RST, Q => 
                           n8732, QN => n_4193);
   clk_r_REG14529_S9 : DFFS_X1 port map( D => n6908, CK => CLK, SN => RST, Q =>
                           n8731, QN => n_4194);
   clk_r_REG13651_S2 : DFF_X1 port map( D => n6907, CK => CLK, Q => n8730, QN 
                           => n_4195);
   clk_r_REG14762_S5 : DFFS_X1 port map( D => n9559, CK => CLK, SN => RST, Q =>
                           n_4196, QN => n8729);
   clk_r_REG16682_S1 : DFFS_X1 port map( D => n9180, CK => CLK, SN => RST, Q =>
                           n_4197, QN => n8728);
   clk_r_REG16684_S2 : DFFR_X1 port map( D => n8728, CK => CLK, RN => RST, Q =>
                           n8727, QN => n_4198);
   clk_r_REG16836_S7 : DFFR_X1 port map( D => n6881, CK => CLK, RN => RST, Q =>
                           n8726, QN => n_4199);
   clk_r_REG16965_S1 : DFFR_X1 port map( D => n9544, CK => CLK, RN => RST, Q =>
                           n_4200, QN => n8725);
   clk_r_REG16991_S7 : DFFR_X1 port map( D => n6900, CK => CLK, RN => RST, Q =>
                           n8724, QN => n9203);
   clk_r_REG16993_S7 : DFFR_X1 port map( D => n6898, CK => CLK, RN => RST, Q =>
                           n8723, QN => n_4201);
   clk_r_REG16994_S7 : DFFR_X1 port map( D => n6889, CK => CLK, RN => RST, Q =>
                           n8722, QN => n_4202);
   clk_r_REG16893_S7 : DFFR_X1 port map( D => n6892, CK => CLK, RN => RST, Q =>
                           n8721, QN => n_4203);
   clk_r_REG16894_S7 : DFFR_X1 port map( D => n6890, CK => CLK, RN => RST, Q =>
                           n8720, QN => n_4204);
   clk_r_REG16895_S7 : DFFS_X1 port map( D => n9583, CK => CLK, SN => RST, Q =>
                           n_4205, QN => n8719);
   clk_r_REG16832_S4 : DFFS_X1 port map( D => n6894, CK => CLK, SN => RST, Q =>
                           n8718, QN => n_4206);
   clk_r_REG16930_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_20_port,
                           CK => CLK, RN => RST, Q => n8717, QN => n_4207);
   clk_r_REG16933_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_16_port,
                           CK => CLK, RN => RST, Q => n8715, QN => n_4208);
   clk_r_REG16958_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_17_port,
                           CK => CLK, RN => RST, Q => n8714, QN => n_4209);
   clk_r_REG14901_S5 : DFFS_X1 port map( D => n9584, CK => CLK, SN => RST, Q =>
                           n_4210, QN => IRAM_ADDRESS_2_port);
   clk_r_REG14761_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_4211);
   clk_r_REG14431_S4 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_4212);
   clk_r_REG14445_S9 : DFFR_X1 port map( D => n1453, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_6_port, QN => n_4213);
   clk_r_REG16741_S2 : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK => CLK, 
                           RN => RST, Q => n8709, QN => n_4214);
   clk_r_REG16740_S2 : DFFR_X1 port map( D => n9526, CK => CLK, RN => RST, Q =>
                           n_4215, QN => IRAM_ENABLE);
   clk_r_REG14612_S7 : DFFS_X1 port map( D => n9608, CK => CLK, SN => RST, Q =>
                           n_4216, QN => IRAM_ADDRESS_11_port);
   clk_r_REG14596_S8 : DFFS_X1 port map( D => n9602, CK => CLK, SN => RST, Q =>
                           n_4217, QN => IRAM_ADDRESS_13_port);
   clk_r_REG16959_S7 : DFFR_X1 port map( D => n6902, CK => CLK, RN => RST, Q =>
                           n8705, QN => n_4218);
   clk_r_REG16736_S2 : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK => CLK, 
                           RN => RST, Q => n8704, QN => n_4219);
   clk_r_REG16735_S3 : DFFR_X1 port map( D => n6879, CK => CLK, RN => RST, Q =>
                           n8703, QN => n_4220);
   clk_r_REG16695_S3 : DFFR_X1 port map( D => n6878, CK => CLK, RN => RST, Q =>
                           n8702, QN => n_4221);
   clk_r_REG16791_S2 : DFFR_X1 port map( D => n6877, CK => CLK, RN => RST, Q =>
                           n8701, QN => n_4222);
   clk_r_REG16995_S7 : DFFR_X1 port map( D => n6876, CK => CLK, RN => RST, Q =>
                           n8700, QN => n_4223);
   clk_r_REG16997_S7 : DFFR_X1 port map( D => n6875, CK => CLK, RN => RST, Q =>
                           n8699, QN => n_4224);
   clk_r_REG16960_S7 : DFFR_X1 port map( D => n6874, CK => CLK, RN => RST, Q =>
                           n8698, QN => n_4225);
   clk_r_REG17000_S7 : DFFR_X1 port map( D => n6873, CK => CLK, RN => RST, Q =>
                           n8697, QN => n_4226);
   clk_r_REG17001_S7 : DFFR_X1 port map( D => n6872, CK => CLK, RN => RST, Q =>
                           n8696, QN => n_4227);
   clk_r_REG17002_S7 : DFFR_X1 port map( D => n6871, CK => CLK, RN => RST, Q =>
                           n8695, QN => n_4228);
   clk_r_REG17003_S7 : DFFR_X1 port map( D => n6870, CK => CLK, RN => RST, Q =>
                           n8694, QN => n_4229);
   clk_r_REG17004_S7 : DFFR_X1 port map( D => n6869, CK => CLK, RN => RST, Q =>
                           n8693, QN => n_4230);
   clk_r_REG16796_S3 : DFFR_X1 port map( D => n6868, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8692, QN => n_4231);
   clk_r_REG16797_S3 : DFFR_X1 port map( D => n6867, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8691, QN => n_4232);
   clk_r_REG16815_S3 : DFFR_X1 port map( D => n6866, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8690, QN => n_4233);
   clk_r_REG16816_S3 : DFFR_X1 port map( D => n6865, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8689, QN => n_4234);
   clk_r_REG16798_S3 : DFFR_X1 port map( D => n6864, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8688, QN => n_4235);
   clk_r_REG16799_S3 : DFFR_X1 port map( D => n6863, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8687, QN => n_4236);
   clk_r_REG16817_S3 : DFFR_X1 port map( D => n6862, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8686, QN => n_4237);
   clk_r_REG16818_S3 : DFFR_X1 port map( D => n6861, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8685, QN => n_4238);
   clk_r_REG16800_S3 : DFFR_X1 port map( D => n6860, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8684, QN => n_4239);
   clk_r_REG16801_S3 : DFFR_X1 port map( D => n6859, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8683, QN => n_4240);
   clk_r_REG16819_S3 : DFFR_X1 port map( D => n6858, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8682, QN => n_4241);
   clk_r_REG16820_S3 : DFFR_X1 port map( D => n6857, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8681, QN => n_4242);
   clk_r_REG16802_S3 : DFFR_X1 port map( D => n6856, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8680, QN => n_4243);
   clk_r_REG16803_S3 : DFFR_X1 port map( D => n6855, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8679, QN => n_4244);
   clk_r_REG16821_S3 : DFFR_X1 port map( D => n6854, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8678, QN => n_4245);
   clk_r_REG16822_S3 : DFFR_X1 port map( D => n6853, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8677, QN => n_4246);
   clk_r_REG16804_S3 : DFFR_X1 port map( D => n6852, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8676, QN => n_4247);
   clk_r_REG16805_S3 : DFFR_X1 port map( D => n6851, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8675, QN => n_4248);
   clk_r_REG16823_S3 : DFFR_X1 port map( D => n6850, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8674, QN => n_4249);
   clk_r_REG16824_S3 : DFFR_X1 port map( D => n6849, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8673, QN => n_4250);
   clk_r_REG16806_S3 : DFFR_X1 port map( D => n6848, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8672, QN => n_4251);
   clk_r_REG16807_S3 : DFFR_X1 port map( D => n6847, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8671, QN => n_4252);
   clk_r_REG16825_S3 : DFFR_X1 port map( D => n6846, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8670, QN => n_4253);
   clk_r_REG16826_S3 : DFFR_X1 port map( D => n6845, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8669, QN => n_4254);
   clk_r_REG16808_S3 : DFFR_X1 port map( D => n6844, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8668, QN => n_4255);
   clk_r_REG16809_S3 : DFFR_X1 port map( D => n6843, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8667, QN => n_4256);
   clk_r_REG16827_S3 : DFFR_X1 port map( D => n6842, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8666, QN => n_4257);
   clk_r_REG16810_S3 : DFFR_X1 port map( D => n6841, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8665, QN => n_4258);
   clk_r_REG16811_S3 : DFFR_X1 port map( D => n6840, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8664, QN => n_4259);
   clk_r_REG16812_S3 : DFFR_X1 port map( D => n6839, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8663, QN => n_4260);
   clk_r_REG16813_S3 : DFFR_X1 port map( D => n6838, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8662, QN => n_4261);
   clk_r_REG16814_S3 : DFFR_X1 port map( D => n6837, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n8661, QN => n_4262);
   clk_r_REG16792_S3 : DFFR_X1 port map( D => n6836, CK => CLK, RN => RST, Q =>
                           n8660, QN => n_4263);
   clk_r_REG16972_S1 : DFFS_X1 port map( D => n6790, CK => CLK, SN => RST, Q =>
                           n8659, QN => n_4264);
   clk_r_REG16700_S4 : DFFS_X1 port map( D => n6835, CK => CLK, SN => RST, Q =>
                           n8658, QN => n_4265);
   clk_r_REG14515_S8 : DFFS_X1 port map( D => n9596, CK => CLK, SN => RST, Q =>
                           n_4266, QN => IRAM_ADDRESS_27_port);
   clk_r_REG14521_S8 : DFFS_X1 port map( D => n9598, CK => CLK, SN => RST, Q =>
                           n_4267, QN => IRAM_ADDRESS_29_port);
   clk_r_REG14509_S8 : DFFS_X1 port map( D => n9590, CK => CLK, SN => RST, Q =>
                           n_4268, QN => IRAM_ADDRESS_25_port);
   clk_r_REG14502_S8 : DFFS_X1 port map( D => n9588, CK => CLK, SN => RST, Q =>
                           n_4269, QN => IRAM_ADDRESS_23_port);
   clk_r_REG14483_S8 : DFFS_X1 port map( D => n9594, CK => CLK, SN => RST, Q =>
                           n_4270, QN => IRAM_ADDRESS_17_port);
   clk_r_REG14495_S8 : DFFS_X1 port map( D => n9586, CK => CLK, SN => RST, Q =>
                           n_4271, QN => IRAM_ADDRESS_21_port);
   clk_r_REG14489_S8 : DFFS_X1 port map( D => n9592, CK => CLK, SN => RST, Q =>
                           n_4272, QN => IRAM_ADDRESS_19_port);
   clk_r_REG14476_S8 : DFFS_X1 port map( D => n9600, CK => CLK, SN => RST, Q =>
                           n_4273, QN => IRAM_ADDRESS_15_port);
   clk_r_REG16698_S3 : DFFS_X1 port map( D => n9536, CK => CLK, SN => RST, Q =>
                           n_4274, QN => n8649);
   clk_r_REG16977_S7 : DFFR_X1 port map( D => n9605, CK => CLK, RN => RST, Q =>
                           n9890, QN => n8648);
   clk_r_REG16979_S7 : DFFR_X1 port map( D => n9606, CK => CLK, RN => RST, Q =>
                           n_4275, QN => n8647);
   clk_r_REG16986_S7 : DFFR_X1 port map( D => n9603, CK => CLK, RN => RST, Q =>
                           n9201, QN => n8646);
   clk_r_REG16988_S7 : DFFR_X1 port map( D => n9604, CK => CLK, RN => RST, Q =>
                           n9200, QN => n8645);
   clk_r_REG16974_S1 : DFFR_X1 port map( D => n4060, CK => CLK, RN => RST, Q =>
                           n_4276, QN => n9208);
   clk_r_REG16680_S1 : DFFR_X1 port map( D => n6896, CK => CLK, RN => RST, Q =>
                           n8643, QN => n_4277);
   clk_r_REG16689_S2 : DFFR_X1 port map( D => n9533, CK => CLK, RN => RST, Q =>
                           n_4278, QN => n8642);
   clk_r_REG16681_S1 : DFFR_X1 port map( D => n4052, CK => CLK, RN => RST, Q =>
                           n8641, QN => n_4279);
   clk_r_REG14615_S6 : DFFS_X1 port map( D => n6823, CK => CLK, SN => RST, Q =>
                           n8640, QN => n_4280);
   clk_r_REG14446_S5 : DFFR_X1 port map( D => n6821, CK => CLK, RN => RST, Q =>
                           n8639, QN => n_4281);
   clk_r_REG13654_S5 : DFFR_X1 port map( D => n6820, CK => CLK, RN => RST, Q =>
                           n8638, QN => n_4282);
   clk_r_REG14456_S5 : DFFR_X1 port map( D => n6819, CK => CLK, RN => RST, Q =>
                           n8637, QN => n_4283);
   clk_r_REG14606_S5 : DFFR_X1 port map( D => n6818, CK => CLK, RN => RST, Q =>
                           n8636, QN => n_4284);
   clk_r_REG14600_S6 : DFFR_X1 port map( D => n6817, CK => CLK, RN => RST, Q =>
                           n8635, QN => n_4285);
   clk_r_REG14585_S9 : DFFR_X1 port map( D => n6816, CK => CLK, RN => RST, Q =>
                           n8634, QN => n_4286);
   clk_r_REG14578_S9 : DFFR_X1 port map( D => n6815, CK => CLK, RN => RST, Q =>
                           n8633, QN => n_4287);
   clk_r_REG14571_S9 : DFFR_X1 port map( D => n6814, CK => CLK, RN => RST, Q =>
                           n8632, QN => n_4288);
   clk_r_REG14563_S9 : DFFR_X1 port map( D => n6813, CK => CLK, RN => RST, Q =>
                           n8631, QN => n_4289);
   clk_r_REG14555_S9 : DFFR_X1 port map( D => n6812, CK => CLK, RN => RST, Q =>
                           n8630, QN => n_4290);
   clk_r_REG14548_S9 : DFFR_X1 port map( D => n6811, CK => CLK, RN => RST, Q =>
                           n8629, QN => n_4291);
   clk_r_REG14541_S9 : DFFR_X1 port map( D => n6810, CK => CLK, RN => RST, Q =>
                           n8628, QN => n_4292);
   clk_r_REG14534_S9 : DFFR_X1 port map( D => n6809, CK => CLK, RN => RST, Q =>
                           n8627, QN => n_4293);
   clk_r_REG14766_S5 : DFFS_X1 port map( D => n6806, CK => CLK, SN => RST, Q =>
                           n8625, QN => n_4294);
   clk_r_REG14432_S4 : DFFS_X1 port map( D => n6805, CK => CLK, SN => RST, Q =>
                           n8624, QN => n_4295);
   clk_r_REG14437_S5 : DFFS_X1 port map( D => n6804, CK => CLK, SN => RST, Q =>
                           n8623, QN => n_4296);
   clk_r_REG14452_S5 : DFFS_X1 port map( D => n6803, CK => CLK, SN => RST, Q =>
                           n8622, QN => n_4297);
   clk_r_REG14463_S5 : DFFS_X1 port map( D => n6802, CK => CLK, SN => RST, Q =>
                           n8621, QN => n_4298);
   clk_r_REG14469_S5 : DFFS_X1 port map( D => n6801, CK => CLK, SN => RST, Q =>
                           n8620, QN => n_4299);
   clk_r_REG14592_S9 : DFFS_X1 port map( D => n6800, CK => CLK, SN => RST, Q =>
                           n8619, QN => n_4300);
   clk_r_REG14479_S9 : DFFS_X1 port map( D => n6799, CK => CLK, SN => RST, Q =>
                           n8618, QN => n_4301);
   clk_r_REG14575_S9 : DFFS_X1 port map( D => n6798, CK => CLK, SN => RST, Q =>
                           n8617, QN => n_4302);
   clk_r_REG14568_S9 : DFFS_X1 port map( D => n6797, CK => CLK, SN => RST, Q =>
                           n8616, QN => n_4303);
   clk_r_REG14560_S9 : DFFS_X1 port map( D => n6796, CK => CLK, SN => RST, Q =>
                           n8615, QN => n_4304);
   clk_r_REG14552_S9 : DFFS_X1 port map( D => n6795, CK => CLK, SN => RST, Q =>
                           n8614, QN => n_4305);
   clk_r_REG14545_S9 : DFFS_X1 port map( D => n6794, CK => CLK, SN => RST, Q =>
                           n8613, QN => n_4306);
   clk_r_REG14538_S9 : DFFS_X1 port map( D => n6793, CK => CLK, SN => RST, Q =>
                           n8612, QN => n_4307);
   clk_r_REG14531_S9 : DFFS_X1 port map( D => n6792, CK => CLK, SN => RST, Q =>
                           n8611, QN => n_4308);
   clk_r_REG14906_S5 : DFFR_X1 port map( D => n6791, CK => CLK, RN => RST, Q =>
                           n8610, QN => n_4309);
   clk_r_REG14902_S5 : DFFS_X1 port map( D => n9560, CK => CLK, SN => RST, Q =>
                           n_4310, QN => n8609);
   clk_r_REG16790_S1 : DFFR_X1 port map( D => n302, CK => CLK, RN => RST, Q => 
                           n8608, QN => n_4311);
   clk_r_REG14455_S7 : DFFR_X1 port map( D => n1449, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_8_port, QN => n_4312);
   clk_r_REG14467_S7 : DFFR_X1 port map( D => n1447, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_10_port, QN => n_4313);
   clk_r_REG14528_S8 : DFFR_X1 port map( D => n6772, CK => CLK, RN => RST, Q =>
                           n9209, QN => n_4314);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => n9525, ADD_WR(3) => n9522, ADD_WR(2) =>
                           n4953, ADD_WR(1) => n9523, ADD_WR(0) => n9524, 
                           ADD_RD1(4) => n6876, ADD_RD1(3) => n6875, ADD_RD1(2)
                           => n6881, ADD_RD1(1) => n6902, ADD_RD1(0) => n6874, 
                           ADD_RD2(4) => curr_instruction_to_cu_i_20_port, 
                           ADD_RD2(3) => curr_instruction_to_cu_i_19_port, 
                           ADD_RD2(2) => n9537, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n43, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n44, OUT1(31) => n1673, 
                           OUT1(30) => n1671, OUT1(29) => n1669, OUT1(28) => 
                           n1667, OUT1(27) => n1665, OUT1(26) => n1663, 
                           OUT1(25) => n1661, OUT1(24) => n1659, OUT1(23) => 
                           n1657, OUT1(22) => n1655, OUT1(21) => n1653, 
                           OUT1(20) => n1651, OUT1(19) => n1649, OUT1(18) => 
                           n1647, OUT1(17) => n1645, OUT1(16) => n1643, 
                           OUT1(15) => n1641, OUT1(14) => n1639, OUT1(13) => 
                           n1637, OUT1(12) => n1635, OUT1(11) => n1633, 
                           OUT1(10) => n1631, OUT1(9) => n1629, OUT1(8) => 
                           n1627, OUT1(7) => n1625, OUT1(6) => n1623, OUT1(5) 
                           => n1621, OUT1(4) => n1619, OUT1(3) => n1617, 
                           OUT1(2) => n1615, OUT1(1) => n1614, OUT1(0) => n1613
                           , OUT2(31) => n7039, OUT2(30) => n7036, OUT2(29) => 
                           n7033, OUT2(28) => n7030, OUT2(27) => n7027, 
                           OUT2(26) => n7024, OUT2(25) => n7021, OUT2(24) => 
                           n7018, OUT2(23) => n7015, OUT2(22) => n7012, 
                           OUT2(21) => n7009, OUT2(20) => n7006, OUT2(19) => 
                           n7003, OUT2(18) => n7000, OUT2(17) => n6997, 
                           OUT2(16) => n6994, OUT2(15) => n6991, OUT2(14) => 
                           n6988, OUT2(13) => n6985, OUT2(12) => n6982, 
                           OUT2(11) => n6979, OUT2(10) => n6976, OUT2(9) => 
                           n6973, OUT2(8) => n6970, OUT2(7) => n6967, OUT2(6) 
                           => n6964, OUT2(5) => n6961, OUT2(4) => n6958, 
                           OUT2(3) => n6955, OUT2(2) => n6952, OUT2(1) => n6949
                           , OUT2(0) => n6946, RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_4315, mul_exeception => 
                           n_4316, FUNC(0) => n9529, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_4317, 
                           OUTALU(31) => datapath_i_alu_output_val_i_31_port, 
                           OUTALU(30) => datapath_i_alu_output_val_i_30_port, 
                           OUTALU(29) => datapath_i_alu_output_val_i_29_port, 
                           OUTALU(28) => datapath_i_alu_output_val_i_28_port, 
                           OUTALU(27) => datapath_i_alu_output_val_i_27_port, 
                           OUTALU(26) => datapath_i_alu_output_val_i_26_port, 
                           OUTALU(25) => datapath_i_alu_output_val_i_25_port, 
                           OUTALU(24) => datapath_i_alu_output_val_i_24_port, 
                           OUTALU(23) => datapath_i_alu_output_val_i_23_port, 
                           OUTALU(22) => datapath_i_alu_output_val_i_22_port, 
                           OUTALU(21) => datapath_i_alu_output_val_i_21_port, 
                           OUTALU(20) => datapath_i_alu_output_val_i_20_port, 
                           OUTALU(19) => datapath_i_alu_output_val_i_19_port, 
                           OUTALU(18) => datapath_i_alu_output_val_i_18_port, 
                           OUTALU(17) => datapath_i_alu_output_val_i_17_port, 
                           OUTALU(16) => datapath_i_alu_output_val_i_16_port, 
                           OUTALU(15) => datapath_i_alu_output_val_i_15_port, 
                           OUTALU(14) => datapath_i_alu_output_val_i_14_port, 
                           OUTALU(13) => datapath_i_alu_output_val_i_13_port, 
                           OUTALU(12) => datapath_i_alu_output_val_i_12_port, 
                           OUTALU(11) => datapath_i_alu_output_val_i_11_port, 
                           OUTALU(10) => datapath_i_alu_output_val_i_10_port, 
                           OUTALU(9) => datapath_i_alu_output_val_i_9_port, 
                           OUTALU(8) => datapath_i_alu_output_val_i_8_port, 
                           OUTALU(7) => datapath_i_alu_output_val_i_7_port, 
                           OUTALU(6) => datapath_i_alu_output_val_i_6_port, 
                           OUTALU(5) => datapath_i_alu_output_val_i_5_port, 
                           OUTALU(4) => datapath_i_alu_output_val_i_4_port, 
                           OUTALU(3) => datapath_i_alu_output_val_i_3_port, 
                           OUTALU(2) => datapath_i_alu_output_val_i_2_port, 
                           OUTALU(1) => datapath_i_alu_output_val_i_1_port, 
                           OUTALU(0) => datapath_i_alu_output_val_i_0_port, 
                           rst_BAR => RST);
   U3692 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_31_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(31), ZN => n9346
                           );
   U3694 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_30_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(30), ZN => n9347
                           );
   U3696 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_29_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(29), ZN => n9348
                           );
   U3698 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_28_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(28), ZN => n9349
                           );
   U3700 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_27_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(27), ZN => n9350
                           );
   U3702 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_26_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(26), ZN => n9351
                           );
   U3704 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_25_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(25), ZN => n9352
                           );
   U3706 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_24_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(24), ZN => n9353
                           );
   U3708 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_23_port, A2 => 
                           n9893, B1 => n9894, B2 => DRAM_DATA(23), ZN => n9354
                           );
   U3710 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(22), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_22_port, ZN => n9355)
                           ;
   U3712 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(21), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_21_port, ZN => n9356)
                           ;
   U3714 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(20), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_20_port, ZN => n9357)
                           ;
   U3716 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(19), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_19_port, ZN => n9358)
                           ;
   U3718 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(18), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_18_port, ZN => n9359)
                           ;
   U3720 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(17), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_17_port, ZN => n9360)
                           ;
   U3722 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(16), B1 => n9378, B2
                           => datapath_i_alu_output_val_i_16_port, ZN => n9361)
                           ;
   U3724 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(15), B1 => n9893, B2
                           => datapath_i_alu_output_val_i_15_port, ZN => n9362)
                           ;
   U3726 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_14_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(14), ZN => n9363
                           );
   U3728 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_13_port, A2 => 
                           n9893, B1 => n9377, B2 => DRAM_DATA(13), ZN => n9364
                           );
   U3730 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_12_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(12), ZN => n9365
                           );
   U3732 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_11_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(11), ZN => n9366
                           );
   U3734 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_10_port, A2 => 
                           n9893, B1 => n9377, B2 => DRAM_DATA(10), ZN => n9367
                           );
   U3736 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_9_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(9), ZN => n9368)
                           ;
   U3738 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_8_port, A2 => 
                           n9893, B1 => n9377, B2 => DRAM_DATA(8), ZN => n9369)
                           ;
   U3740 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_7_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(7), ZN => n9370)
                           ;
   U3742 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_6_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(6), ZN => n9371)
                           ;
   U3744 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_5_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(5), ZN => n9372)
                           ;
   U3746 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_4_port, A2 => 
                           n9893, B1 => n9377, B2 => DRAM_DATA(4), ZN => n9373)
                           ;
   U3748 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_3_port, A2 => 
                           n9893, B1 => n9377, B2 => DRAM_DATA(3), ZN => n9374)
                           ;
   U3750 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_2_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(2), ZN => n9375)
                           ;
   U3752 : AOI22_X1 port map( A1 => n9377, A2 => DRAM_DATA(1), B1 => n9893, B2 
                           => datapath_i_alu_output_val_i_1_port, ZN => n9376);
   U3754 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_0_port, A2 => 
                           n9378, B1 => n9377, B2 => DRAM_DATA(0), ZN => n9379)
                           ;
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => n4417);
   clk_r_REG14604_S7 : DFFR_X1 port map( D => n1445, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_12_port, QN => n_4318);
   clk_r_REG16751_S2 : DFFS_X1 port map( D => n6808, CK => CLK, SN => RST, Q =>
                           n9122, QN => n_4319);
   clk_r_REG13715_S2 : DFF_X1 port map( D => n1673, CK => CLK, Q => n8930, QN 
                           => n_4320);
   clk_r_REG16835_S6 : DFFR_X1 port map( D => n5388, CK => CLK, RN => RST, Q =>
                           n9054, QN => n9887);
   clk_r_REG16691_S2 : DFFR_X1 port map( D => n9532, CK => CLK, RN => RST, Q =>
                           n_4321, QN => n9141);
   clk_r_REG16756_S4 : DFFR_X1 port map( D => n9173, CK => CLK, RN => RST, Q =>
                           n_4322, QN => n8945);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => n8718, Q => 
                           n5388);
   clk_r_REG16932_S7 : DFFR_X1 port map( D => n6887, CK => CLK, RN => RST, Q =>
                           n8716, QN => n_4323);
   clk_r_REG16609_S4 : DFFS_X1 port map( D => n9610, CK => CLK, SN => RST, Q =>
                           n9052, QN => n_4324);
   clk_r_REG16608_S4 : DFFS_X1 port map( D => n9610, CK => CLK, SN => RST, Q =>
                           n_4325, QN => n9073);
   clk_r_REG16592_S4 : DFFS_X1 port map( D => n9194, CK => CLK, SN => RST, Q =>
                           n9053, QN => n_4326);
   clk_r_REG16750_S2 : DFFS_X1 port map( D => n6808, CK => CLK, SN => RST, Q =>
                           n8626, QN => n_4327);
   clk_r_REG16745_S2 : DFFS_X1 port map( D => n9531, CK => CLK, SN => RST, Q =>
                           n9013, QN => n_4328);
   clk_r_REG16833_S6 : DFFS_X1 port map( D => n9535, CK => CLK, SN => RST, Q =>
                           n9883, QN => n8773);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X2 port map( A => 
                           n8847, EN => n9891, Z => DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X2 port map( A => 
                           n8844, EN => n9141, Z => DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X2 port map( A => 
                           n8784, EN => n8999, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X2 port map( A => 
                           n8835, EN => n9891, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X2 port map( A => 
                           n8829, EN => n9891, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X2 port map( A => 
                           n8841, EN => n9141, Z => DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X2 port map( A => 
                           n8838, EN => n9141, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X2 port map( A => 
                           n8826, EN => n9141, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X2 port map( A => 
                           n8832, EN => n8999, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X2 port map( A => 
                           n8874, EN => n9891, Z => DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X2 port map( A => 
                           n8868, EN => n9891, Z => DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X2 port map( A => 
                           n8865, EN => n9891, Z => DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X2 port map( A => 
                           n8859, EN => n9891, Z => DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X2 port map( A => 
                           n8850, EN => n9891, Z => DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X2 port map( A => 
                           n8814, EN => n9891, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X2 port map( A => 
                           n8808, EN => n9891, Z => DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X2 port map( A => 
                           n8802, EN => n9891, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X2 port map( A => 
                           n8796, EN => n9891, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X2 port map( A => 
                           n8781, EN => n9891, Z => DRAM_DATA(0));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X2 port map( A => 
                           n8871, EN => n9141, Z => DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X2 port map( A => 
                           n8862, EN => n9141, Z => DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X2 port map( A => 
                           n8853, EN => n9141, Z => DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X2 port map( A => 
                           n8820, EN => n9141, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X2 port map( A => 
                           n8805, EN => n9141, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X2 port map( A => 
                           n8793, EN => n9141, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X2 port map( A => 
                           n8856, EN => n8999, Z => DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X2 port map( A => 
                           n8823, EN => n8999, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X2 port map( A => 
                           n8817, EN => n8999, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X2 port map( A => 
                           n8811, EN => n8999, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X2 port map( A => 
                           n8799, EN => n8999, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X2 port map( A => 
                           n8790, EN => n8999, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X2 port map( A => 
                           n8787, EN => n8999, Z => DRAM_DATA(2));
   U3981 : OAI21_X2 port map( B1 => n8742, B2 => n8982, A => n9725, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U3982 : INV_X1 port map( A => n4337, ZN => n9609);
   U3983 : INV_X1 port map( A => n9609, ZN => n9610);
   U3984 : AOI22_X2 port map( A1 => n5388, A2 => n9542, B1 => n9074, B2 => 
                           n9535, ZN => n9531);
   U3985 : BUF_X1 port map( A => n9209, Z => IRAM_ADDRESS_31_port);
   U3986 : AOI22_X1 port map( A1 => n9054, A2 => cu_i_cmd_alu_op_type_2_port, 
                           B1 => n9121, B2 => n8776, ZN => n9675);
   U3987 : NOR2_X1 port map( A1 => n9675, A2 => n9671, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U3988 : NOR2_X1 port map( A1 => n9674, A2 => n9670, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U3989 : NOR2_X1 port map( A1 => n9677, A2 => n9676, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U3990 : CLKBUF_X1 port map( A => n8945, Z => n9841);
   U3991 : MUX2_X1 port map( A => IRAM_DATA(22), B => n8705, S => n9054, Z => 
                           n6902);
   U3992 : INV_X1 port map( A => n5388, ZN => n9535);
   U3993 : AOI22_X1 port map( A1 => n8773, A2 => n8998, B1 => n8931, B2 => 
                           IRAM_DATA(1), ZN => n9807);
   U3994 : INV_X1 port map( A => n9807, ZN => n9603);
   U3995 : AOI22_X1 port map( A1 => n8773, A2 => n8997, B1 => n8931, B2 => 
                           IRAM_DATA(2), ZN => n9808);
   U3996 : INV_X1 port map( A => n9808, ZN => n9604);
   U3997 : AOI22_X1 port map( A1 => n8773, A2 => n9119, B1 => n8931, B2 => 
                           IRAM_DATA(29), ZN => n9840);
   U3998 : INV_X1 port map( A => n9840, ZN => n9540);
   U3999 : AOI22_X1 port map( A1 => n8773, A2 => n9118, B1 => n8931, B2 => 
                           IRAM_DATA(30), ZN => n9615);
   U4000 : INV_X1 port map( A => n9615, ZN => n9545);
   U4001 : AOI22_X1 port map( A1 => n8773, A2 => n9110, B1 => n8931, B2 => 
                           IRAM_DATA(31), ZN => n9627);
   U4002 : NAND3_X1 port map( A1 => n9540, A2 => n9545, A3 => n9627, ZN => 
                           n9626);
   U4003 : INV_X1 port map( A => n9626, ZN => n9539);
   U4004 : NOR2_X1 port map( A1 => n8771, A2 => n9048, ZN => n9722);
   U4005 : NAND2_X1 port map( A1 => n9722, A2 => n9026, ZN => n9717);
   U4006 : OAI211_X1 port map( C1 => n9722, C2 => n9026, A => n9072, B => n9717
                           , ZN => n9612);
   U4007 : NAND2_X1 port map( A1 => n8618, A2 => n9612, ZN => n9766);
   U4008 : INV_X1 port map( A => n9766, ZN => n9571);
   U4009 : NOR2_X1 port map( A1 => n9046, A2 => n9717, ZN => n9716);
   U4010 : NAND2_X1 port map( A1 => n9716, A2 => n9027, ZN => n9711);
   U4011 : OAI211_X1 port map( C1 => n9716, C2 => n9027, A => n9072, B => n9711
                           , ZN => n9613);
   U4012 : NAND2_X1 port map( A1 => n8617, A2 => n9613, ZN => n9727);
   U4013 : INV_X1 port map( A => n9727, ZN => n9570);
   U4014 : AOI22_X1 port map( A1 => n8773, A2 => n9104, B1 => n8931, B2 => 
                           IRAM_DATA(27), ZN => n9616);
   U4015 : INV_X1 port map( A => n9616, ZN => n9550);
   U4016 : INV_X1 port map( A => n9627, ZN => n9547);
   U4017 : AOI22_X1 port map( A1 => n8773, A2 => n8995, B1 => n8931, B2 => 
                           IRAM_DATA(26), ZN => n9869);
   U4018 : AOI22_X1 port map( A1 => n8773, A2 => n8996, B1 => n8931, B2 => 
                           IRAM_DATA(28), ZN => n9631);
   U4019 : NAND2_X1 port map( A1 => n9631, A2 => n9550, ZN => n9810);
   U4020 : NOR3_X1 port map( A1 => n9869, A2 => n9545, A3 => n9810, ZN => n9614
                           );
   U4021 : NAND2_X1 port map( A1 => n9614, A2 => n9547, ZN => n9636);
   U4022 : NOR2_X1 port map( A1 => n9888, A2 => n9636, ZN => n9546);
   U4023 : INV_X1 port map( A => n9546, ZN => n9839);
   U4024 : NOR2_X1 port map( A1 => n9540, A2 => n9839, ZN => 
                           cu_i_cmd_word_3_port);
   U4025 : OAI22_X1 port map( A1 => n9535, A2 => cu_i_cmd_word_3_port, B1 => 
                           n8703, B2 => n5388, ZN => n9633);
   U4026 : INV_X1 port map( A => n9633, ZN => n9534);
   U4027 : NAND2_X1 port map( A1 => n9616, A2 => n9869, ZN => n7739);
   U4028 : INV_X1 port map( A => n9631, ZN => n9605);
   U4029 : INV_X1 port map( A => n7739, ZN => n9622);
   U4030 : NAND2_X1 port map( A1 => n9622, A2 => n9605, ZN => n9637);
   U4031 : NAND2_X1 port map( A1 => n9627, A2 => n9615, ZN => n9630);
   U4032 : NOR2_X1 port map( A1 => n9540, A2 => n9630, ZN => n9621);
   U4033 : NAND2_X1 port map( A1 => n9621, A2 => n9882, ZN => n9620);
   U4034 : AOI21_X1 port map( B1 => n9810, B2 => n9637, A => n9620, ZN => 
                           cu_i_cmd_word_6_port);
   U4035 : INV_X1 port map( A => n9869, ZN => n9606);
   U4036 : NAND2_X1 port map( A1 => n9616, A2 => n9606, ZN => n474);
   U4037 : NOR3_X1 port map( A1 => n9631, A2 => n9620, A3 => n474, ZN => n8055)
                           ;
   U4038 : AOI22_X1 port map( A1 => n5388, A2 => cu_i_cmd_word_6_port, B1 => 
                           n8709, B2 => n9535, ZN => n9619);
   U4039 : AOI22_X1 port map( A1 => n5388, A2 => n8055, B1 => n9001, B2 => 
                           n9535, ZN => n9617);
   U4040 : NAND2_X1 port map( A1 => n8730, A2 => n9617, ZN => n9618);
   U4041 : OAI22_X1 port map( A1 => n9619, A2 => n9618, B1 => n8730, B2 => 
                           n9617, ZN => n9530);
   U4042 : NOR2_X1 port map( A1 => n9810, A2 => n9620, ZN => n9541);
   U4043 : NAND3_X1 port map( A1 => n9622, A2 => n9631, A3 => n9621, ZN => 
                           n9544);
   U4044 : INV_X1 port map( A => n9544, ZN => n9693);
   U4045 : NAND2_X1 port map( A1 => n9693, A2 => n9882, ZN => n9543);
   U4046 : NOR2_X1 port map( A1 => n8773, A2 => IRAM_DATA(4), ZN => n9623);
   U4047 : AOI21_X1 port map( B1 => n9203, B2 => n8773, A => n9623, ZN => n6900
                           );
   U4048 : MUX2_X1 port map( A => IRAM_DATA(3), B => n8723, S => n8773, Z => 
                           n6898);
   U4049 : AOI22_X1 port map( A1 => n8773, A2 => n9105, B1 => n8931, B2 => 
                           IRAM_DATA(5), ZN => n9624);
   U4050 : INV_X1 port map( A => n9624, ZN => n9549);
   U4051 : NAND2_X1 port map( A1 => n8931, A2 => IRAM_DATA(0), ZN => n9625);
   U4052 : OAI21_X1 port map( B1 => n9883, B2 => n9174, A => n9625, ZN => n9548
                           );
   U4053 : AOI211_X1 port map( C1 => n9631, C2 => n9869, A => n9550, B => n9626
                           , ZN => n4060);
   U4054 : NAND2_X1 port map( A1 => n9627, A2 => n9545, ZN => n9628);
   U4055 : NOR4_X1 port map( A1 => n9631, A2 => n9606, A3 => n9540, A4 => n9628
                           , ZN => n6896);
   U4056 : INV_X1 port map( A => n9541, ZN => n9872);
   U4057 : NAND4_X1 port map( A1 => n6900, A2 => n6898, A3 => n9549, A4 => 
                           n9548, ZN => n9629);
   U4058 : NOR3_X1 port map( A1 => n9807, A2 => n9808, A3 => n9629, ZN => n9656
                           );
   U4059 : NOR2_X1 port map( A1 => n9840, A2 => n9630, ZN => n9868);
   U4060 : OAI21_X1 port map( B1 => n9631, B2 => n9550, A => n9606, ZN => n9632
                           );
   U4061 : AOI211_X1 port map( C1 => n9868, C2 => n9632, A => n4060, B => n6896
                           , ZN => n9695);
   U4062 : OAI222_X1 port map( A1 => n9872, A2 => n9869, B1 => n9543, B2 => 
                           n9656, C1 => n9695, C2 => n8745, ZN => n302);
   U4063 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n302, ZN => n6933
                           );
   U4064 : OAI22_X1 port map( A1 => n9535, A2 => n9546, B1 => n8702, B2 => 
                           n5388, ZN => n7193);
   U4065 : INV_X1 port map( A => n7193, ZN => n9533);
   U4066 : NAND2_X1 port map( A1 => n9533, A2 => n9633, ZN => n7215);
   U4067 : INV_X1 port map( A => n7215, ZN => n9532);
   U4068 : AOI22_X1 port map( A1 => n9054, A2 => n9099, B1 => n9121, B2 => 
                           IRAM_DATA(13), ZN => n9873);
   U4069 : INV_X1 port map( A => n9873, ZN => n9538);
   U4070 : AOI22_X1 port map( A1 => n9054, A2 => n9098, B1 => n9121, B2 => 
                           IRAM_DATA(18), ZN => n9875);
   U4071 : INV_X1 port map( A => n9875, ZN => n9537);
   U4072 : AOI22_X1 port map( A1 => n9054, A2 => n8719, B1 => IRAM_DATA(19), B2
                           => n9887, ZN => n9583);
   U4073 : INV_X1 port map( A => n9583, ZN => curr_instruction_to_cu_i_19_port)
                           ;
   U4074 : MUX2_X1 port map( A => IRAM_DATA(20), B => n8717, S => n9054, Z => 
                           curr_instruction_to_cu_i_20_port);
   U4075 : NOR2_X1 port map( A1 => n9044, A2 => n9711, ZN => n9710);
   U4076 : NAND2_X1 port map( A1 => n9710, A2 => n9028, ZN => n9714);
   U4077 : OAI211_X1 port map( C1 => n9710, C2 => n9028, A => n9072, B => n9714
                           , ZN => n9634);
   U4078 : NAND2_X1 port map( A1 => n8616, A2 => n9634, ZN => n9775);
   U4079 : INV_X1 port map( A => n9775, ZN => n9568);
   U4080 : INV_X1 port map( A => cu_i_n151, ZN => n9528);
   U4081 : NOR2_X1 port map( A1 => n4417, A2 => n3284, ZN => n9635);
   U4082 : NOR2_X1 port map( A1 => n9635, A2 => n9528, ZN => n9527);
   U4083 : NAND3_X1 port map( A1 => cu_i_n151, A2 => n9635, A3 => n6942, ZN => 
                           n6894);
   U4084 : MUX2_X1 port map( A => IRAM_DATA(14), B => n8720, S => n9054, Z => 
                           n6890);
   U4085 : INV_X1 port map( A => n9872, ZN => n9892);
   U4086 : INV_X1 port map( A => n9527, ZN => n9645);
   U4087 : NAND2_X1 port map( A1 => n9645, A2 => n6894, ZN => n9657);
   U4088 : AOI21_X1 port map( B1 => n9656, B2 => n9657, A => n9543, ZN => n9876
                           );
   U4089 : INV_X1 port map( A => n9876, ZN => n9874);
   U4090 : AOI221_X1 port map( B1 => n9874, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n9876, C2 =>
                           n6890, A => n9892, ZN => n9878);
   U4091 : INV_X1 port map( A => n9878, ZN => n9522);
   U4092 : OAI211_X1 port map( C1 => n9637, C2 => n9547, A => n9695, B => n9636
                           , ZN => n9692);
   U4093 : AOI21_X1 port map( B1 => n9882, B2 => n9692, A => n8055, ZN => n9641
                           );
   U4094 : NAND2_X1 port map( A1 => n9641, A2 => n9872, ZN => n7737);
   U4095 : CLKBUF_X1 port map( A => n7737, Z => n9895);
   U4096 : NOR2_X1 port map( A1 => n9042, A2 => n9714, ZN => n9713);
   U4097 : NAND2_X1 port map( A1 => n9713, A2 => n9029, ZN => n9720);
   U4098 : OAI211_X1 port map( C1 => n9713, C2 => n9029, A => n9072, B => n9720
                           , ZN => n9638);
   U4099 : NAND2_X1 port map( A1 => n8615, A2 => n9638, ZN => n9854);
   U4100 : INV_X1 port map( A => n9854, ZN => n9567);
   U4101 : MUX2_X1 port map( A => IRAM_DATA(15), B => n8716, S => n9054, Z => 
                           n6887);
   U4102 : AOI221_X1 port map( B1 => n9874, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n9876, C2 =>
                           n6887, A => n9892, ZN => n9639);
   U4103 : INV_X1 port map( A => n9639, ZN => n9525);
   U4104 : MUX2_X1 port map( A => IRAM_DATA(16), B => n8715, S => n9054, Z => 
                           curr_instruction_to_cu_i_16_port);
   U4105 : MUX2_X1 port map( A => IRAM_DATA(11), B => n8722, S => n8773, Z => 
                           n6889);
   U4106 : AOI221_X1 port map( B1 => n9874, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n9876, C2 =>
                           n6889, A => n9892, ZN => n9640);
   U4107 : INV_X1 port map( A => n9640, ZN => n9524);
   U4108 : MUX2_X1 port map( A => IRAM_DATA(12), B => n8721, S => n9054, Z => 
                           n6892);
   U4109 : MUX2_X1 port map( A => IRAM_DATA(17), B => n8714, S => n9054, Z => 
                           curr_instruction_to_cu_i_17_port);
   U4110 : NAND2_X1 port map( A1 => n9641, A2 => n9874, ZN => enable_rf_i);
   U4111 : INV_X1 port map( A => n9543, ZN => n9642);
   U4112 : NAND2_X1 port map( A1 => n9642, A2 => n9656, ZN => n6928);
   U4113 : OAI21_X1 port map( B1 => n9645, B2 => n6928, A => n8658, ZN => 
                           write_rf_i);
   U4114 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U4115 : AOI22_X1 port map( A1 => n8989, A2 => n8983, B1 => n8948, B2 => 
                           n8744, ZN => n9643);
   U4116 : INV_X1 port map( A => n9643, ZN => n9644);
   U4117 : AOI21_X1 port map( B1 => n8991, B2 => 
                           datapath_i_alu_output_val_i_9_port, A => n9644, ZN 
                           => n9782);
   U4118 : INV_X1 port map( A => n9782, ZN => n9607);
   U4119 : NOR2_X1 port map( A1 => n9645, A2 => n6928, ZN => n9646);
   U4120 : NOR2_X1 port map( A1 => n9646, A2 => n8660, ZN => n9650);
   U4121 : AND3_X1 port map( A1 => n9650, A2 => n9841, A3 => DRAM_READY, ZN => 
                           n9377);
   U4122 : CLKBUF_X1 port map( A => n9377, Z => n9894);
   U4123 : NOR2_X1 port map( A1 => n9040, A2 => n9720, ZN => n9719);
   U4124 : NAND2_X1 port map( A1 => n9719, A2 => n9030, ZN => n9702);
   U4125 : OAI211_X1 port map( C1 => n9719, C2 => n9030, A => n9072, B => n9702
                           , ZN => n9647);
   U4126 : NAND2_X1 port map( A1 => n8614, A2 => n9647, ZN => n9759);
   U4127 : INV_X1 port map( A => n9759, ZN => n9566);
   U4128 : AOI22_X1 port map( A1 => n8989, A2 => n9056, B1 => n8948, B2 => 
                           n8746, ZN => n9648);
   U4129 : INV_X1 port map( A => n9648, ZN => n9649);
   U4130 : AOI21_X1 port map( B1 => n8991, B2 => 
                           datapath_i_alu_output_val_i_7_port, A => n9649, ZN 
                           => n9780);
   U4131 : INV_X1 port map( A => n9780, ZN => n9582);
   U4132 : NOR2_X1 port map( A1 => n9650, A2 => n8947, ZN => n9378);
   U4133 : CLKBUF_X1 port map( A => n9378, Z => n9893);
   U4134 : NOR2_X1 port map( A1 => n9038, A2 => n9702, ZN => n9701);
   U4135 : NAND2_X1 port map( A1 => n9701, A2 => n9031, ZN => n9708);
   U4136 : OAI211_X1 port map( C1 => n9701, C2 => n9031, A => n9072, B => n9708
                           , ZN => n9651);
   U4137 : NAND2_X1 port map( A1 => n8613, A2 => n9651, ZN => n9756);
   U4138 : INV_X1 port map( A => n9756, ZN => n9565);
   U4139 : AOI21_X1 port map( B1 => n8991, B2 => 
                           datapath_i_alu_output_val_i_5_port, A => n9078, ZN 
                           => n9781);
   U4140 : INV_X1 port map( A => n9781, ZN => n9552);
   U4141 : NOR2_X1 port map( A1 => n9036, A2 => n9708, ZN => n9707);
   U4142 : NAND2_X1 port map( A1 => n9707, A2 => n9032, ZN => n9705);
   U4143 : OAI211_X1 port map( C1 => n9707, C2 => n9032, A => n9072, B => n9705
                           , ZN => n9652);
   U4144 : NAND2_X1 port map( A1 => n8612, A2 => n9652, ZN => n9754);
   U4145 : INV_X1 port map( A => n9754, ZN => n9564);
   U4146 : NOR2_X1 port map( A1 => n9034, A2 => n9705, ZN => n9704);
   U4147 : NAND2_X1 port map( A1 => n9704, A2 => n9033, ZN => n9654);
   U4148 : XOR2_X1 port map( A => n9209, B => n9654, Z => n9653);
   U4149 : AOI22_X1 port map( A1 => n9072, A2 => n9653, B1 => n9051, B2 => 
                           n8731, ZN => n9860);
   U4150 : INV_X1 port map( A => n9860, ZN => n9562);
   U4151 : OAI211_X1 port map( C1 => n9704, C2 => n9033, A => n9072, B => n9654
                           , ZN => n9655);
   U4152 : NAND2_X1 port map( A1 => n8611, A2 => n9655, ZN => n9752);
   U4153 : INV_X1 port map( A => n9752, ZN => n9563);
   U4154 : NAND2_X1 port map( A1 => n9693, A2 => n9656, ZN => n477);
   U4155 : INV_X1 port map( A => n9657, ZN => n9658);
   U4156 : OAI21_X1 port map( B1 => n9658, B2 => n9543, A => n8737, ZN => n9659
                           );
   U4157 : OAI221_X1 port map( B1 => n9659, B2 => n9011, C1 => n9659, C2 => 
                           n477, A => n9535, ZN => n9526);
   U4158 : INV_X1 port map( A => datapath_i_alu_output_val_i_2_port, ZN => 
                           n9660);
   U4159 : OAI22_X1 port map( A1 => n9053, A2 => n8932, B1 => n9660, B2 => 
                           n9884, ZN => n9661);
   U4160 : AOI21_X1 port map( B1 => n8948, B2 => n8609, A => n9661, ZN => n9584
                           );
   U4161 : INV_X1 port map( A => n9584, ZN => n9862);
   U4162 : AOI22_X1 port map( A1 => n8610, A2 => n9052, B1 => n9073, B2 => 
                           n9862, ZN => n9864);
   U4163 : INV_X1 port map( A => n9864, ZN => n9560);
   U4164 : AOI22_X1 port map( A1 => n8948, A2 => n8729, B1 => n8951, B2 => 
                           datapath_i_alu_output_val_i_3_port, ZN => n9662);
   U4165 : OAI21_X1 port map( B1 => n9053, B2 => n8935, A => n9662, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U4166 : NAND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_3_port,
                           A2 => n9862, ZN => n9779);
   U4167 : OAI211_X1 port map( C1 => n9862, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n9073, B => n9779, ZN => n9663);
   U4168 : NAND2_X1 port map( A1 => n8625, A2 => n9663, ZN => n9866);
   U4169 : INV_X1 port map( A => n9866, ZN => n9559);
   U4170 : AOI22_X1 port map( A1 => n8991, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n8948, B2 
                           => n8738, ZN => n9664);
   U4171 : OAI21_X1 port map( B1 => n9053, B2 => n8938, A => n9664, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U4172 : INV_X1 port map( A => n9779, ZN => n9665);
   U4173 : NAND2_X1 port map( A1 => n9665, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n9679);
   U4174 : OAI211_X1 port map( C1 => n9665, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n9073, B => n9679, ZN => n9666);
   U4175 : NAND2_X1 port map( A1 => n8624, A2 => n9666, ZN => n9777);
   U4176 : INV_X1 port map( A => n9777, ZN => n9561);
   U4177 : INV_X1 port map( A => n9152, ZN => IRAM_ADDRESS_1_port);
   U4178 : AOI22_X1 port map( A1 => n8948, A2 => n9079, B1 => n8951, B2 => 
                           datapath_i_alu_output_val_i_1_port, ZN => n9667);
   U4179 : OAI21_X1 port map( B1 => n9053, B2 => n9015, A => n9667, ZN => n5478
                           );
   U4180 : AOI22_X1 port map( A1 => n9052, A2 => IRAM_ADDRESS_1_port, B1 => 
                           n9073, B2 => n5478, ZN => n7839);
   U4181 : AOI22_X1 port map( A1 => n8991, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n8948, B2 
                           => n8739, ZN => n9668);
   U4182 : OAI21_X1 port map( B1 => n9053, B2 => n8941, A => n9668, ZN => n1453
                           );
   U4183 : NOR2_X1 port map( A1 => n9781, A2 => n9679, ZN => n9678);
   U4184 : NAND2_X1 port map( A1 => n9678, A2 => n1453, ZN => n9686);
   U4185 : OAI211_X1 port map( C1 => n9678, C2 => n1453, A => n9073, B => n9686
                           , ZN => n9669);
   U4186 : NAND2_X1 port map( A1 => n8623, A2 => n9669, ZN => n9761);
   U4187 : INV_X1 port map( A => n9761, ZN => n9558);
   U4188 : AOI22_X1 port map( A1 => n9054, A2 => cu_i_cmd_alu_op_type_0_port, 
                           B1 => n9121, B2 => n8778, ZN => n9674);
   U4189 : AOI22_X1 port map( A1 => n9054, A2 => cu_i_cmd_alu_op_type_1_port, 
                           B1 => n9121, B2 => n8777, ZN => n9677);
   U4190 : AOI22_X1 port map( A1 => n9054, A2 => cu_i_cmd_alu_op_type_3_port, 
                           B1 => n9121, B2 => n8775, ZN => n9673);
   U4191 : AOI21_X1 port map( B1 => n9675, B2 => n9677, A => n9673, ZN => n9670
                           );
   U4192 : INV_X1 port map( A => n9673, ZN => n9671);
   U4193 : OAI211_X1 port map( C1 => n9674, C2 => n9677, A => n9671, B => n9675
                           , ZN => n9672);
   U4194 : INV_X1 port map( A => n9672, ZN => n9529);
   U4195 : AOI21_X1 port map( B1 => n9675, B2 => n9674, A => n9673, ZN => n9676
                           );
   U4196 : AOI211_X1 port map( C1 => n9781, C2 => n9679, A => n9052, B => n9678
                           , ZN => n9680);
   U4197 : NOR2_X1 port map( A1 => n8638, A2 => n9680, ZN => n9553);
   U4198 : INV_X1 port map( A => n9553, ZN => n9773);
   U4199 : AOI22_X1 port map( A1 => n9010, A2 => n8988, B1 => n9008, B2 => 
                           n9773, ZN => n9681);
   U4200 : INV_X1 port map( A => n9681, ZN => n9554);
   U4201 : INV_X1 port map( A => datapath_i_alu_output_val_i_8_port, ZN => 
                           n9682);
   U4202 : OAI222_X1 port map( A1 => n9682, A2 => n8993, B1 => n9053, B2 => 
                           n9075, C1 => n9077, C2 => n8950, ZN => n1449);
   U4203 : NOR2_X1 port map( A1 => n9780, A2 => n9686, ZN => n9685);
   U4204 : NAND2_X1 port map( A1 => n9685, A2 => n1449, ZN => n9688);
   U4205 : OAI211_X1 port map( C1 => n9685, C2 => n1449, A => n9073, B => n9688
                           , ZN => n9683);
   U4206 : NAND2_X1 port map( A1 => n8622, A2 => n9683, ZN => n9769);
   U4207 : INV_X1 port map( A => n9769, ZN => n9555);
   U4208 : INV_X1 port map( A => n9153, ZN => IRAM_ADDRESS_0_port);
   U4209 : AOI22_X1 port map( A1 => n8991, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n8948, B2 
                           => n9070, ZN => n9684);
   U4210 : OAI21_X1 port map( B1 => n9053, B2 => n9018, A => n9684, ZN => n5479
                           );
   U4211 : AOI22_X1 port map( A1 => n9052, A2 => IRAM_ADDRESS_0_port, B1 => 
                           n9073, B2 => n5479, ZN => n7852);
   U4212 : AOI211_X1 port map( C1 => n9780, C2 => n9686, A => n9052, B => n9685
                           , ZN => n9687);
   U4213 : NOR2_X1 port map( A1 => n8639, A2 => n9687, ZN => n9557);
   U4214 : OR2_X1 port map( A1 => n8055, A2 => cu_i_cmd_word_6_port, ZN => 
                           n9542);
   U4215 : AOI221_X1 port map( B1 => n9012, B2 => n9535, C1 => n9542, C2 => 
                           n5388, A => n9021, ZN => n4337);
   U4216 : NOR2_X1 port map( A1 => n9782, A2 => n9688, ZN => n9880);
   U4217 : AOI211_X1 port map( C1 => n9782, C2 => n9688, A => n9052, B => n9880
                           , ZN => n9689);
   U4218 : NOR2_X1 port map( A1 => n8637, A2 => n9689, ZN => n9556);
   U4219 : OAI211_X1 port map( C1 => n9025, C2 => n8740, A => n9072, B => n8771
                           , ZN => n9690);
   U4220 : NAND2_X1 port map( A1 => n8619, A2 => n9690, ZN => n9747);
   U4221 : INV_X1 port map( A => n9747, ZN => n9569);
   U4222 : INV_X1 port map( A => n9530, ZN => n9700);
   U4223 : AND2_X1 port map( A1 => n8994, A2 => n9700, ZN => n9170);
   U4224 : OR3_X1 port map( A1 => n9537, A2 => curr_instruction_to_cu_i_19_port
                           , A3 => curr_instruction_to_cu_i_20_port, ZN => 
                           n9691);
   U4225 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_16_port, A2 => 
                           curr_instruction_to_cu_i_17_port, A3 => n9691, ZN =>
                           n9694);
   U4226 : OAI22_X1 port map( A1 => n9695, A2 => n9694, B1 => n9693, B2 => 
                           n9692, ZN => n9699);
   U4227 : INV_X1 port map( A => n6892, ZN => n9870);
   U4228 : NOR4_X1 port map( A1 => n6889, A2 => n6890, A3 => n6887, A4 => n9538
                           , ZN => n9697);
   U4229 : AOI211_X1 port map( C1 => n8727, C2 => n8641, A => n9546, B => n9542
                           , ZN => n9696);
   U4230 : OAI221_X1 port map( B1 => n9543, B2 => n9870, C1 => n9543, C2 => 
                           n9697, A => n9696, ZN => n9698);
   U4231 : AOI21_X1 port map( B1 => n9882, B2 => n9699, A => n9698, ZN => n4052
                           );
   U4232 : OR2_X1 port map( A1 => n4052, A2 => n9003, ZN => n9180);
   U4233 : AND2_X1 port map( A1 => n8769, A2 => n9700, ZN => n9169);
   U4234 : CLKBUF_X1 port map( A => n9141, Z => n9891);
   U4235 : AOI211_X1 port map( C1 => n9039, C2 => n9702, A => n9051, B => n9701
                           , ZN => n9703);
   U4236 : OR2_X1 port map( A1 => n8629, A2 => n9703, ZN => n9589);
   U4237 : AOI211_X1 port map( C1 => n9035, C2 => n9705, A => n9051, B => n9704
                           , ZN => n9706);
   U4238 : OR2_X1 port map( A1 => n8627, A2 => n9706, ZN => n9597);
   U4239 : AOI211_X1 port map( C1 => n9037, C2 => n9708, A => n9051, B => n9707
                           , ZN => n9709);
   U4240 : OR2_X1 port map( A1 => n8628, A2 => n9709, ZN => n9595);
   U4241 : AOI211_X1 port map( C1 => n9045, C2 => n9711, A => n9051, B => n9710
                           , ZN => n9712);
   U4242 : OR2_X1 port map( A1 => n8632, A2 => n9712, ZN => n9591);
   U4243 : AOI211_X1 port map( C1 => n9043, C2 => n9714, A => n9051, B => n9713
                           , ZN => n9715);
   U4244 : OR2_X1 port map( A1 => n8631, A2 => n9715, ZN => n9585);
   U4245 : AOI211_X1 port map( C1 => n9047, C2 => n9717, A => n9051, B => n9716
                           , ZN => n9718);
   U4246 : OR2_X1 port map( A1 => n8633, A2 => n9718, ZN => n9593);
   U4247 : AOI211_X1 port map( C1 => n9041, C2 => n9720, A => n9051, B => n9719
                           , ZN => n9721);
   U4248 : OR2_X1 port map( A1 => n8630, A2 => n9721, ZN => n9587);
   U4249 : AOI211_X1 port map( C1 => n8771, C2 => n9049, A => n9722, B => n9051
                           , ZN => n9723);
   U4250 : OR2_X1 port map( A1 => n8634, A2 => n9723, ZN => n9599);
   U4251 : AOI211_X1 port map( C1 => n9024, C2 => n8741, A => n8740, B => n9051
                           , ZN => n9724);
   U4252 : OR2_X1 port map( A1 => n8635, A2 => n9724, ZN => n9601);
   U4253 : OR2_X1 port map( A1 => n9095, A2 => n8767, ZN => cu_i_N278);
   U4254 : INV_X1 port map( A => n9145, ZN => IRAM_ADDRESS_14_port);
   U4255 : INV_X1 port map( A => n9142, ZN => IRAM_ADDRESS_16_port);
   U4256 : INV_X1 port map( A => n9148, ZN => IRAM_ADDRESS_18_port);
   U4257 : INV_X1 port map( A => n9150, ZN => IRAM_ADDRESS_20_port);
   U4258 : INV_X1 port map( A => n9147, ZN => IRAM_ADDRESS_22_port);
   U4259 : INV_X1 port map( A => n9143, ZN => IRAM_ADDRESS_24_port);
   U4260 : INV_X1 port map( A => n9146, ZN => IRAM_ADDRESS_26_port);
   U4261 : INV_X1 port map( A => n9149, ZN => IRAM_ADDRESS_28_port);
   U4262 : INV_X1 port map( A => n9144, ZN => IRAM_ADDRESS_30_port);
   U4263 : AOI22_X1 port map( A1 => n9171, A2 => n8743, B1 => n9013, B2 => 
                           n8889, ZN => n9725);
   U4264 : MUX2_X1 port map( A => n8664, B => n8791, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U4265 : MUX2_X1 port map( A => n8665, B => n8788, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U4266 : MUX2_X1 port map( A => n8666, B => n8785, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U4267 : INV_X1 port map( A => n9531, ZN => n9726);
   U4268 : NAND2_X1 port map( A1 => n9115, A2 => n9726, ZN => n6920);
   U4269 : NOR2_X1 port map( A1 => n9115, A2 => n9531, ZN => n6919);
   U4270 : AOI22_X1 port map( A1 => n8743, A2 => n9727, B1 => n9013, B2 => 
                           n8903, ZN => n9728);
   U4271 : OAI21_X1 port map( B1 => n8742, B2 => n9111, A => n9728, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U4272 : OAI21_X1 port map( B1 => n8742, B2 => n8985, A => n8640, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U4273 : MUX2_X1 port map( A => n8663, B => n8794, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U4274 : MUX2_X1 port map( A => IRAM_DATA(23), B => n8726, S => n9054, Z => 
                           n6881);
   U4275 : NAND2_X1 port map( A1 => n9074, A2 => n9535, ZN => n9729);
   U4276 : OAI21_X1 port map( B1 => n9120, B2 => n9535, A => n9729, ZN => n7789
                           );
   U4277 : NAND2_X1 port map( A1 => n9868, A2 => n9605, ZN => n2299);
   U4278 : AOI222_X1 port map( A1 => n9601, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_13_port, B2 => n8951, C1
                           => n8989, C2 => n8977, ZN => n9602);
   U4279 : AOI222_X1 port map( A1 => n9886, A2 => n9171, B1 => n8991, B2 => 
                           datapath_i_alu_output_val_i_11_port, C1 => n8989, C2
                           => n8980, ZN => n9608);
   U4280 : INV_X1 port map( A => datapath_i_alu_output_val_i_10_port, ZN => 
                           n9730);
   U4281 : OAI222_X1 port map( A1 => n9730, A2 => n8993, B1 => n9053, B2 => 
                           n8747, C1 => n8749, C2 => n8950, ZN => n1447);
   U4282 : INV_X1 port map( A => datapath_i_alu_output_val_i_12_port, ZN => 
                           n9731);
   U4283 : OAI222_X1 port map( A1 => n9731, A2 => n8993, B1 => n9053, B2 => 
                           n9068, C1 => n9179, C2 => n8950, ZN => n1445);
   U4284 : NAND2_X1 port map( A1 => n9880, A2 => n1447, ZN => n9879);
   U4285 : NOR2_X1 port map( A1 => n9608, A2 => n9879, ZN => n9742);
   U4286 : NAND2_X1 port map( A1 => n9742, A2 => n1445, ZN => n6917);
   U4287 : NOR2_X1 port map( A1 => n9602, A2 => n6917, ZN => n6916);
   U4288 : INV_X1 port map( A => datapath_i_alu_output_val_i_14_port, ZN => 
                           n9732);
   U4289 : OAI222_X1 port map( A1 => n9732, A2 => n9055, B1 => n9053, B2 => 
                           n9107, C1 => n9569, C2 => n8950, ZN => n1443);
   U4290 : NAND2_X1 port map( A1 => n6916, A2 => n1443, ZN => n7861);
   U4291 : INV_X1 port map( A => datapath_i_alu_output_val_i_16_port, ZN => 
                           n9733);
   U4292 : OAI222_X1 port map( A1 => n9733, A2 => n9055, B1 => n9053, B2 => 
                           n9113, C1 => n9571, C2 => n8950, ZN => n5342);
   U4293 : INV_X1 port map( A => datapath_i_alu_output_val_i_18_port, ZN => 
                           n9734);
   U4294 : OAI222_X1 port map( A1 => n9734, A2 => n9055, B1 => n9053, B2 => 
                           n9111, C1 => n9570, C2 => n8950, ZN => n5343);
   U4295 : INV_X1 port map( A => datapath_i_alu_output_val_i_20_port, ZN => 
                           n9735);
   U4296 : OAI222_X1 port map( A1 => n9735, A2 => n9055, B1 => n9053, B2 => 
                           n9102, C1 => n9568, C2 => n8950, ZN => n5344);
   U4297 : INV_X1 port map( A => datapath_i_alu_output_val_i_22_port, ZN => 
                           n9736);
   U4298 : OAI222_X1 port map( A1 => n9736, A2 => n9055, B1 => n9053, B2 => 
                           n9096, C1 => n9567, C2 => n8950, ZN => n5345);
   U4299 : INV_X1 port map( A => datapath_i_alu_output_val_i_24_port, ZN => 
                           n9737);
   U4300 : OAI222_X1 port map( A1 => n9737, A2 => n9055, B1 => n9053, B2 => 
                           n9093, C1 => n9566, C2 => n8950, ZN => n5346);
   U4301 : INV_X1 port map( A => datapath_i_alu_output_val_i_26_port, ZN => 
                           n9738);
   U4302 : OAI222_X1 port map( A1 => n9738, A2 => n9055, B1 => n9053, B2 => 
                           n9089, C1 => n9565, C2 => n8950, ZN => n5347);
   U4303 : INV_X1 port map( A => datapath_i_alu_output_val_i_28_port, ZN => 
                           n9739);
   U4304 : OAI222_X1 port map( A1 => n9739, A2 => n9055, B1 => n9053, B2 => 
                           n9085, C1 => n9564, C2 => n8950, ZN => n5348);
   U4305 : INV_X1 port map( A => datapath_i_alu_output_val_i_30_port, ZN => 
                           n9740);
   U4306 : OAI222_X1 port map( A1 => n9740, A2 => n9055, B1 => n9053, B2 => 
                           n9083, C1 => n9563, C2 => n8950, ZN => n5349);
   U4307 : OAI211_X1 port map( C1 => n9742, C2 => n1445, A => n9073, B => n6917
                           , ZN => n9741);
   U4308 : NAND2_X1 port map( A1 => n8620, A2 => n9741, ZN => n7912);
   U4309 : AOI211_X1 port map( C1 => n9608, C2 => n9879, A => n9052, B => n9742
                           , ZN => n9743);
   U4310 : NOR2_X1 port map( A1 => n8636, A2 => n9743, ZN => n4128);
   U4311 : MUX2_X1 port map( A => n8662, B => n8797, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U4312 : AOI22_X1 port map( A1 => n8891, A2 => n9013, B1 => n8743, B2 => 
                           n9885, ZN => n9744);
   U4313 : OAI21_X1 port map( B1 => n9068, B2 => n8742, A => n9744, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U4314 : AOI22_X1 port map( A1 => n8893, A2 => n9013, B1 => n8743, B2 => 
                           n9601, ZN => n9745);
   U4315 : OAI21_X1 port map( B1 => n8742, B2 => n8979, A => n9745, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U4316 : AOI22_X1 port map( A1 => n8743, A2 => n9002, B1 => n9013, B2 => 
                           n8887, ZN => n9746);
   U4317 : OAI21_X1 port map( B1 => n8747, B2 => n8742, A => n9746, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U4318 : MUX2_X1 port map( A => n8672, B => n8782, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U4319 : AOI22_X1 port map( A1 => n8895, A2 => n9013, B1 => n8743, B2 => 
                           n9747, ZN => n9748);
   U4320 : OAI21_X1 port map( B1 => n9107, B2 => n8742, A => n9748, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U4321 : AOI22_X1 port map( A1 => n8743, A2 => n9599, B1 => n9013, B2 => 
                           n8897, ZN => n9749);
   U4322 : OAI21_X1 port map( B1 => n8742, B2 => n8976, A => n9749, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U4323 : AOI22_X1 port map( A1 => n8743, A2 => n9591, B1 => n9013, B2 => 
                           n8905, ZN => n9750);
   U4324 : OAI21_X1 port map( B1 => n8742, B2 => n8970, A => n9750, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U4325 : AOI22_X1 port map( A1 => n8743, A2 => n9597, B1 => n9013, B2 => 
                           n8925, ZN => n9751);
   U4326 : OAI21_X1 port map( B1 => n8742, B2 => n8955, A => n9751, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U4327 : AOI22_X1 port map( A1 => n8743, A2 => n9752, B1 => n9013, B2 => 
                           n8927, ZN => n9753);
   U4328 : OAI21_X1 port map( B1 => n8742, B2 => n9083, A => n9753, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U4329 : AOI22_X1 port map( A1 => n8743, A2 => n9754, B1 => n9013, B2 => 
                           n8923, ZN => n9755);
   U4330 : OAI21_X1 port map( B1 => n8742, B2 => n9085, A => n9755, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U4331 : AOI22_X1 port map( A1 => n8743, A2 => n9756, B1 => n9013, B2 => 
                           n8919, ZN => n9757);
   U4332 : OAI21_X1 port map( B1 => n8742, B2 => n9089, A => n9757, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U4333 : AOI22_X1 port map( A1 => n8743, A2 => n9589, B1 => n9013, B2 => 
                           n8917, ZN => n9758);
   U4334 : OAI21_X1 port map( B1 => n8742, B2 => n8961, A => n9758, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U4335 : AOI22_X1 port map( A1 => n8743, A2 => n9759, B1 => n9013, B2 => 
                           n8915, ZN => n9760);
   U4336 : OAI21_X1 port map( B1 => n8742, B2 => n9093, A => n9760, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U4337 : AOI22_X1 port map( A1 => n9531, A2 => n8883, B1 => n6919, B2 => 
                           n9761, ZN => n9762);
   U4338 : OAI21_X1 port map( B1 => n8942, B2 => n6920, A => n9762, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);
   U4339 : INV_X1 port map( A => n9557, ZN => n9763);
   U4340 : AOI22_X1 port map( A1 => n9531, A2 => n8884, B1 => n6919, B2 => 
                           n9763, ZN => n9764);
   U4341 : OAI21_X1 port map( B1 => n9004, B2 => n6920, A => n9764, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U4342 : INV_X1 port map( A => n9556, ZN => n9765);
   U4343 : AOI22_X1 port map( A1 => n9531, A2 => n8886, B1 => n6919, B2 => 
                           n9765, ZN => n6823);
   U4344 : AOI22_X1 port map( A1 => n8743, A2 => n9766, B1 => n9013, B2 => 
                           n8899, ZN => n9767);
   U4345 : OAI21_X1 port map( B1 => n8742, B2 => n9113, A => n9767, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U4346 : NOR2_X1 port map( A1 => n9889, A2 => n9205, ZN => n9804);
   U4347 : INV_X1 port map( A => n9804, ZN => n9806);
   U4348 : NOR2_X1 port map( A1 => n9204, A2 => n9806, ZN => n9805);
   U4349 : NOR2_X1 port map( A1 => n9805, A2 => n9206, ZN => n9768);
   U4350 : AOI211_X1 port map( C1 => n9805, C2 => n9206, A => n8763, B => n9768
                           , ZN => cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U4352 : AOI22_X1 port map( A1 => n9531, A2 => n8885, B1 => n6919, B2 => 
                           n9769, ZN => n9770);
   U4353 : OAI21_X1 port map( B1 => n9076, B2 => n6920, A => n9770, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U4354 : INV_X1 port map( A => n7839, ZN => n9771);
   U4355 : AOI22_X1 port map( A1 => n9531, A2 => n8878, B1 => n6919, B2 => 
                           n9771, ZN => n9772);
   U4356 : OAI21_X1 port map( B1 => n9016, B2 => n6920, A => n9772, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U4357 : AOI22_X1 port map( A1 => n9531, A2 => n8882, B1 => n6919, B2 => 
                           n9773, ZN => n9774);
   U4358 : OAI21_X1 port map( B1 => n8986, B2 => n6920, A => n9774, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U4359 : AOI22_X1 port map( A1 => n8743, A2 => n9775, B1 => n9013, B2 => 
                           n8907, ZN => n9776);
   U4360 : OAI21_X1 port map( B1 => n8742, B2 => n9102, A => n9776, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U4361 : AOI22_X1 port map( A1 => n9531, A2 => n8881, B1 => n6919, B2 => 
                           n9777, ZN => n9778);
   U4362 : OAI21_X1 port map( B1 => n8939, B2 => n6920, A => n9778, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U4363 : NAND2_X1 port map( A1 => n8728, A2 => n4052, ZN => n6914);
   U4364 : NOR2_X1 port map( A1 => n9779, A2 => n9526, ZN => n9815);
   U4365 : NAND2_X1 port map( A1 => n9815, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n9814);
   U4366 : NOR2_X1 port map( A1 => n9781, A2 => n9814, ZN => n9817);
   U4367 : NAND2_X1 port map( A1 => n9817, A2 => n1453, ZN => n9816);
   U4368 : NOR2_X1 port map( A1 => n9780, A2 => n9816, ZN => n9819);
   U4369 : AOI211_X1 port map( C1 => n9780, C2 => n9816, A => n9819, B => n9609
                           , ZN => n6821);
   U4370 : AOI211_X1 port map( C1 => n9781, C2 => n9814, A => n9817, B => n9609
                           , ZN => n6820);
   U4371 : NAND2_X1 port map( A1 => n9819, A2 => n1449, ZN => n9818);
   U4372 : NOR2_X1 port map( A1 => n9782, A2 => n9818, ZN => n9821);
   U4373 : AOI211_X1 port map( C1 => n9782, C2 => n9818, A => n9821, B => n9609
                           , ZN => n6819);
   U4374 : NAND2_X1 port map( A1 => n9821, A2 => n1447, ZN => n9820);
   U4375 : NOR2_X1 port map( A1 => n9608, A2 => n9820, ZN => n9822);
   U4376 : AOI211_X1 port map( C1 => n9608, C2 => n9820, A => n9822, B => n9609
                           , ZN => n6818);
   U4377 : AOI211_X1 port map( C1 => n8736, C2 => n9023, A => n9073, B => n8735
                           , ZN => n6817);
   U4378 : NAND2_X1 port map( A1 => n9822, A2 => n1445, ZN => n6910);
   U4379 : NOR2_X1 port map( A1 => n9602, A2 => n6910, ZN => n8001);
   U4380 : NAND2_X1 port map( A1 => n8001, A2 => n1443, ZN => n8000);
   U4381 : NOR2_X1 port map( A1 => n9048, A2 => n8734, ZN => n9824);
   U4382 : AOI211_X1 port map( C1 => n8734, C2 => n9048, A => n9824, B => n9073
                           , ZN => n6816);
   U4383 : NAND2_X1 port map( A1 => n9026, A2 => n9824, ZN => n9823);
   U4384 : NOR2_X1 port map( A1 => n9046, A2 => n9823, ZN => n9826);
   U4385 : AOI211_X1 port map( C1 => n9046, C2 => n9823, A => n9826, B => n9073
                           , ZN => n6815);
   U4386 : NAND2_X1 port map( A1 => n9027, A2 => n9826, ZN => n9825);
   U4387 : NOR2_X1 port map( A1 => n9044, A2 => n9825, ZN => n9828);
   U4388 : AOI211_X1 port map( C1 => n9044, C2 => n9825, A => n9828, B => n9073
                           , ZN => n6814);
   U4389 : NAND2_X1 port map( A1 => n9028, A2 => n9828, ZN => n9827);
   U4390 : NOR2_X1 port map( A1 => n9042, A2 => n9827, ZN => n9830);
   U4391 : AOI211_X1 port map( C1 => n9042, C2 => n9827, A => n9830, B => n9073
                           , ZN => n6813);
   U4392 : NAND2_X1 port map( A1 => n9029, A2 => n9830, ZN => n9829);
   U4393 : NOR2_X1 port map( A1 => n9040, A2 => n9829, ZN => n9832);
   U4394 : AOI211_X1 port map( C1 => n9040, C2 => n9829, A => n9832, B => n9073
                           , ZN => n6812);
   U4395 : NAND2_X1 port map( A1 => n9030, A2 => n9832, ZN => n9831);
   U4396 : NOR2_X1 port map( A1 => n9038, A2 => n9831, ZN => n9834);
   U4397 : AOI211_X1 port map( C1 => n9038, C2 => n9831, A => n9834, B => n9073
                           , ZN => n6811);
   U4398 : NAND2_X1 port map( A1 => n9031, A2 => n9834, ZN => n9833);
   U4399 : NOR2_X1 port map( A1 => n9036, A2 => n9833, ZN => n9836);
   U4400 : AOI211_X1 port map( C1 => n9036, C2 => n9833, A => n9836, B => n9073
                           , ZN => n6810);
   U4401 : NAND2_X1 port map( A1 => n9032, A2 => n9836, ZN => n9835);
   U4402 : NOR2_X1 port map( A1 => n9034, A2 => n9835, ZN => n9837);
   U4403 : AOI211_X1 port map( C1 => n9034, C2 => n9835, A => n9837, B => n9073
                           , ZN => n6809);
   U4404 : AOI22_X1 port map( A1 => n5388, A2 => n9895, B1 => n9095, B2 => 
                           n9535, ZN => n6808);
   U4405 : INV_X1 port map( A => datapath_i_alu_output_val_i_31_port, ZN => 
                           n9783);
   U4406 : OAI222_X1 port map( A1 => n9562, A2 => n8950, B1 => n9783, B2 => 
                           n8993, C1 => n9081, C2 => n9053, ZN => n6772);
   U4407 : NAND3_X1 port map( A1 => n9203, A2 => n9105, A3 => n8725, ZN => 
                           n9784);
   U4408 : NOR2_X1 port map( A1 => n8723, A2 => n9784, ZN => n9796);
   U4409 : NOR2_X1 port map( A1 => n8645, A2 => n9106, ZN => n9795);
   U4410 : NAND2_X1 port map( A1 => n8725, A2 => n8732, ZN => n9790);
   U4411 : INV_X1 port map( A => n9796, ZN => n9802);
   U4412 : INV_X1 port map( A => n9784, ZN => n9785);
   U4413 : NAND3_X1 port map( A1 => n8723, A2 => n9785, A3 => n8646, ZN => 
                           n9803);
   U4414 : OAI211_X1 port map( C1 => n8646, C2 => n9790, A => n9802, B => n9803
                           , ZN => n9786);
   U4415 : AOI22_X1 port map( A1 => n9796, A2 => n8733, B1 => n9795, B2 => 
                           n9786, ZN => n9789);
   U4416 : NAND3_X1 port map( A1 => n9117, A2 => n9177, A3 => n9890, ZN => 
                           n9788);
   U4417 : NAND2_X1 port map( A1 => n9104, A2 => n8643, ZN => n9787);
   U4418 : NAND4_X1 port map( A1 => n8659, A2 => n9789, A3 => n9788, A4 => 
                           n9787, ZN => cu_i_N264);
   U4419 : NOR2_X1 port map( A1 => n9790, A2 => n9105, ZN => n9791);
   U4420 : AOI21_X1 port map( B1 => n9791, B2 => n9795, A => n8643, ZN => n9800
                           );
   U4421 : NOR3_X1 port map( A1 => n9174, A2 => n9200, A3 => n9803, ZN => n9794
                           );
   U4422 : NAND3_X1 port map( A1 => n8648, A2 => n9175, A3 => n9117, ZN => 
                           n9792);
   U4423 : NAND2_X1 port map( A1 => n9792, A2 => n8762, ZN => n9793);
   U4424 : AOI211_X1 port map( C1 => n9177, C2 => n9207, A => n9794, B => n9793
                           , ZN => n9798);
   U4425 : NAND3_X1 port map( A1 => n9796, A2 => n9795, A3 => n8646, ZN => 
                           n9797);
   U4426 : NAND3_X1 port map( A1 => n9800, A2 => n9798, A3 => n9797, ZN => 
                           cu_i_N265);
   U4427 : OAI221_X1 port map( B1 => n8733, B2 => n8646, C1 => n8733, C2 => 
                           n9106, A => n9200, ZN => n9801);
   U4428 : OAI221_X1 port map( B1 => n9175, B2 => n9104, C1 => n9175, C2 => 
                           n8647, A => n9207, ZN => n9799);
   U4429 : OAI211_X1 port map( C1 => n9802, C2 => n9801, A => n9800, B => n9799
                           , ZN => cu_i_N266);
   U4430 : OAI221_X1 port map( B1 => n9803, B2 => n8645, C1 => n9803, C2 => 
                           n9174, A => n9208, ZN => cu_i_N267);
   U4431 : NAND2_X1 port map( A1 => n9054, A2 => n8763, ZN => cu_i_N274);
   U4432 : AOI211_X1 port map( C1 => n9205, C2 => n9889, A => n8763, B => n9804
                           , ZN => cu_i_N275);
   U4433 : NOR2_X1 port map( A1 => n8763, A2 => n8779, ZN => cu_i_N273);
   U4434 : AOI211_X1 port map( C1 => n9204, C2 => n9806, A => n8763, B => n9805
                           , ZN => cu_i_N276);
   U4435 : AOI211_X1 port map( C1 => n9054, C2 => n8718, A => n8763, B => n9000
                           , ZN => cu_i_N279);
   U4436 : NOR2_X1 port map( A1 => n9807, A2 => n9548, ZN => n6932);
   U4437 : NOR2_X1 port map( A1 => n6900, A2 => n6898, ZN => n492);
   U4438 : NAND4_X1 port map( A1 => n9808, A2 => n6932, A3 => n492, A4 => n9549
                           , ZN => n9811);
   U4439 : NAND3_X1 port map( A1 => n9869, A2 => n9011, A3 => n9868, ZN => 
                           n9809);
   U4440 : OAI22_X1 port map( A1 => n9543, A2 => n9811, B1 => n9810, B2 => 
                           n9809, ZN => cu_i_cmd_word_8_port);
   U4441 : MUX2_X1 port map( A => n8704, B => cu_i_cmd_word_8_port, S => n5388,
                           Z => alu_cin_i);
   U4442 : MUX2_X1 port map( A => n8770, B => n8703, S => n5388, Z => n6879);
   U4443 : MUX2_X1 port map( A => n9101, B => n8702, S => n5388, Z => n6878);
   U4444 : MUX2_X1 port map( A => n8608, B => n8701, S => n5388, Z => n6877);
   U4445 : MUX2_X1 port map( A => IRAM_DATA(25), B => n8700, S => n8773, Z => 
                           n6876);
   U4446 : MUX2_X1 port map( A => IRAM_DATA(24), B => n8699, S => n8773, Z => 
                           n6875);
   U4447 : MUX2_X1 port map( A => IRAM_DATA(21), B => n8698, S => n9054, Z => 
                           n6874);
   U4448 : MUX2_X1 port map( A => IRAM_DATA(10), B => n8697, S => n8773, Z => 
                           n6873);
   U4449 : MUX2_X1 port map( A => IRAM_DATA(9), B => n8696, S => n8773, Z => 
                           n6872);
   U4450 : MUX2_X1 port map( A => IRAM_DATA(8), B => n8695, S => n8773, Z => 
                           n6871);
   U4451 : MUX2_X1 port map( A => IRAM_DATA(7), B => n8694, S => n8773, Z => 
                           n6870);
   U4452 : MUX2_X1 port map( A => IRAM_DATA(6), B => n8693, S => n8773, Z => 
                           n6869);
   U4453 : NOR2_X1 port map( A1 => n9584, A2 => n9526, ZN => n9813);
   U4454 : INV_X1 port map( A => n9815, ZN => n9812);
   U4455 : OAI211_X1 port map( C1 => n9813, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n9610, B => n9812, ZN => n6806);
   U4456 : OAI211_X1 port map( C1 => n9815, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n9610, B => n9814, ZN => n6805);
   U4457 : OAI211_X1 port map( C1 => n9817, C2 => n1453, A => n9610, B => n9816
                           , ZN => n6804);
   U4458 : OAI211_X1 port map( C1 => n9819, C2 => n1449, A => n9610, B => n9818
                           , ZN => n6803);
   U4459 : OAI211_X1 port map( C1 => n9821, C2 => n1447, A => n9610, B => n9820
                           , ZN => n6802);
   U4460 : OAI211_X1 port map( C1 => n9822, C2 => n1445, A => n9610, B => n6910
                           , ZN => n6801);
   U4461 : OAI211_X1 port map( C1 => n8735, C2 => IRAM_ADDRESS_14_port, A => 
                           n8734, B => n9052, ZN => n6800);
   U4462 : OAI211_X1 port map( C1 => n9824, C2 => IRAM_ADDRESS_16_port, A => 
                           n9052, B => n9823, ZN => n6799);
   U4463 : OAI211_X1 port map( C1 => n9826, C2 => IRAM_ADDRESS_18_port, A => 
                           n9052, B => n9825, ZN => n6798);
   U4464 : OAI211_X1 port map( C1 => n9828, C2 => IRAM_ADDRESS_20_port, A => 
                           n9052, B => n9827, ZN => n6797);
   U4465 : OAI211_X1 port map( C1 => n9830, C2 => IRAM_ADDRESS_22_port, A => 
                           n9052, B => n9829, ZN => n6796);
   U4466 : OAI211_X1 port map( C1 => n9832, C2 => IRAM_ADDRESS_24_port, A => 
                           n9052, B => n9831, ZN => n6795);
   U4467 : OAI211_X1 port map( C1 => n9834, C2 => IRAM_ADDRESS_26_port, A => 
                           n9052, B => n9833, ZN => n6794);
   U4468 : OAI211_X1 port map( C1 => n9836, C2 => IRAM_ADDRESS_28_port, A => 
                           n9052, B => n9835, ZN => n6793);
   U4469 : NAND2_X1 port map( A1 => n9033, A2 => n9837, ZN => n9838);
   U4470 : OAI211_X1 port map( C1 => n9837, C2 => IRAM_ADDRESS_30_port, A => 
                           n9052, B => n9838, ZN => n6792);
   U4471 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n9838, Z => n6908)
                           ;
   U4472 : AND2_X1 port map( A1 => n9095, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U4473 : OAI21_X1 port map( B1 => n9840, B2 => n9839, A => n9874, ZN => 
                           read_rf_p2_i);
   U4474 : OAI21_X1 port map( B1 => n9019, B2 => n9841, A => n9379, ZN => 
                           datapath_i_decode_stage_dp_n44);
   U4475 : OAI21_X1 port map( B1 => n9016, B2 => n9841, A => n9376, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U4476 : OAI21_X1 port map( B1 => n8933, B2 => n9841, A => n9375, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U4477 : OAI21_X1 port map( B1 => n8936, B2 => n9841, A => n9374, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U4478 : OAI21_X1 port map( B1 => n8939, B2 => n8945, A => n9373, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U4479 : OAI21_X1 port map( B1 => n8986, B2 => n9841, A => n9372, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U4480 : OAI21_X1 port map( B1 => n8942, B2 => n9841, A => n9371, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U4481 : OAI21_X1 port map( B1 => n9004, B2 => n9841, A => n9370, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U4482 : OAI21_X1 port map( B1 => n9076, B2 => n9841, A => n9369, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U4483 : OAI21_X1 port map( B1 => n9841, B2 => n9006, A => n9368, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U4484 : OAI21_X1 port map( B1 => n9841, B2 => n8748, A => n9367, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U4485 : OAI21_X1 port map( B1 => n8945, B2 => n8759, A => n9366, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U4486 : OAI21_X1 port map( B1 => n8945, B2 => n9069, A => n9365, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U4487 : OAI21_X1 port map( B1 => n9841, B2 => n8758, A => n9364, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U4488 : OAI21_X1 port map( B1 => n9841, B2 => n9108, A => n9363, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U4489 : OAI21_X1 port map( B1 => n8945, B2 => n8757, A => n9362, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U4490 : OAI21_X1 port map( B1 => n8945, B2 => n9114, A => n9361, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U4491 : OAI21_X1 port map( B1 => n9841, B2 => n8754, A => n9360, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U4492 : OAI21_X1 port map( B1 => n9841, B2 => n9112, A => n9359, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U4493 : OAI21_X1 port map( B1 => n8945, B2 => n8753, A => n9358, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U4494 : OAI21_X1 port map( B1 => n8945, B2 => n9103, A => n9357, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U4495 : OAI21_X1 port map( B1 => n9841, B2 => n8750, A => n9356, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U4496 : OAI21_X1 port map( B1 => n9841, B2 => n9097, A => n9355, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U4497 : OAI21_X1 port map( B1 => n8945, B2 => n8751, A => n9354, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U4498 : OAI21_X1 port map( B1 => n8945, B2 => n9094, A => n9353, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U4499 : OAI21_X1 port map( B1 => n9841, B2 => n8752, A => n9352, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U4500 : OAI21_X1 port map( B1 => n9841, B2 => n9090, A => n9351, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U4501 : OAI21_X1 port map( B1 => n8945, B2 => n8755, A => n9350, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U4502 : OAI21_X1 port map( B1 => n8945, B2 => n9086, A => n9349, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U4503 : OAI21_X1 port map( B1 => n9841, B2 => n8756, A => n9348, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U4504 : OAI21_X1 port map( B1 => n9841, B2 => n9084, A => n9347, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U4505 : OAI21_X1 port map( B1 => n8945, B2 => n9082, A => n9346, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U4506 : NOR4_X1 port map( A1 => n1641, A2 => n1643, A3 => n1645, A4 => n1647
                           , ZN => n9845);
   U4507 : NOR4_X1 port map( A1 => n1649, A2 => n1651, A3 => n1653, A4 => n1655
                           , ZN => n9844);
   U4508 : NOR4_X1 port map( A1 => n1625, A2 => n1627, A3 => n1629, A4 => n1631
                           , ZN => n9843);
   U4509 : NOR4_X1 port map( A1 => n1633, A2 => n1635, A3 => n1637, A4 => n1639
                           , ZN => n9842);
   U4510 : NAND4_X1 port map( A1 => n9845, A2 => n9844, A3 => n9843, A4 => 
                           n9842, ZN => n9851);
   U4511 : NOR4_X1 port map( A1 => n1663, A2 => n1617, A3 => n1619, A4 => n1621
                           , ZN => n9849);
   U4512 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1661
                           , ZN => n9848);
   U4513 : NOR4_X1 port map( A1 => n1667, A2 => n1669, A3 => n1657, A4 => n1659
                           , ZN => n9847);
   U4514 : NOR4_X1 port map( A1 => n1623, A2 => n1671, A3 => n1673, A4 => n1665
                           , ZN => n9846);
   U4515 : NAND4_X1 port map( A1 => n9849, A2 => n9848, A3 => n9847, A4 => 
                           n9846, ZN => n9850);
   U4516 : NOR2_X1 port map( A1 => n9851, A2 => n9850, ZN => n6907);
   U4517 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n9116, Z => n6868);
   U4518 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n9116, Z => n6867);
   U4519 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n9050, Z => n6866);
   U4520 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n9050, Z => n6865);
   U4521 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n9116, Z => n6864);
   U4522 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n9116, Z => n6863);
   U4523 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n9050, Z => n6862);
   U4524 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n9050, Z => n6861);
   U4525 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, S 
                           => n9116, Z => n6860);
   U4526 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, S 
                           => n9116, Z => n6859);
   U4527 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, S 
                           => n9050, Z => n6858);
   U4528 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, S 
                           => n9050, Z => n6857);
   U4529 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, S 
                           => n9116, Z => n6856);
   U4530 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, S 
                           => n9116, Z => n6855);
   U4531 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, S 
                           => n9050, Z => n6854);
   U4532 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, S 
                           => n9050, Z => n6853);
   U4533 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, S 
                           => n9116, Z => n6852);
   U4534 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, S 
                           => n9116, Z => n6851);
   U4535 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, S 
                           => n9050, Z => n6850);
   U4536 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, S 
                           => n9050, Z => n6849);
   U4537 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n9116, Z => n6848);
   U4538 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, S 
                           => n9116, Z => n6847);
   U4539 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, S 
                           => n9050, Z => n6846);
   U4540 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, S 
                           => n9050, Z => n6845);
   U4541 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, S 
                           => n9116, Z => n6844);
   U4542 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, S 
                           => n9116, Z => n6843);
   U4543 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n9050, Z => n6842);
   U4544 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n9116, Z => n6841);
   U4545 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n9116, Z => n6840);
   U4546 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n9116, Z => n6839);
   U4547 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n9116, Z => n6838);
   U4548 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n9116, Z => n6837);
   U4549 : MUX2_X1 port map( A => n8692, B => n8803, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U4550 : MUX2_X1 port map( A => n8691, B => n8806, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U4551 : MUX2_X1 port map( A => n8690, B => n8809, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U4552 : MUX2_X1 port map( A => n8689, B => n8812, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U4553 : MUX2_X1 port map( A => n8688, B => n8815, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U4554 : MUX2_X1 port map( A => n8687, B => n8818, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U4555 : MUX2_X1 port map( A => n8686, B => n8821, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U4556 : MUX2_X1 port map( A => n8685, B => n8824, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U4557 : MUX2_X1 port map( A => n8684, B => n8827, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U4558 : MUX2_X1 port map( A => n8683, B => n8830, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U4559 : MUX2_X1 port map( A => n8682, B => n8833, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U4560 : MUX2_X1 port map( A => n8681, B => n8836, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U4561 : MUX2_X1 port map( A => n8680, B => n8839, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U4562 : MUX2_X1 port map( A => n8679, B => n8842, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U4563 : MUX2_X1 port map( A => n8678, B => n8845, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U4564 : MUX2_X1 port map( A => n8677, B => n8848, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U4565 : MUX2_X1 port map( A => n8676, B => n8851, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U4566 : MUX2_X1 port map( A => n8675, B => n8854, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U4567 : MUX2_X1 port map( A => n8674, B => n8857, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U4568 : MUX2_X1 port map( A => n8673, B => n8860, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U4569 : MUX2_X1 port map( A => n8671, B => n8863, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U4570 : MUX2_X1 port map( A => n8670, B => n8866, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U4571 : MUX2_X1 port map( A => n8669, B => n8869, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U4572 : MUX2_X1 port map( A => n8668, B => n8872, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U4573 : MUX2_X1 port map( A => n8667, B => n8875, S => n8626, Z => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U4574 : MUX2_X1 port map( A => n8661, B => n8800, S => n9122, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U4575 : AOI22_X1 port map( A1 => n8743, A2 => n9593, B1 => n9013, B2 => 
                           n8901, ZN => n9852);
   U4576 : OAI21_X1 port map( B1 => n8742, B2 => n8973, A => n9852, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U4577 : AOI22_X1 port map( A1 => n8743, A2 => n9585, B1 => n9013, B2 => 
                           n8909, ZN => n9853);
   U4578 : OAI21_X1 port map( B1 => n8742, B2 => n8967, A => n9853, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U4579 : AOI22_X1 port map( A1 => n8743, A2 => n9854, B1 => n9013, B2 => 
                           n8911, ZN => n9855);
   U4580 : OAI21_X1 port map( B1 => n8742, B2 => n9096, A => n9855, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U4581 : AOI22_X1 port map( A1 => n8743, A2 => n9587, B1 => n9013, B2 => 
                           n8913, ZN => n9856);
   U4582 : OAI21_X1 port map( B1 => n8742, B2 => n8964, A => n9856, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U4583 : INV_X1 port map( A => n7852, ZN => n9857);
   U4584 : AOI22_X1 port map( A1 => n9531, A2 => n8877, B1 => n6919, B2 => 
                           n9857, ZN => n9858);
   U4585 : OAI21_X1 port map( B1 => n9019, B2 => n6920, A => n9858, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U4586 : AOI22_X1 port map( A1 => n8743, A2 => n9595, B1 => n9013, B2 => 
                           n8921, ZN => n9859);
   U4587 : OAI21_X1 port map( B1 => n8742, B2 => n8958, A => n9859, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U4588 : AOI22_X1 port map( A1 => n9860, A2 => n8743, B1 => n9013, B2 => 
                           n8929, ZN => n9861);
   U4589 : OAI21_X1 port map( B1 => n9081, B2 => n8742, A => n9861, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U4590 : INV_X1 port map( A => n9526, ZN => n9863);
   U4591 : AOI22_X1 port map( A1 => n9584, A2 => n9863, B1 => n9526, B2 => 
                           n9862, ZN => n6791);
   U4592 : AOI22_X1 port map( A1 => n9531, A2 => n8879, B1 => n6919, B2 => 
                           n9864, ZN => n9865);
   U4593 : OAI21_X1 port map( B1 => n8933, B2 => n6920, A => n9865, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U4594 : AOI22_X1 port map( A1 => n9531, A2 => n8880, B1 => n6919, B2 => 
                           n9866, ZN => n9867);
   U4595 : OAI21_X1 port map( B1 => n8936, B2 => n6920, A => n9867, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U4596 : MUX2_X1 port map( A => n8701, B => n8660, S => n5388, Z => n6836);
   U4597 : OAI211_X1 port map( C1 => n9550, C2 => n9605, A => n9869, B => n9868
                           , ZN => n6790);
   U4598 : MUX2_X1 port map( A => n9022, B => n8658, S => n5388, Z => n6835);
   U4599 : INV_X1 port map( A => curr_instruction_to_cu_i_17_port, ZN => n9871)
                           ;
   U4600 : OAI221_X1 port map( B1 => n9876, B2 => n9871, C1 => n9874, C2 => 
                           n9870, A => n9872, ZN => n9523);
   U4601 : OAI221_X1 port map( B1 => n9876, B2 => n9875, C1 => n9874, C2 => 
                           n9873, A => n9872, ZN => n4953);
   U4602 : NAND4_X1 port map( A1 => n9523, A2 => n9524, A3 => n9525, A4 => 
                           n4953, ZN => n9877);
   U4603 : NOR2_X1 port map( A1 => n9878, A2 => n9877, ZN => n9168);
   U4604 : OAI211_X1 port map( C1 => n9880, C2 => n1447, A => n9073, B => n9879
                           , ZN => n9881);
   U4605 : NAND2_X1 port map( A1 => n8621, A2 => n9881, ZN => n9178);
   U4606 : NOR2_X1 port map( A1 => n8728, A2 => n4052, ZN => n9182);
   U4607 : AOI222_X1 port map( A1 => n9599, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_15_port, B2 => n8951, C1
                           => n8989, C2 => n8974, ZN => n9600);
   U4608 : AOI222_X1 port map( A1 => n9597, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_29_port, B2 => n8951, C1
                           => n8989, C2 => n8953, ZN => n9598);
   U4609 : AOI222_X1 port map( A1 => n9595, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_27_port, B2 => n8951, C1
                           => n8989, C2 => n8956, ZN => n9596);
   U4610 : AOI222_X1 port map( A1 => n9593, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_17_port, B2 => n8951, C1
                           => n8989, C2 => n8971, ZN => n9594);
   U4611 : AOI222_X1 port map( A1 => n9591, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_19_port, B2 => n8951, C1
                           => n8989, C2 => n8968, ZN => n9592);
   U4612 : AOI222_X1 port map( A1 => n9589, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_25_port, B2 => n8951, C1
                           => n8989, C2 => n8959, ZN => n9590);
   U4613 : AOI222_X1 port map( A1 => n9587, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_23_port, B2 => n8951, C1
                           => n8989, C2 => n8962, ZN => n9588);
   U4614 : AOI222_X1 port map( A1 => n9585, A2 => n9886, B1 => 
                           datapath_i_alu_output_val_i_21_port, B2 => n8951, C1
                           => n8989, C2 => n8965, ZN => n9586);
   U4615 : AOI22_X1 port map( A1 => n5388, A2 => n8649, B1 => n8766, B2 => 
                           n9535, ZN => n9536);

end SYN_dlx_rtl;
