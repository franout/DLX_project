--------------------------------------------------------------------------------
-- Title       : execute stage of datapath
-- Project     : DLX for Microelectronic Systems
--------------------------------------------------------------------------------
-- File        : a.b.c-Execute.stage.vhd
-- Author      : Francesco Angione <s262620@studenti.polito.it>
-- Company     : Politecnico di Torino, Italy
-- Created     : Wed Jul 22 20:59:12 2020
-- Last update : Wed Jul 22 20:59:20 2020
-- Platform    : Default Part Number
-- Standard    : VHDL-2008 
--------------------------------------------------------------------------------
-- Copyright (c) 2020 Politecnico di Torino, Italy
-------------------------------------------------------------------------------
-- Description: 
--------------------------------------------------------------------------------

library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity execute_stage is
  port (
	clock
  ) ;
end entity ; -- execute_stage

architecture arch of execute_stage is

begin

end architecture ; -- arch