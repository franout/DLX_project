
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, 
      boothmul_pipelined_i_muxes_in_7_233_port, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_1_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_7_15_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n3076, 
      n3077, n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
      n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
      n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n_1004, n_1005, 
      n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, 
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, 
      n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, 
      n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, 
      n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, 
      n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, 
      n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, 
      n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, 
      n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, 
      n_1348 : std_logic;

begin
   
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n5140, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n5140, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n5139, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n5139, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n5139, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n5140, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n5139, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n5139, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n5140, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n5139, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n5140, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n5139, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n5140, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n5140, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n5140, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n5139, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n5140, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n5140, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n5140, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n5139, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n5140, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n5140, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n5140, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n5140, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n5140, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n5139, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n5139, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n5140, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n5139, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n5139, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => n5138, GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => n5137, GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => n5136, GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => n5135, GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, QN 
                           => n5125);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => n3111, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => n3103, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => n3105, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => n3107, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => n3107, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3080);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => n3112, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => n3108, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => n3111, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => n3113, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => n3110, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => n3104, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3079);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => n3105, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => n3105, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => n3105, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => n3101, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => n3111, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => n3101, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3078);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => n3104, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => n3108, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => n3109, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => n3110, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => n3113, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => n3115, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => n3105, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => n3104, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => n3109, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3082);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => n3113, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => n3103, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => n3101, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => n3115, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => n3108, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => n3104, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => n3108, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => n3112, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => n3109, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => n3108, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => n3103, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3076);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => n3103, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => n3113, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => n3108, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => n3104, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => n3113, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => n3104, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => n3104, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => n3111, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => n3101, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => n3115, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => n3107, Q => n_1060, QN => n5126);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => n3101, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3095, CK => clk, RN => rst_BAR, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => n3107, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => n3112, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => n3106, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => n3113, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => n3113, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => n3101, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => n3113, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => n3109, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => n3109, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => n3111, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => n3113, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => n3113, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_7_233_port, QN => 
                           n5134);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1106);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => n3108, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => n3115, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => n3106, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => n3111, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => n3109, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => n3103, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => n3106, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => n3114, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => n3107, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => n3106, Q => n_1120, QN => n5133);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => n3107, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1121
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3094, CK => clk, RN => n3115, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1122
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => n3113, Q => boothmul_pipelined_i_sum_out_6_9_port
                           , QN => n_1123);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => n3103, Q => boothmul_pipelined_i_sum_out_6_8_port
                           , QN => n_1124);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => n3115, Q => boothmul_pipelined_i_sum_out_6_7_port
                           , QN => n_1125);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => n3111, Q => boothmul_pipelined_i_sum_out_6_6_port
                           , QN => n_1126);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => n3107, Q => boothmul_pipelined_i_sum_out_6_5_port
                           , QN => n_1127);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => n3101, Q => boothmul_pipelined_i_sum_out_6_4_port
                           , QN => n_1128);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_3_port, QN => n_1129)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => n3107, Q => boothmul_pipelined_i_sum_out_6_2_port
                           , QN => n_1130);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => n3111, Q => boothmul_pipelined_i_sum_out_6_1_port
                           , QN => n_1131);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => n3112, Q => boothmul_pipelined_i_sum_out_6_0_port
                           , QN => n_1132);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => n5129
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1133);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => n5123
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1156);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1157);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1158);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1159);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1160);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1161);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1162);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => n3108, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1163);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1164);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => n3114, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1165);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1166);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => n3103, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1167);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => n3112, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => n3109, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => n3109, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => n3103, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => n3113, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => n3102, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => n3113, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => n3102, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => n3108, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => n3114, Q => n_1177, QN => n5132);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => n3110, Q => boothmul_pipelined_i_sum_out_5_9_port
                           , QN => n_1178);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3093, CK => clk, RN => n3101, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1179)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => n3104, Q => boothmul_pipelined_i_sum_out_5_7_port
                           , QN => n_1180);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_6_port, QN => n_1181)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => n3114, Q => boothmul_pipelined_i_sum_out_5_5_port
                           , QN => n_1182);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => n3106, Q => boothmul_pipelined_i_sum_out_5_4_port
                           , QN => n_1183);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => n3114, Q => boothmul_pipelined_i_sum_out_5_3_port
                           , QN => n_1184);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => n3112, Q => boothmul_pipelined_i_sum_out_5_2_port
                           , QN => n_1185);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => n3109, Q => boothmul_pipelined_i_sum_out_5_1_port
                           , QN => n_1186);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => n3107, Q => boothmul_pipelined_i_sum_out_5_0_port
                           , QN => n_1187);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => n5128
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1188);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1189);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1190);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1191);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n5122);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => n3108, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => n3111, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => n3114, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => n3108, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => n3102, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => n3101, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => n3109, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => n3101, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => n3101, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => n3104, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1231
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => n3107, Q => n_1232, QN => n5131);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => n3114, Q => boothmul_pipelined_i_sum_out_4_7_port
                           , QN => n_1233);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3092, CK => clk, RN => n3110, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1234)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => n3111, Q => boothmul_pipelined_i_sum_out_4_5_port
                           , QN => n_1235);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => n3107, Q => boothmul_pipelined_i_sum_out_4_4_port
                           , QN => n_1236);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => n3107, Q => boothmul_pipelined_i_sum_out_4_3_port
                           , QN => n_1237);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => n3101, Q => boothmul_pipelined_i_sum_out_4_2_port
                           , QN => n_1238);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => n3104, Q => boothmul_pipelined_i_sum_out_4_1_port
                           , QN => n_1239);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => n3112, Q => boothmul_pipelined_i_sum_out_4_0_port
                           , QN => n_1240);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => n5127
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1241);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1242);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1243);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1244);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1245);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1246);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1249);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1250);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1251);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1252);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1253);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1254);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => n5121
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1255);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => n3103, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1256);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1257);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1258);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => n3110, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => n3103, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => n3107, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => n3102, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => n3113, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => n3109, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => n3112, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => n3104, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1282
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1283
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => n3114, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1284
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => n3110, Q => n_1285, QN => n5124);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => n3102, Q => boothmul_pipelined_i_sum_out_3_5_port
                           , QN => n_1286);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3091, CK => clk, RN => n3112, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1287)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => n3106, Q => boothmul_pipelined_i_sum_out_3_3_port
                           , QN => n_1288);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => n3109, Q => boothmul_pipelined_i_sum_out_3_2_port
                           , QN => n_1289);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => n3114, Q => boothmul_pipelined_i_sum_out_3_1_port
                           , QN => n_1290);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => n3114, Q => boothmul_pipelined_i_sum_out_3_0_port
                           , QN => n_1291);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => 
                           n_1292);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => n3108, Q => 
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1293);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1294);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1295);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1296);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1297);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1298);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => n3106, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => n3114, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => n3107, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => n3115, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => n3104, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => n3113, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => n3111, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => n3109, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => n3105, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => n3112, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => n3102, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => n3113, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => n3115, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => n3105, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => n3114, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => n3112, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => n3110, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => n3114, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => n3111, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1332
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => n3107, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1333
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1334
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => n3103, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1335
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => n3107, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1336
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => n3104, Q => n_1337, QN => n5130);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => n3114, Q => boothmul_pipelined_i_sum_out_2_3_port
                           , QN => n_1338);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3086, CK => clk, RN => n3102, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1339)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_1_port, CK => clk, RN
                           => n3109, Q => boothmul_pipelined_i_sum_out_2_1_port
                           , QN => n_1340);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => n3108, Q => boothmul_pipelined_i_sum_out_2_0_port
                           , QN => n_1341);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => n3101, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n3077);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n5140, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1993, B => n1994, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1992, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1991, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1990, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1989, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1988, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1987, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1986, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1985, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1984, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1983, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1982, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1981, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1980, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1979, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3083,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1342, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3085,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1343, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3084,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n1998, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1344, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3090,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n1997, B => boothmul_pipelined_i_sum_B_in_4_24_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1345, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3089
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n1996, B => boothmul_pipelined_i_sum_B_in_5_26_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1346, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3088
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n1995, B => boothmul_pipelined_i_sum_B_in_6_28_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1347, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3087
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1348, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n5140, Q => 
                           DATA2_I_30_port);
   U3 : CLKBUF_X1 port map( A => n3104, Z => n3101);
   U4 : CLKBUF_X1 port map( A => n3104, Z => n3102);
   U5 : CLKBUF_X1 port map( A => n3104, Z => n3103);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n3104);
   U7 : CLKBUF_X1 port map( A => n3108, Z => n3105);
   U8 : CLKBUF_X1 port map( A => n3101, Z => n3106);
   U9 : CLKBUF_X1 port map( A => n3102, Z => n3107);
   U10 : CLKBUF_X1 port map( A => n3102, Z => n3108);
   U11 : CLKBUF_X1 port map( A => n3102, Z => n3109);
   U12 : CLKBUF_X1 port map( A => n3102, Z => n3110);
   U13 : CLKBUF_X1 port map( A => n3103, Z => n3111);
   U14 : CLKBUF_X1 port map( A => n3103, Z => n3112);
   U15 : CLKBUF_X1 port map( A => n3103, Z => n3113);
   U16 : CLKBUF_X1 port map( A => n3103, Z => n3114);
   U17 : CLKBUF_X1 port map( A => n3103, Z => n3115);
   U18 : NOR2_X2 port map( A1 => DATA2(4), A2 => DATA2(5), ZN => n4555);
   U19 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => n4834, ZN => n3135);
   U20 : CLKBUF_X1 port map( A => n4832, Z => n4822);
   U21 : NOR2_X1 port map( A1 => FUNC(1), A2 => FUNC(0), ZN => n3147);
   U22 : INV_X1 port map( A => FUNC(2), ZN => n4724);
   U23 : AND2_X1 port map( A1 => n3147, A2 => n4724, ZN => n4797);
   U24 : INV_X1 port map( A => n4797, ZN => n5140);
   U25 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n3116);
   U26 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, A
                           => n3116, ZN => n3140);
   U27 : NOR2_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_3_7_port
                           , A2 => n3140, ZN => n4952);
   U28 : CLKBUF_X1 port map( A => n4952, Z => n4946);
   U29 : NAND3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n4919);
   U30 : INV_X1 port map( A => n4919, ZN => n4950);
   U31 : NOR3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n4949);
   U32 : NOR2_X1 port map( A1 => n3082, A2 => n3140, ZN => n4932);
   U33 : CLKBUF_X1 port map( A => n4932, Z => n4951);
   U34 : AOI22_X1 port map( A1 => n4949, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, B1 => 
                           n4951, B2 => 
                           boothmul_pipelined_i_muxes_in_3_161_port, ZN => 
                           n3117);
   U35 : INV_X1 port map( A => n3117, ZN => n3118);
   U36 : AOI221_X1 port map( B1 => boothmul_pipelined_i_muxes_in_3_46_port, B2 
                           => n4946, C1 => 
                           boothmul_pipelined_i_muxes_in_3_46_port, C2 => n4950
                           , A => n3118, ZN => n3119);
   U37 : INV_X1 port map( A => n3119, ZN => n1998);
   U38 : INV_X1 port map( A => data1_mul_0_port, ZN => n1994);
   U39 : AND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n5102);
   U40 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n4834);
   U41 : CLKBUF_X1 port map( A => n3135, Z => n3132);
   U42 : AND2_X1 port map( A1 => n4834, A2 => data2_mul_1_port, ZN => n5103);
   U43 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, A2
                           => n5102, B1 => data1_mul_14_port, B2 => n3132, C1 
                           => boothmul_pipelined_i_muxes_in_0_104_port, C2 => 
                           n5103, ZN => n3120);
   U44 : INV_X1 port map( A => n3120, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U45 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, A2
                           => n5102, B1 => data1_mul_13_port, B2 => n3135, C1 
                           => boothmul_pipelined_i_muxes_in_0_105_port, C2 => 
                           n5103, ZN => n3121);
   U46 : INV_X1 port map( A => n3121, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U47 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, A2
                           => n5102, B1 => data1_mul_12_port, B2 => n3135, C1 
                           => boothmul_pipelined_i_muxes_in_0_106_port, C2 => 
                           n5103, ZN => n3122);
   U48 : INV_X1 port map( A => n3122, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U49 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, A2
                           => n5102, B1 => data1_mul_11_port, B2 => n3132, C1 
                           => boothmul_pipelined_i_muxes_in_0_107_port, C2 => 
                           n5103, ZN => n3123);
   U50 : INV_X1 port map( A => n3123, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U51 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, A2
                           => n5102, B1 => data1_mul_10_port, B2 => n3132, C1 
                           => boothmul_pipelined_i_muxes_in_0_108_port, C2 => 
                           n5103, ZN => n3124);
   U52 : INV_X1 port map( A => n3124, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U53 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, A2
                           => n5102, B1 => data1_mul_9_port, B2 => n3135, C1 =>
                           boothmul_pipelined_i_muxes_in_0_109_port, C2 => 
                           n5103, ZN => n3125);
   U54 : INV_X1 port map( A => n3125, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U55 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, A2
                           => n5102, B1 => data1_mul_8_port, B2 => n3132, C1 =>
                           boothmul_pipelined_i_muxes_in_0_110_port, C2 => 
                           n5103, ZN => n3126);
   U56 : INV_X1 port map( A => n3126, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U57 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, A2
                           => n5102, B1 => data1_mul_7_port, B2 => n3135, C1 =>
                           boothmul_pipelined_i_muxes_in_0_111_port, C2 => 
                           n5103, ZN => n3127);
   U58 : INV_X1 port map( A => n3127, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U59 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, A2
                           => n5102, B1 => data1_mul_6_port, B2 => n3135, C1 =>
                           boothmul_pipelined_i_muxes_in_0_112_port, C2 => 
                           n5103, ZN => n3128);
   U60 : INV_X1 port map( A => n3128, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U61 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, A2
                           => n5102, B1 => data1_mul_5_port, B2 => n3132, C1 =>
                           boothmul_pipelined_i_muxes_in_0_113_port, C2 => 
                           n5103, ZN => n3129);
   U62 : INV_X1 port map( A => n3129, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U63 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, A2
                           => n5102, B1 => data1_mul_4_port, B2 => n3132, C1 =>
                           boothmul_pipelined_i_muxes_in_0_114_port, C2 => 
                           n5103, ZN => n3130);
   U64 : INV_X1 port map( A => n3130, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U65 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, A2
                           => n5102, B1 => data1_mul_3_port, B2 => n3132, C1 =>
                           boothmul_pipelined_i_muxes_in_0_115_port, C2 => 
                           n5103, ZN => n3131);
   U66 : INV_X1 port map( A => n3131, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U67 : AOI222_X1 port map( A1 => n5102, A2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B1 => 
                           data1_mul_1_port, B2 => n3132, C1 => 
                           data1_mul_0_port, C2 => n5103, ZN => n3133);
   U68 : INV_X1 port map( A => n3133, ZN => 
                           boothmul_pipelined_i_sum_out_1_1_port);
   U69 : CLKBUF_X1 port map( A => DATA1(4), Z => n5136);
   U70 : CLKBUF_X1 port map( A => DATA1(14), Z => n5138);
   U71 : CLKBUF_X1 port map( A => DATA1(10), Z => n5137);
   U72 : CLKBUF_X1 port map( A => DATA1(3), Z => n5135);
   U73 : INV_X1 port map( A => n4797, ZN => n5139);
   U74 : INV_X1 port map( A => data1_mul_15_port, ZN => n1979);
   U75 : XNOR2_X1 port map( A => data1_mul_15_port, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
                           ZN => boothmul_pipelined_i_muxes_in_0_119_port);
   U76 : INV_X1 port map( A => n3135, ZN => n5105);
   U77 : AOI22_X1 port map( A1 => n5103, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n5102, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n3134);
   U78 : OAI21_X1 port map( B1 => n5105, B2 => n1979, A => n3134, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U79 : INV_X1 port map( A => data1_mul_14_port, ZN => n1980);
   U80 : INV_X1 port map( A => data1_mul_13_port, ZN => n1981);
   U81 : INV_X1 port map( A => data1_mul_12_port, ZN => n1982);
   U82 : INV_X1 port map( A => data1_mul_11_port, ZN => n1983);
   U83 : INV_X1 port map( A => data1_mul_10_port, ZN => n1984);
   U84 : INV_X1 port map( A => data1_mul_9_port, ZN => n1985);
   U85 : INV_X1 port map( A => data1_mul_8_port, ZN => n1986);
   U86 : INV_X1 port map( A => data1_mul_7_port, ZN => n1987);
   U87 : INV_X1 port map( A => data1_mul_6_port, ZN => n1988);
   U88 : INV_X1 port map( A => data1_mul_5_port, ZN => n1989);
   U89 : INV_X1 port map( A => data1_mul_4_port, ZN => n1990);
   U90 : INV_X1 port map( A => data1_mul_3_port, ZN => n1991);
   U91 : INV_X1 port map( A => data1_mul_2_port, ZN => n1992);
   U92 : INV_X1 port map( A => data1_mul_1_port, ZN => n1993);
   U93 : AOI222_X1 port map( A1 => n3135, A2 => data1_mul_2_port, B1 => n5103, 
                           B2 => boothmul_pipelined_i_muxes_in_0_116_port, C1 
                           => n5102, C2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, ZN => 
                           n3137);
   U94 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n4875);
   U95 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n4875, ZN => n4835);
   U96 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n4835, ZN => n3136);
   U97 : NOR2_X1 port map( A1 => n3137, A2 => n3136, ZN => n3083);
   U98 : AOI21_X1 port map( B1 => n3137, B2 => n3136, A => n3083, ZN => n3086);
   U99 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n3138);
   U100 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n3138, ZN => n4877);
   U101 : NOR3_X1 port map( A1 => n1994, A2 => n4877, A3 => n5130, ZN => n3085)
                           ;
   U102 : OR2_X1 port map( A1 => n1994, A2 => n4877, ZN => n3139);
   U103 : AOI21_X1 port map( B1 => n3139, B2 => n5130, A => n3085, ZN => n3091)
                           ;
   U104 : NOR3_X1 port map( A1 => n3077, A2 => n3140, A3 => n5124, ZN => n3084)
                           ;
   U105 : AOI221_X1 port map( B1 => n3077, B2 => n5124, C1 => n3140, C2 => 
                           n5124, A => n3084, ZN => n3092);
   U106 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n3141);
   U107 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, A
                           => n3141, ZN => n4956);
   U108 : NOR3_X1 port map( A1 => n4956, A2 => n5121, A3 => n5131, ZN => n3090)
                           ;
   U109 : INV_X1 port map( A => n4956, ZN => n4955);
   U110 : NAND2_X1 port map( A1 => n4955, A2 => 
                           boothmul_pipelined_i_muxes_in_4_65_port, ZN => n3142
                           );
   U111 : AOI21_X1 port map( B1 => n3142, B2 => n5131, A => n3090, ZN => n3093)
                           ;
   U112 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n3143);
   U113 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           A => n3143, ZN => n4992);
   U114 : NOR3_X1 port map( A1 => n4992, A2 => n5122, A3 => n5132, ZN => n3089)
                           ;
   U115 : INV_X1 port map( A => n4992, ZN => n4991);
   U116 : NAND2_X1 port map( A1 => n4991, A2 => 
                           boothmul_pipelined_i_muxes_in_5_205_port, ZN => 
                           n3144);
   U117 : AOI21_X1 port map( B1 => n3144, B2 => n5132, A => n3089, ZN => n3094)
                           ;
   U118 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n3145);
   U119 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           A => n3145, ZN => n5028);
   U120 : NOR3_X1 port map( A1 => n5028, A2 => n5123, A3 => n5133, ZN => n3088)
                           ;
   U121 : INV_X1 port map( A => n5028, ZN => n5027);
   U122 : NAND2_X1 port map( A1 => n5027, A2 => 
                           boothmul_pipelined_i_muxes_in_6_73_port, ZN => n3146
                           );
   U123 : AOI21_X1 port map( B1 => n3146, B2 => n5133, A => n3088, ZN => n3095)
                           ;
   U124 : NOR2_X1 port map( A1 => FUNC(3), A2 => n4724, ZN => n4770);
   U125 : NAND2_X1 port map( A1 => n4770, A2 => n3147, ZN => n553);
   U126 : INV_X1 port map( A => DATA1(9), ZN => n3617);
   U127 : NOR2_X1 port map( A1 => DATA2(9), A2 => n3617, ZN => n4613);
   U128 : INV_X1 port map( A => n4613, ZN => n4679);
   U129 : NAND2_X1 port map( A1 => DATA2(9), A2 => n3617, ZN => n4674);
   U130 : AND2_X1 port map( A1 => n4679, A2 => n4674, ZN => n4768);
   U131 : INV_X1 port map( A => FUNC(0), ZN => n4773);
   U132 : NAND2_X1 port map( A1 => n4773, A2 => FUNC(1), ZN => n3174);
   U133 : NOR2_X1 port map( A1 => FUNC(2), A2 => n3174, ZN => n4778);
   U134 : CLKBUF_X1 port map( A => n4778, Z => n4372);
   U135 : INV_X1 port map( A => n4372, ZN => n4479);
   U136 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(8), A3 => DATA2(6), A4 
                           => DATA2(7), ZN => n3155);
   U137 : INV_X1 port map( A => DATA2(3), ZN => n4828);
   U138 : NAND2_X1 port map( A1 => n4555, A2 => n4828, ZN => n3167);
   U139 : INV_X1 port map( A => n3167, ZN => n3169);
   U140 : INV_X1 port map( A => DATA2(2), ZN => n4829);
   U141 : AND2_X1 port map( A1 => n3169, A2 => n4829, ZN => n3658);
   U142 : NOR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n3510);
   U143 : NAND2_X1 port map( A1 => n3658, A2 => n3510, ZN => n4248);
   U144 : INV_X1 port map( A => DATA2(12), ZN => n4817);
   U145 : INV_X1 port map( A => DATA2(10), ZN => n4819);
   U146 : INV_X1 port map( A => DATA2(11), ZN => n4818);
   U147 : INV_X1 port map( A => DATA2(13), ZN => n4816);
   U148 : NAND4_X1 port map( A1 => n4817, A2 => n4819, A3 => n4818, A4 => n4816
                           , ZN => n3148);
   U149 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n4248, A4 
                           => n3148, ZN => n3154);
   U150 : NOR4_X1 port map( A1 => DATA1(13), A2 => DATA1(12), A3 => DATA1(11), 
                           A4 => DATA1(10), ZN => n3152);
   U151 : NOR4_X1 port map( A1 => DATA1(15), A2 => n5138, A3 => DATA1(9), A4 =>
                           DATA1(7), ZN => n3151);
   U152 : CLKBUF_X1 port map( A => DATA1(8), Z => n3619);
   U153 : NOR4_X1 port map( A1 => n3619, A2 => DATA1(6), A3 => DATA1(5), A4 => 
                           n5136, ZN => n3150);
   U154 : CLKBUF_X1 port map( A => DATA1(0), Z => n4780);
   U155 : NOR4_X1 port map( A1 => DATA1(3), A2 => DATA1(2), A3 => DATA1(1), A4 
                           => n4780, ZN => n3149);
   U156 : AND4_X1 port map( A1 => n3152, A2 => n3151, A3 => n3150, A4 => n3149,
                           ZN => n3153);
   U157 : AOI211_X1 port map( C1 => n3155, C2 => n3154, A => n3153, B => n553, 
                           ZN => n4476);
   U158 : INV_X1 port map( A => n4476, ZN => n4403);
   U159 : INV_X1 port map( A => n4403, ZN => n4491);
   U160 : NAND2_X1 port map( A1 => FUNC(3), A2 => FUNC(2), ZN => n3156);
   U161 : NOR3_X1 port map( A1 => FUNC(1), A2 => FUNC(0), A3 => n3156, ZN => 
                           n4781);
   U162 : CLKBUF_X1 port map( A => n4781, Z => n4510);
   U163 : INV_X1 port map( A => n4510, ZN => n4471);
   U164 : INV_X1 port map( A => FUNC(3), ZN => n4796);
   U165 : NAND2_X1 port map( A1 => n4778, A2 => n4796, ZN => n4470);
   U166 : NAND2_X1 port map( A1 => n4471, A2 => n4470, ZN => n4450);
   U167 : INV_X1 port map( A => n4450, ZN => n4111);
   U168 : INV_X1 port map( A => DATA2(9), ZN => n4820);
   U169 : NOR3_X1 port map( A1 => n4111, A2 => n4820, A3 => n3617, ZN => n3178)
                           ;
   U170 : INV_X1 port map( A => n4555, ZN => n4028);
   U171 : NOR2_X1 port map( A1 => DATA2(2), A2 => n4028, ZN => n3194);
   U172 : NAND3_X1 port map( A1 => DATA2(3), A2 => n3194, A3 => n3510, ZN => 
                           n4531);
   U173 : INV_X1 port map( A => n4531, ZN => n4160);
   U174 : CLKBUF_X1 port map( A => n4160, Z => n4196);
   U175 : INV_X1 port map( A => DATA2(1), ZN => n4830);
   U176 : OAI21_X1 port map( B1 => n4829, B2 => n4830, A => n3169, ZN => n4529)
                           ;
   U177 : INV_X1 port map( A => n4529, ZN => n3852);
   U178 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(0), ZN => n3192);
   U179 : AND2_X1 port map( A1 => n3852, A2 => n3192, ZN => n4527);
   U180 : INV_X1 port map( A => n4527, ZN => n4113);
   U181 : CLKBUF_X1 port map( A => n3658, Z => n4255);
   U182 : INV_X1 port map( A => n4255, ZN => n4009);
   U183 : INV_X1 port map( A => DATA1(7), ZN => n3471);
   U184 : NOR2_X1 port map( A1 => n4248, A2 => n3471, ZN => n3158);
   U185 : INV_X1 port map( A => DATA2(0), ZN => n4831);
   U186 : NOR2_X1 port map( A1 => n4831, A2 => DATA2(1), ZN => n3949);
   U187 : NAND2_X1 port map( A1 => n4255, A2 => n3949, ZN => n4242);
   U188 : INV_X1 port map( A => n4242, ZN => n4074);
   U189 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(6), ZN => n3433);
   U190 : OR3_X1 port map( A1 => DATA2(0), A2 => n4830, A3 => n4009, ZN => 
                           n4007);
   U191 : INV_X1 port map( A => n4007, ZN => n4520);
   U192 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(5), ZN => n3512);
   U193 : NOR2_X1 port map( A1 => n4830, A2 => n4831, ZN => n3454);
   U194 : NAND2_X1 port map( A1 => n3454, A2 => n3658, ZN => n4077);
   U195 : INV_X1 port map( A => n4077, ZN => n3785);
   U196 : CLKBUF_X1 port map( A => n3785, Z => n3810);
   U197 : NAND2_X1 port map( A1 => n3810, A2 => DATA1(4), ZN => n4253);
   U198 : NAND3_X1 port map( A1 => n3433, A2 => n3512, A3 => n4253, ZN => n3157
                           );
   U199 : AOI211_X1 port map( C1 => n5135, C2 => n4009, A => n3158, B => n3157,
                           ZN => n3168);
   U200 : NAND4_X1 port map( A1 => DATA2(2), A2 => DATA2(0), A3 => n3169, A4 =>
                           n4830, ZN => n3768);
   U201 : INV_X1 port map( A => n3768, ZN => n4525);
   U202 : INV_X1 port map( A => n4525, ZN => n4115);
   U203 : INV_X1 port map( A => n4248, ZN => n4258);
   U204 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(6), ZN => n3399);
   U205 : INV_X1 port map( A => n3399, ZN => n3160);
   U206 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(5), ZN => n3472);
   U207 : INV_X1 port map( A => n4007, ZN => n4073);
   U208 : NAND2_X1 port map( A1 => n4073, A2 => n5136, ZN => n4010);
   U209 : NAND2_X1 port map( A1 => n3810, A2 => n5135, ZN => n4522);
   U210 : NAND3_X1 port map( A1 => n3472, A2 => n4010, A3 => n4522, ZN => n3159
                           );
   U211 : AOI211_X1 port map( C1 => DATA1(2), C2 => n4009, A => n3160, B => 
                           n3159, ZN => n3173);
   U212 : INV_X1 port map( A => DATA1(5), ZN => n4254);
   U213 : NOR2_X1 port map( A1 => n4248, A2 => n4254, ZN => n3162);
   U214 : INV_X1 port map( A => DATA1(2), ZN => n4008);
   U215 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(4), ZN => n3514);
   U216 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(3), ZN => n4252);
   U217 : OAI211_X1 port map( C1 => n4077, C2 => n4008, A => n3514, B => n4252,
                           ZN => n3161);
   U218 : AOI211_X1 port map( C1 => DATA1(1), C2 => n4009, A => n3162, B => 
                           n3161, ZN => n3455);
   U219 : CLKBUF_X1 port map( A => n3852, Z => n3900);
   U220 : OAI222_X1 port map( A1 => n4113, A2 => n3168, B1 => n4115, B2 => 
                           n3173, C1 => n3455, C2 => n3900, ZN => n3965);
   U221 : CLKBUF_X1 port map( A => n4529, Z => n4260);
   U222 : OAI21_X1 port map( B1 => DATA2(0), B2 => n3167, A => n4260, ZN => 
                           n4193);
   U223 : INV_X1 port map( A => n4527, ZN => n3871);
   U224 : CLKBUF_X1 port map( A => n4258, Z => n4519);
   U225 : NOR2_X1 port map( A1 => n4007, A2 => n3471, ZN => n3435);
   U226 : NOR2_X1 port map( A1 => n4255, A2 => n4254, ZN => n3163);
   U227 : AOI211_X1 port map( C1 => DATA1(9), C2 => n4519, A => n3435, B => 
                           n3163, ZN => n3164);
   U228 : NAND2_X1 port map( A1 => n4074, A2 => n3619, ZN => n3372);
   U229 : NAND2_X1 port map( A1 => n3810, A2 => DATA1(6), ZN => n3513);
   U230 : NAND3_X1 port map( A1 => n3164, A2 => n3372, A3 => n3513, ZN => n3673
                           );
   U231 : INV_X1 port map( A => n3673, ZN => n3680);
   U232 : NOR2_X1 port map( A1 => n4242, A2 => n3471, ZN => n3401);
   U233 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(8), ZN => n3165);
   U234 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(6), ZN => n3473);
   U235 : NAND2_X1 port map( A1 => n3785, A2 => DATA1(5), ZN => n4011);
   U236 : INV_X1 port map( A => n3658, ZN => n3809);
   U237 : NAND2_X1 port map( A1 => n5136, A2 => n3809, ZN => n4521);
   U238 : NAND4_X1 port map( A1 => n3165, A2 => n3473, A3 => n4011, A4 => n4521
                           , ZN => n3166);
   U239 : NOR2_X1 port map( A1 => n3401, A2 => n3166, ZN => n3679);
   U240 : OAI222_X1 port map( A1 => n3871, A2 => n3680, B1 => n3768, B2 => 
                           n3679, C1 => n3168, C2 => n3900, ZN => n3715);
   U241 : AOI22_X1 port map( A1 => n4196, A2 => n3965, B1 => n4193, B2 => n3715
                           , ZN => n3176);
   U242 : INV_X1 port map( A => n4193, ZN => n4534);
   U243 : INV_X1 port map( A => n4534, ZN => n4161);
   U244 : OR2_X1 port map( A1 => n3167, A2 => n4161, ZN => n4535);
   U245 : INV_X1 port map( A => n4535, ZN => n4147);
   U246 : OAI222_X1 port map( A1 => n3871, A2 => n3679, B1 => n3768, B2 => 
                           n3168, C1 => n3173, C2 => n3852, ZN => n3963);
   U247 : OAI21_X1 port map( B1 => n4829, B2 => n4828, A => n4555, ZN => n3199)
                           ;
   U248 : AOI21_X1 port map( B1 => DATA2(1), B2 => DATA2(3), A => n3199, ZN => 
                           n3792);
   U249 : INV_X1 port map( A => n3792, ZN => n4542);
   U250 : OR3_X1 port map( A1 => n4542, A2 => n3169, A3 => n3510, ZN => n4537);
   U251 : INV_X1 port map( A => n4537, ZN => n3403);
   U252 : NOR2_X1 port map( A1 => n4007, A2 => n4008, ZN => n3172);
   U253 : INV_X1 port map( A => DATA1(0), ZN => n4750);
   U254 : NAND2_X1 port map( A1 => n4074, A2 => n5135, ZN => n4012);
   U255 : NAND2_X1 port map( A1 => n4519, A2 => n5136, ZN => n3170);
   U256 : OAI211_X1 port map( C1 => n3658, C2 => n4750, A => n4012, B => n3170,
                           ZN => n3171);
   U257 : AOI211_X1 port map( C1 => DATA1(1), C2 => n3785, A => n3172, B => 
                           n3171, ZN => n3466);
   U258 : OAI222_X1 port map( A1 => n3871, A2 => n3173, B1 => n3768, B2 => 
                           n3455, C1 => n3466, C2 => n3900, ZN => n3964);
   U259 : AOI22_X1 port map( A1 => n3837, A2 => n3963, B1 => n3403, B2 => n3964
                           , ZN => n3175);
   U260 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(4), ZN => n3344);
   U261 : NOR2_X1 port map( A1 => n4828, A2 => n3344, ZN => n3950);
   U262 : NAND2_X1 port map( A1 => n3950, A2 => DATA2(1), ZN => n4597);
   U263 : INV_X1 port map( A => n4597, ZN => n4288);
   U264 : OR2_X1 port map( A1 => n3174, A2 => DATA2(5), ZN => n3960);
   U265 : AOI211_X1 port map( C1 => DATA2(0), C2 => n4288, A => n4724, B => 
                           n3960, ZN => n3179);
   U266 : NAND2_X1 port map( A1 => n3179, A2 => n4796, ZN => n4467);
   U267 : AOI21_X1 port map( B1 => n3176, B2 => n3175, A => n4467, ZN => n3177)
                           ;
   U268 : AOI211_X1 port map( C1 => dataout_mul_9_port, C2 => n4491, A => n3178
                           , B => n3177, ZN => n3326);
   U269 : NAND2_X1 port map( A1 => FUNC(3), A2 => n3179, ZN => n4794);
   U270 : INV_X1 port map( A => n4794, ZN => n4506);
   U271 : INV_X1 port map( A => n3344, ZN => n3289);
   U272 : NOR2_X1 port map( A1 => n4555, A2 => n4828, ZN => n4279);
   U273 : INV_X1 port map( A => n4279, ZN => n4583);
   U274 : NAND4_X1 port map( A1 => DATA2(1), A2 => n3289, A3 => n4831, A4 => 
                           n4583, ZN => n4199);
   U275 : OAI221_X1 port map( B1 => n4829, B2 => n4555, C1 => n4830, C2 => 
                           n4555, A => n4583, ZN => n3272);
   U276 : NAND2_X1 port map( A1 => DATA2(4), A2 => n3454, ZN => n3286);
   U277 : NAND2_X1 port map( A1 => n3344, A2 => n4583, ZN => n4276);
   U278 : INV_X1 port map( A => n4276, ZN => n4572);
   U279 : NAND3_X1 port map( A1 => n3272, A2 => n3286, A3 => n4572, ZN => n4455
                           );
   U280 : INV_X1 port map( A => n4455, ZN => n4564);
   U281 : INV_X1 port map( A => DATA1(19), ZN => n4315);
   U282 : NOR2_X1 port map( A1 => n4242, A2 => n4315, ZN => n3571);
   U283 : INV_X1 port map( A => DATA1(22), ZN => n4202);
   U284 : NAND2_X1 port map( A1 => n4519, A2 => DATA1(18), ZN => n3568);
   U285 : NAND2_X1 port map( A1 => DATA1(20), A2 => n4520, ZN => n3649);
   U286 : OAI211_X1 port map( C1 => n4255, C2 => n4202, A => n3568, B => n3649,
                           ZN => n3180);
   U287 : AOI211_X1 port map( C1 => DATA1(21), C2 => n3810, A => n3571, B => 
                           n3180, ZN => n3196);
   U288 : INV_X1 port map( A => DATA1(18), ZN => n4324);
   U289 : NOR2_X1 port map( A1 => n4242, A2 => n4324, ZN => n3576);
   U290 : INV_X1 port map( A => DATA1(21), ZN => n4218);
   U291 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(17), ZN => n3582);
   U292 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(19), ZN => n3634);
   U293 : OAI211_X1 port map( C1 => n4255, C2 => n4218, A => n3582, B => n3634,
                           ZN => n3181);
   U294 : AOI211_X1 port map( C1 => DATA1(20), C2 => n3810, A => n3576, B => 
                           n3181, ZN => n3201);
   U295 : INV_X1 port map( A => DATA1(20), ZN => n4240);
   U296 : NOR2_X1 port map( A1 => n4242, A2 => n4240, ZN => n3633);
   U297 : INV_X1 port map( A => DATA1(23), ZN => n4163);
   U298 : NAND2_X1 port map( A1 => n4519, A2 => DATA1(19), ZN => n3578);
   U299 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(21), ZN => n3728);
   U300 : OAI211_X1 port map( C1 => n4255, C2 => n4163, A => n3578, B => n3728,
                           ZN => n3182);
   U301 : AOI211_X1 port map( C1 => DATA1(22), C2 => n3810, A => n3633, B => 
                           n3182, ZN => n3185);
   U302 : OAI222_X1 port map( A1 => n4115, A2 => n3196, B1 => n4113, B2 => 
                           n3201, C1 => n3185, C2 => n3900, ZN => n3233);
   U303 : NOR2_X1 port map( A1 => n4202, A2 => n4007, ZN => n3750);
   U304 : INV_X1 port map( A => DATA1(24), ZN => n4636);
   U305 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(21), ZN => n3646);
   U306 : NAND2_X1 port map( A1 => DATA1(20), A2 => n4519, ZN => n3572);
   U307 : OAI211_X1 port map( C1 => n4255, C2 => n4636, A => n3646, B => n3572,
                           ZN => n3183);
   U308 : AOI211_X1 port map( C1 => DATA1(23), C2 => n3785, A => n3750, B => 
                           n3183, ZN => n3189);
   U309 : OAI222_X1 port map( A1 => n3768, A2 => n3185, B1 => n3871, B2 => 
                           n3196, C1 => n3189, C2 => n3900, ZN => n3223);
   U310 : INV_X1 port map( A => n3223, ZN => n3204);
   U311 : AOI22_X1 port map( A1 => n3810, A2 => DATA1(24), B1 => DATA1(21), B2 
                           => n4519, ZN => n3184);
   U312 : NAND2_X1 port map( A1 => DATA1(22), A2 => n4074, ZN => n3727);
   U313 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(23), ZN => n3766);
   U314 : NAND2_X1 port map( A1 => DATA1(25), A2 => n3809, ZN => n3850);
   U315 : AND4_X1 port map( A1 => n3184, A2 => n3727, A3 => n3766, A4 => n3850,
                           ZN => n3188);
   U316 : OAI222_X1 port map( A1 => n3188, A2 => n3852, B1 => n3185, B2 => 
                           n4113, C1 => n3189, C2 => n4115, ZN => n3208);
   U317 : INV_X1 port map( A => n3208, ZN => n3215);
   U318 : OAI22_X1 port map( A1 => n3204, A2 => n4535, B1 => n3215, B2 => n4531
                           , ZN => n3191);
   U319 : CLKBUF_X1 port map( A => n3792, Z => n4263);
   U320 : AOI22_X1 port map( A1 => DATA1(23), A2 => n4258, B1 => DATA1(27), B2 
                           => n3809, ZN => n3186);
   U321 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(25), ZN => n3812);
   U322 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(24), ZN => n3765);
   U323 : NAND2_X1 port map( A1 => n3810, A2 => DATA1(26), ZN => n3849);
   U324 : AND4_X1 port map( A1 => n3186, A2 => n3812, A3 => n3765, A4 => n3849,
                           ZN => n3212);
   U325 : AOI22_X1 port map( A1 => n3785, A2 => DATA1(25), B1 => DATA1(22), B2 
                           => n4258, ZN => n3187);
   U326 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(23), ZN => n3746);
   U327 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(24), ZN => n3788);
   U328 : NAND2_X1 port map( A1 => DATA1(26), A2 => n4009, ZN => n3866);
   U329 : AND4_X1 port map( A1 => n3187, A2 => n3746, A3 => n3788, A4 => n3866,
                           ZN => n3207);
   U330 : OAI222_X1 port map( A1 => n3212, A2 => n3852, B1 => n3188, B2 => 
                           n4113, C1 => n3207, C2 => n3768, ZN => n3245);
   U331 : INV_X1 port map( A => n3245, ZN => n3214);
   U332 : OAI222_X1 port map( A1 => n3207, A2 => n3852, B1 => n3189, B2 => 
                           n4113, C1 => n3188, C2 => n3768, ZN => n3239);
   U333 : INV_X1 port map( A => n3239, ZN => n3213);
   U334 : OAI22_X1 port map( A1 => n4263, A2 => n3214, B1 => n3213, B2 => n4537
                           , ZN => n3190);
   U335 : AOI211_X1 port map( C1 => n3233, C2 => n4161, A => n3191, B => n3190,
                           ZN => n3249);
   U336 : NOR2_X1 port map( A1 => n4828, A2 => n3192, ZN => n3228);
   U337 : INV_X1 port map( A => n3228, ZN => n3205);
   U338 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(1), ZN => n3193);
   U339 : OAI21_X1 port map( B1 => n4829, B2 => n3193, A => n4555, ZN => n4020)
                           ;
   U340 : CLKBUF_X1 port map( A => n4020, Z => n3969);
   U341 : INV_X1 port map( A => n3969, ZN => n4550);
   U342 : NAND3_X1 port map( A1 => n3205, A2 => n4550, A3 => n3199, ZN => n4545
                           );
   U343 : NAND3_X1 port map( A1 => DATA2(3), A2 => n3454, A3 => n3194, ZN => 
                           n4547);
   U344 : INV_X1 port map( A => n4547, ZN => n4441);
   U345 : AOI22_X1 port map( A1 => DATA1(16), A2 => n4258, B1 => DATA1(20), B2 
                           => n4009, ZN => n3195);
   U346 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(18), ZN => n3573);
   U347 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(17), ZN => n3567);
   U348 : NAND2_X1 port map( A1 => n3810, A2 => DATA1(19), ZN => n3648);
   U349 : AND4_X1 port map( A1 => n3195, A2 => n3573, A3 => n3567, A4 => n3648,
                           ZN => n3221);
   U350 : OAI222_X1 port map( A1 => n3871, A2 => n3221, B1 => n4115, B2 => 
                           n3201, C1 => n3196, C2 => n3900, ZN => n3222);
   U351 : INV_X1 port map( A => n3222, ZN => n3263);
   U352 : OAI22_X1 port map( A1 => n4534, A2 => n3263, B1 => n3204, B2 => n4531
                           , ZN => n3198);
   U353 : OAI22_X1 port map( A1 => n3792, A2 => n3213, B1 => n3215, B2 => n4537
                           , ZN => n3197);
   U354 : AOI211_X1 port map( C1 => n4147, C2 => n3233, A => n3198, B => n3197,
                           ZN => n3265);
   U355 : INV_X1 port map( A => n3265, ZN => n3254);
   U356 : AOI21_X1 port map( B1 => n3454, B2 => DATA2(3), A => n3199, ZN => 
                           n4426);
   U357 : INV_X1 port map( A => n4426, ZN => n4543);
   U358 : INV_X1 port map( A => n4543, ZN => n4508);
   U359 : AOI22_X1 port map( A1 => DATA1(18), A2 => n3810, B1 => DATA1(19), B2 
                           => n4009, ZN => n3200);
   U360 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(16), ZN => n3581);
   U361 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(17), ZN => n3577);
   U362 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(15), ZN => n3591);
   U363 : AND4_X1 port map( A1 => n3200, A2 => n3581, A3 => n3577, A4 => n3591,
                           ZN => n3230);
   U364 : OAI222_X1 port map( A1 => n3871, A2 => n3230, B1 => n3768, B2 => 
                           n3221, C1 => n3201, C2 => n3900, ZN => n3260);
   U365 : AOI22_X1 port map( A1 => n4161, A2 => n3260, B1 => n3222, B2 => n4147
                           , ZN => n3203);
   U366 : AOI22_X1 port map( A1 => n3233, A2 => n4160, B1 => n4542, B2 => n3208
                           , ZN => n3202);
   U367 : OAI211_X1 port map( C1 => n4537, C2 => n3204, A => n3203, B => n3202,
                           ZN => n3234);
   U368 : AOI22_X1 port map( A1 => n4441, A2 => n3254, B1 => n4508, B2 => n3234
                           , ZN => n3219);
   U369 : NOR2_X1 port map( A1 => n4020, A2 => n3205, ZN => n4022);
   U370 : CLKBUF_X1 port map( A => n4542, Z => n4018);
   U371 : NOR2_X1 port map( A1 => n4248, A2 => n4636, ZN => n3749);
   U372 : INV_X1 port map( A => DATA1(25), ZN => n4708);
   U373 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(26), ZN => n3833);
   U374 : NAND2_X1 port map( A1 => n3785, A2 => DATA1(27), ZN => n3867);
   U375 : OAI211_X1 port map( C1 => n4708, C2 => n4242, A => n3833, B => n3867,
                           ZN => n3206);
   U376 : AOI211_X1 port map( C1 => DATA1(28), C2 => n4009, A => n3749, B => 
                           n3206, ZN => n3238);
   U377 : OAI222_X1 port map( A1 => n3871, A2 => n3207, B1 => n3768, B2 => 
                           n3212, C1 => n3238, C2 => n3852, ZN => n4192);
   U378 : AOI22_X1 port map( A1 => n3837, A2 => n3208, B1 => n4018, B2 => n4192
                           , ZN => n3210);
   U379 : AOI22_X1 port map( A1 => n3403, A2 => n3245, B1 => n4161, B2 => n3223
                           , ZN => n3209);
   U380 : OAI211_X1 port map( C1 => n3213, C2 => n4531, A => n3210, B => n3209,
                           ZN => n4318);
   U381 : AOI22_X1 port map( A1 => DATA1(28), A2 => n3785, B1 => DATA1(29), B2 
                           => n4009, ZN => n3211);
   U382 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(27), ZN => n3848);
   U383 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(26), ZN => n3811);
   U384 : NAND2_X1 port map( A1 => n4519, A2 => DATA1(25), ZN => n3764);
   U385 : AND4_X1 port map( A1 => n3211, A2 => n3848, A3 => n3811, A4 => n3764,
                           ZN => n3244);
   U386 : OAI222_X1 port map( A1 => n3244, A2 => n3900, B1 => n3212, B2 => 
                           n4113, C1 => n3238, C2 => n3768, ZN => n4194);
   U387 : INV_X1 port map( A => n4194, ZN => n3242);
   U388 : OAI22_X1 port map( A1 => n3792, A2 => n3242, B1 => n3213, B2 => n4535
                           , ZN => n3217);
   U389 : OAI22_X1 port map( A1 => n4534, A2 => n3215, B1 => n3214, B2 => n4531
                           , ZN => n3216);
   U390 : AOI211_X1 port map( C1 => n3403, C2 => n4192, A => n3217, B => n3216,
                           ZN => n3257);
   U391 : INV_X1 port map( A => n3257, ZN => n4319);
   U392 : AOI22_X1 port map( A1 => n4022, A2 => n4318, B1 => n3969, B2 => n4319
                           , ZN => n3218);
   U393 : OAI211_X1 port map( C1 => n3249, C2 => n4545, A => n3219, B => n3218,
                           ZN => n3285);
   U394 : INV_X1 port map( A => n3234, ZN => n3279);
   U395 : OAI22_X1 port map( A1 => n3265, A2 => n4545, B1 => n3279, B2 => n4547
                           , ZN => n3227);
   U396 : INV_X1 port map( A => n3260, ZN => n3278);
   U397 : INV_X1 port map( A => DATA1(15), ZN => n4621);
   U398 : NOR2_X1 port map( A1 => n4242, A2 => n4621, ZN => n3588);
   U399 : INV_X1 port map( A => DATA1(14), ZN => n4405);
   U400 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(16), ZN => n3566);
   U401 : NAND2_X1 port map( A1 => DATA1(18), A2 => n3809, ZN => n3647);
   U402 : OAI211_X1 port map( C1 => n4248, C2 => n4405, A => n3566, B => n3647,
                           ZN => n3220);
   U403 : AOI211_X1 port map( C1 => DATA1(17), C2 => n3785, A => n3588, B => 
                           n3220, ZN => n3259);
   U404 : OAI222_X1 port map( A1 => n3221, A2 => n3852, B1 => n3259, B2 => 
                           n4113, C1 => n3230, C2 => n4115, ZN => n3275);
   U405 : AOI22_X1 port map( A1 => n4160, A2 => n3222, B1 => n4161, B2 => n3275
                           , ZN => n3225);
   U406 : AOI22_X1 port map( A1 => n3403, A2 => n3233, B1 => n4018, B2 => n3223
                           , ZN => n3224);
   U407 : OAI211_X1 port map( C1 => n3278, C2 => n4535, A => n3225, B => n3224,
                           ZN => n3296);
   U408 : INV_X1 port map( A => n3296, ZN => n3264);
   U409 : INV_X1 port map( A => n4022, ZN => n4429);
   U410 : OAI22_X1 port map( A1 => n3264, A2 => n4543, B1 => n3249, B2 => n4429
                           , ZN => n3226);
   U411 : AOI211_X1 port map( C1 => n4020, C2 => n4318, A => n3227, B => n3226,
                           ZN => n3270);
   U412 : INV_X1 port map( A => n3270, ZN => n3284);
   U413 : AOI21_X1 port map( B1 => DATA2(1), B2 => n3228, A => n4028, ZN => 
                           n4026);
   U414 : CLKBUF_X1 port map( A => n4026, Z => n4407);
   U415 : NOR2_X1 port map( A1 => n4407, A2 => n4028, ZN => n4357);
   U416 : INV_X1 port map( A => n4545, ZN => n4440);
   U417 : AOI22_X1 port map( A1 => DATA1(16), A2 => n3810, B1 => DATA1(17), B2 
                           => n3809, ZN => n3229);
   U418 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(14), ZN => n3590);
   U419 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(15), ZN => n3580);
   U420 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(13), ZN => n3614);
   U421 : AND4_X1 port map( A1 => n3229, A2 => n3590, A3 => n3580, A4 => n3614,
                           ZN => n3274);
   U422 : OAI222_X1 port map( A1 => n3230, A2 => n3900, B1 => n3274, B2 => 
                           n4113, C1 => n3259, C2 => n3768, ZN => n3292);
   U423 : INV_X1 port map( A => n3292, ZN => n3307);
   U424 : OAI22_X1 port map( A1 => n4534, A2 => n3307, B1 => n3278, B2 => n4531
                           , ZN => n3232);
   U425 : INV_X1 port map( A => n3275, ZN => n3295);
   U426 : OAI22_X1 port map( A1 => n3295, A2 => n4535, B1 => n3263, B2 => n4537
                           , ZN => n3231);
   U427 : AOI211_X1 port map( C1 => n4018, C2 => n3233, A => n3232, B => n3231,
                           ZN => n3308);
   U428 : INV_X1 port map( A => n3308, ZN => n3268);
   U429 : AOI22_X1 port map( A1 => n4440, A2 => n3234, B1 => n4508, B2 => n3268
                           , ZN => n3236);
   U430 : CLKBUF_X1 port map( A => n4441, Z => n4425);
   U431 : CLKBUF_X1 port map( A => n4022, Z => n4554);
   U432 : AOI22_X1 port map( A1 => n4425, A2 => n3296, B1 => n4554, B2 => n3254
                           , ZN => n3235);
   U433 : OAI211_X1 port map( C1 => n4550, C2 => n3249, A => n3236, B => n3235,
                           ZN => n3269);
   U434 : AOI222_X1 port map( A1 => n3285, A2 => n4028, B1 => n3284, B2 => 
                           n4357, C1 => n3269, C2 => n4407, ZN => n4462);
   U435 : INV_X1 port map( A => n4462, ZN => n3312);
   U436 : INV_X1 port map( A => DATA1(28), ZN => n4642);
   U437 : NOR2_X1 port map( A1 => n4007, A2 => n4642, ZN => n3869);
   U438 : INV_X1 port map( A => DATA1(30), ZN => n4721);
   U439 : NAND2_X1 port map( A1 => n4519, A2 => DATA1(26), ZN => n3786);
   U440 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(27), ZN => n3832);
   U441 : OAI211_X1 port map( C1 => n3658, C2 => n4721, A => n3786, B => n3832,
                           ZN => n3237);
   U442 : AOI211_X1 port map( C1 => DATA1(29), C2 => n3785, A => n3869, B => 
                           n3237, ZN => n4112);
   U443 : OAI222_X1 port map( A1 => n3871, A2 => n3238, B1 => n4115, B2 => 
                           n3244, C1 => n4112, C2 => n3852, ZN => n4195);
   U444 : AOI22_X1 port map( A1 => n4160, A2 => n4192, B1 => n4542, B2 => n4195
                           , ZN => n3241);
   U445 : AOI22_X1 port map( A1 => n3837, A2 => n3245, B1 => n4161, B2 => n3239
                           , ZN => n3240);
   U446 : OAI211_X1 port map( C1 => n3242, C2 => n4537, A => n3241, B => n3240,
                           ZN => n4321);
   U447 : INV_X1 port map( A => n4321, ZN => n3252);
   U448 : INV_X1 port map( A => n4192, ZN => n3248);
   U449 : INV_X1 port map( A => DATA1(27), ZN => n4097);
   U450 : NOR2_X1 port map( A1 => n4248, A2 => n4097, ZN => n3816);
   U451 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(29), ZN => n3897);
   U452 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(28), ZN => n3847);
   U453 : OAI211_X1 port map( C1 => n4721, C2 => n4077, A => n3897, B => n3847,
                           ZN => n3243);
   U454 : AOI211_X1 port map( C1 => DATA1(31), C2 => n4009, A => n3816, B => 
                           n3243, ZN => n4114);
   U455 : OAI222_X1 port map( A1 => n3871, A2 => n3244, B1 => n3768, B2 => 
                           n4112, C1 => n4114, C2 => n3900, ZN => n4197);
   U456 : AOI22_X1 port map( A1 => n4160, A2 => n4194, B1 => n4018, B2 => n4197
                           , ZN => n3247);
   U457 : AOI22_X1 port map( A1 => n3403, A2 => n4195, B1 => n4161, B2 => n3245
                           , ZN => n3246);
   U458 : OAI211_X1 port map( C1 => n3248, C2 => n4535, A => n3247, B => n3246,
                           ZN => n4320);
   U459 : AOI22_X1 port map( A1 => n4440, A2 => n4319, B1 => n3969, B2 => n4320
                           , ZN => n3251);
   U460 : INV_X1 port map( A => n3249, ZN => n3253);
   U461 : AOI22_X1 port map( A1 => n4425, A2 => n4318, B1 => n4426, B2 => n3253
                           , ZN => n3250);
   U462 : OAI211_X1 port map( C1 => n3252, C2 => n4429, A => n3251, B => n3250,
                           ZN => n4356);
   U463 : AOI22_X1 port map( A1 => n4441, A2 => n3253, B1 => n3969, B2 => n4321
                           , ZN => n3256);
   U464 : AOI22_X1 port map( A1 => n4440, A2 => n4318, B1 => n4426, B2 => n3254
                           , ZN => n3255);
   U465 : OAI211_X1 port map( C1 => n3257, C2 => n4429, A => n3256, B => n3255,
                           ZN => n4358);
   U466 : CLKBUF_X1 port map( A => n4357, Z => n4370);
   U467 : AOI222_X1 port map( A1 => n4356, A2 => n4028, B1 => n4358, B2 => 
                           n4370, C1 => n3285, C2 => n4407, ZN => n4460);
   U468 : INV_X1 port map( A => n4407, ZN => n4558);
   U469 : AOI22_X1 port map( A1 => DATA1(15), A2 => n3785, B1 => DATA1(16), B2 
                           => n3809, ZN => n3258);
   U470 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(13), ZN => n3594);
   U471 : NAND2_X1 port map( A1 => n4520, A2 => n5138, ZN => n3585);
   U472 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(12), ZN => n3622);
   U473 : AND4_X1 port map( A1 => n3258, A2 => n3594, A3 => n3585, A4 => n3622,
                           ZN => n3291);
   U474 : OAI222_X1 port map( A1 => n3871, A2 => n3291, B1 => n3768, B2 => 
                           n3274, C1 => n3259, C2 => n3852, ZN => n3332);
   U475 : AOI22_X1 port map( A1 => n3275, A2 => n4160, B1 => n4161, B2 => n3332
                           , ZN => n3262);
   U476 : AOI22_X1 port map( A1 => n3292, A2 => n4147, B1 => n3260, B2 => n3403
                           , ZN => n3261);
   U477 : OAI211_X1 port map( C1 => n4263, C2 => n3263, A => n3262, B => n3261,
                           ZN => n3336);
   U478 : INV_X1 port map( A => n3336, ZN => n3280);
   U479 : OAI22_X1 port map( A1 => n3279, A2 => n4429, B1 => n3280, B2 => n4543
                           , ZN => n3267);
   U480 : OAI22_X1 port map( A1 => n4550, A2 => n3265, B1 => n3264, B2 => n4545
                           , ZN => n3266);
   U481 : AOI211_X1 port map( C1 => n4425, C2 => n3268, A => n3267, B => n3266,
                           ZN => n3300);
   U482 : INV_X1 port map( A => n4357, ZN => n4560);
   U483 : INV_X1 port map( A => n3269, ZN => n3283);
   U484 : OAI222_X1 port map( A1 => n4558, A2 => n3300, B1 => n4560, B2 => 
                           n3283, C1 => n3270, C2 => n4555, ZN => n3341);
   U485 : INV_X1 port map( A => n3341, ZN => n4458);
   U486 : OAI21_X1 port map( B1 => DATA2(3), B2 => DATA2(2), A => n4028, ZN => 
                           n3271);
   U487 : OAI21_X1 port map( B1 => n4555, B2 => n3510, A => n3271, ZN => n4457)
                           ;
   U488 : INV_X1 port map( A => n4457, ZN => n4562);
   U489 : NOR2_X1 port map( A1 => n3272, A2 => n4562, ZN => n4566);
   U490 : INV_X1 port map( A => n4566, ZN => n4461);
   U491 : OAI22_X1 port map( A1 => n4572, A2 => n4460, B1 => n4458, B2 => n4461
                           , ZN => n3288);
   U492 : AOI22_X1 port map( A1 => DATA1(14), A2 => n3785, B1 => DATA1(15), B2 
                           => n3809, ZN => n3273);
   U493 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(12), ZN => n3613);
   U494 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(13), ZN => n3589);
   U495 : NAND2_X1 port map( A1 => n4519, A2 => DATA1(11), ZN => n3610);
   U496 : AND4_X1 port map( A1 => n3273, A2 => n3613, A3 => n3589, A4 => n3610,
                           ZN => n3304);
   U497 : OAI222_X1 port map( A1 => n3274, A2 => n3852, B1 => n3304, B2 => 
                           n4113, C1 => n3291, C2 => n3768, ZN => n3376);
   U498 : AOI22_X1 port map( A1 => n3275, A2 => n3403, B1 => n4161, B2 => n3376
                           , ZN => n3277);
   U499 : CLKBUF_X1 port map( A => n4147, Z => n3837);
   U500 : AOI22_X1 port map( A1 => n3292, A2 => n4196, B1 => n3332, B2 => n3837
                           , ZN => n3276);
   U501 : OAI211_X1 port map( C1 => n4263, C2 => n3278, A => n3277, B => n3276,
                           ZN => n3335);
   U502 : INV_X1 port map( A => n3335, ZN => n3382);
   U503 : OAI22_X1 port map( A1 => n4550, A2 => n3279, B1 => n3382, B2 => n4543
                           , ZN => n3282);
   U504 : OAI22_X1 port map( A1 => n3308, A2 => n4545, B1 => n3280, B2 => n4547
                           , ZN => n3281);
   U505 : AOI211_X1 port map( C1 => n4554, C2 => n3296, A => n3282, B => n3281,
                           ZN => n3311);
   U506 : OAI222_X1 port map( A1 => n3283, A2 => n4555, B1 => n3300, B2 => 
                           n4560, C1 => n3311, C2 => n4558, ZN => n3340);
   U507 : INV_X1 port map( A => n3340, ZN => n3387);
   U508 : CLKBUF_X1 port map( A => n4457, Z => n4419);
   U509 : AOI222_X1 port map( A1 => n4358, A2 => n4028, B1 => n3285, B2 => 
                           n4357, C1 => n3284, C2 => n4407, ZN => n4456);
   U510 : NOR2_X1 port map( A1 => n4276, A2 => n3286, ZN => n3826);
   U511 : INV_X1 port map( A => n3826, ZN => n4459);
   U512 : OAI22_X1 port map( A1 => n3387, A2 => n4419, B1 => n4456, B2 => n4459
                           , ZN => n3287);
   U513 : AOI211_X1 port map( C1 => n4564, C2 => n3312, A => n3288, B => n3287,
                           ZN => n4493);
   U514 : NAND3_X1 port map( A1 => n4828, A2 => n3289, A3 => n3949, ZN => n4492
                           );
   U515 : INV_X1 port map( A => DATA1(11), ZN => n4473);
   U516 : NOR2_X1 port map( A1 => n4242, A2 => n4473, ZN => n3618);
   U517 : NAND2_X1 port map( A1 => n3785, A2 => DATA1(13), ZN => n3586);
   U518 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(12), ZN => n3595);
   U519 : OAI211_X1 port map( C1 => n4255, C2 => n4405, A => n3586, B => n3595,
                           ZN => n3290);
   U520 : AOI211_X1 port map( C1 => n4519, C2 => DATA1(10), A => n3618, B => 
                           n3290, ZN => n3331);
   U521 : OAI222_X1 port map( A1 => n3291, A2 => n3900, B1 => n3331, B2 => 
                           n4113, C1 => n3304, C2 => n3768, ZN => n3404);
   U522 : AOI22_X1 port map( A1 => n4147, A2 => n3376, B1 => n4161, B2 => n3404
                           , ZN => n3294);
   U523 : AOI22_X1 port map( A1 => n3403, A2 => n3292, B1 => n4196, B2 => n3332
                           , ZN => n3293);
   U524 : OAI211_X1 port map( C1 => n3792, C2 => n3295, A => n3294, B => n3293,
                           ZN => n3407);
   U525 : AOI22_X1 port map( A1 => n4440, A2 => n3336, B1 => n4508, B2 => n3407
                           , ZN => n3298);
   U526 : AOI22_X1 port map( A1 => n4441, A2 => n3335, B1 => n4020, B2 => n3296
                           , ZN => n3297);
   U527 : OAI211_X1 port map( C1 => n3308, C2 => n4429, A => n3298, B => n3297,
                           ZN => n3299);
   U528 : INV_X1 port map( A => n3299, ZN => n3339);
   U529 : OAI222_X1 port map( A1 => n4560, A2 => n3311, B1 => n4558, B2 => 
                           n3339, C1 => n3300, C2 => n4555, ZN => n3413);
   U530 : OAI22_X1 port map( A1 => n3387, A2 => n4461, B1 => n4458, B2 => n4455
                           , ZN => n3302);
   U531 : OAI22_X1 port map( A1 => n4572, A2 => n4456, B1 => n4462, B2 => n4459
                           , ZN => n3301);
   U532 : AOI211_X1 port map( C1 => n4562, C2 => n3413, A => n3302, B => n3301,
                           ZN => n4494);
   U533 : INV_X1 port map( A => n3413, ZN => n3388);
   U534 : INV_X1 port map( A => n3407, ZN => n3381);
   U535 : INV_X1 port map( A => DATA1(10), ZN => n4681);
   U536 : NOR2_X1 port map( A1 => n4242, A2 => n4681, ZN => n3607);
   U537 : INV_X1 port map( A => DATA1(13), ZN => n4423);
   U538 : NAND2_X1 port map( A1 => n3810, A2 => DATA1(12), ZN => n3593);
   U539 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(11), ZN => n3615);
   U540 : OAI211_X1 port map( C1 => n4255, C2 => n4423, A => n3593, B => n3615,
                           ZN => n3303);
   U541 : AOI211_X1 port map( C1 => n4258, C2 => DATA1(9), A => n3607, B => 
                           n3303, ZN => n3374);
   U542 : OAI222_X1 port map( A1 => n3304, A2 => n3852, B1 => n3374, B2 => 
                           n3871, C1 => n3331, C2 => n4115, ZN => n3437);
   U543 : AOI22_X1 port map( A1 => n3837, A2 => n3404, B1 => n4161, B2 => n3437
                           , ZN => n3306);
   U544 : AOI22_X1 port map( A1 => n3403, A2 => n3332, B1 => n4160, B2 => n3376
                           , ZN => n3305);
   U545 : OAI211_X1 port map( C1 => n4263, C2 => n3307, A => n3306, B => n3305,
                           ZN => n3441);
   U546 : INV_X1 port map( A => n3441, ZN => n3380);
   U547 : OAI22_X1 port map( A1 => n3381, A2 => n4547, B1 => n3380, B2 => n4543
                           , ZN => n3310);
   U548 : OAI22_X1 port map( A1 => n3308, A2 => n4550, B1 => n3382, B2 => n4545
                           , ZN => n3309);
   U549 : AOI211_X1 port map( C1 => n4022, C2 => n3336, A => n3310, B => n3309,
                           ZN => n3385);
   U550 : OAI222_X1 port map( A1 => n3311, A2 => n4555, B1 => n3339, B2 => 
                           n4560, C1 => n3385, C2 => n4558, ZN => n3329);
   U551 : AOI22_X1 port map( A1 => n4564, A2 => n3340, B1 => n4562, B2 => n3329
                           , ZN => n3314);
   U552 : CLKBUF_X1 port map( A => n3826, Z => n4568);
   U553 : AOI22_X1 port map( A1 => n4568, A2 => n3341, B1 => n4276, B2 => n3312
                           , ZN => n3313);
   U554 : OAI211_X1 port map( C1 => n3388, C2 => n4461, A => n3314, B => n3313,
                           ZN => n3450);
   U555 : INV_X1 port map( A => n3450, ZN => n3328);
   U556 : AOI21_X1 port map( B1 => n3510, B2 => n4583, A => n4572, ZN => n4472)
                           ;
   U557 : CLKBUF_X1 port map( A => n4472, Z => n4495);
   U558 : OAI222_X1 port map( A1 => n4199, A2 => n4493, B1 => n4492, B2 => 
                           n4494, C1 => n3328, C2 => n4495, ZN => n3324);
   U559 : NOR2_X1 port map( A1 => n3619, A2 => DATA2_I_8_port, ZN => n3327);
   U560 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n4374)
                           ;
   U561 : OAI21_X1 port map( B1 => DATA1(9), B2 => DATA2_I_9_port, A => n4374, 
                           ZN => n3542);
   U562 : NOR2_X1 port map( A1 => n3327, A2 => n3542, ZN => n4375);
   U563 : XNOR2_X1 port map( A => DATA2_I_7_port, B => n3471, ZN => n3397);
   U564 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n3362)
                           ;
   U565 : OAI21_X1 port map( B1 => DATA1(6), B2 => DATA2_I_6_port, A => n3362, 
                           ZN => n3425);
   U566 : NAND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n3361)
                           ;
   U567 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n3316)
                           ;
   U568 : INV_X1 port map( A => n3316, ZN => n3360);
   U569 : XOR2_X1 port map( A => DATA2_I_2_port, B => n4008, Z => n4049);
   U570 : INV_X1 port map( A => n4049, ZN => n4051);
   U571 : XOR2_X1 port map( A => DATA1(1), B => DATA2_I_1_port, Z => n4294);
   U572 : OAI21_X1 port map( B1 => n4780, B2 => DATA2_I_0_port, A => n4294, ZN 
                           => n4292);
   U573 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n4776)
                           ;
   U574 : INV_X1 port map( A => cin, ZN => n3356);
   U575 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n3357)
                           ;
   U576 : OAI221_X1 port map( B1 => n4292, B2 => n4776, C1 => n4292, C2 => 
                           n3356, A => n3357, ZN => n3315);
   U577 : AND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n3358);
   U578 : AOI21_X1 port map( B1 => n4051, B2 => n3315, A => n3358, ZN => n3317)
                           ;
   U579 : NAND2_X1 port map( A1 => n5135, A2 => DATA2_I_3_port, ZN => n3359);
   U580 : OAI21_X1 port map( B1 => DATA1(3), B2 => DATA2_I_3_port, A => n3359, 
                           ZN => n3540);
   U581 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n3316, 
                           ZN => n3355);
   U582 : AOI221_X1 port map( B1 => n3317, B2 => n3359, C1 => n3540, C2 => 
                           n3359, A => n3355, ZN => n3318);
   U583 : XOR2_X1 port map( A => DATA2_I_5_port, B => n4254, Z => n3463);
   U584 : INV_X1 port map( A => n3463, ZN => n3465);
   U585 : OAI21_X1 port map( B1 => n3360, B2 => n3318, A => n3465, ZN => n3319)
                           ;
   U586 : OAI221_X1 port map( B1 => n3425, B2 => n3361, C1 => n3425, C2 => 
                           n3319, A => n3362, ZN => n3320);
   U587 : AOI22_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, B1 => n3397,
                           B2 => n3320, ZN => n3547);
   U588 : INV_X1 port map( A => n3547, ZN => n4418);
   U589 : NAND2_X1 port map( A1 => n4797, A2 => n4418, ZN => n4496);
   U590 : AOI211_X1 port map( C1 => n3327, C2 => n3542, A => n4375, B => n4496,
                           ZN => n3323);
   U591 : NAND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n3321)
                           ;
   U592 : NOR2_X1 port map( A1 => n3542, A2 => n3321, ZN => n3545);
   U593 : NAND2_X1 port map( A1 => n4797, A2 => n3547, ZN => n4499);
   U594 : AOI211_X1 port map( C1 => n3542, C2 => n3321, A => n3545, B => n4499,
                           ZN => n3322);
   U595 : AOI211_X1 port map( C1 => n4506, C2 => n3324, A => n3323, B => n3322,
                           ZN => n3325);
   U596 : OAI211_X1 port map( C1 => n4768, C2 => n4479, A => n3326, B => n3325,
                           ZN => OUTALU(9));
   U597 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => DATA1(8), A => n3327, 
                           ZN => n3544);
   U598 : INV_X1 port map( A => n3544, ZN => n3354);
   U599 : OAI22_X1 port map( A1 => n3328, A2 => n4492, B1 => n4494, B2 => n4199
                           , ZN => n3352);
   U600 : INV_X1 port map( A => n3329, ZN => n3446);
   U601 : INV_X1 port map( A => n3437, ZN => n3375);
   U602 : NOR2_X1 port map( A1 => n4077, A2 => n4473, ZN => n3597);
   U603 : INV_X1 port map( A => DATA1(12), ZN => n4686);
   U604 : NAND2_X1 port map( A1 => n4073, A2 => DATA1(10), ZN => n3621);
   U605 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(9), ZN => n3662);
   U606 : OAI211_X1 port map( C1 => n3658, C2 => n4686, A => n3621, B => n3662,
                           ZN => n3330);
   U607 : AOI211_X1 port map( C1 => n4519, C2 => DATA1(8), A => n3597, B => 
                           n3330, ZN => n3402);
   U608 : OAI222_X1 port map( A1 => n3871, A2 => n3402, B1 => n4115, B2 => 
                           n3374, C1 => n3331, C2 => n3852, ZN => n3476);
   U609 : AOI22_X1 port map( A1 => n4196, A2 => n3404, B1 => n4161, B2 => n3476
                           , ZN => n3334);
   U610 : AOI22_X1 port map( A1 => n3403, A2 => n3376, B1 => n4542, B2 => n3332
                           , ZN => n3333);
   U611 : OAI211_X1 port map( C1 => n3375, C2 => n4535, A => n3334, B => n3333,
                           ZN => n3480);
   U612 : AOI22_X1 port map( A1 => n3407, A2 => n4440, B1 => n3480, B2 => n4426
                           , ZN => n3338);
   U613 : AOI22_X1 port map( A1 => n4020, A2 => n3336, B1 => n3335, B2 => n4022
                           , ZN => n3337);
   U614 : OAI211_X1 port map( C1 => n4547, C2 => n3380, A => n3338, B => n3337,
                           ZN => n3410);
   U615 : INV_X1 port map( A => n3410, ZN => n3386);
   U616 : OAI222_X1 port map( A1 => n3339, A2 => n4555, B1 => n3385, B2 => 
                           n4560, C1 => n3386, C2 => n4558, ZN => n3449);
   U617 : AOI22_X1 port map( A1 => n4568, A2 => n3340, B1 => n4562, B2 => n3449
                           , ZN => n3343);
   U618 : AOI22_X1 port map( A1 => n4564, A2 => n3413, B1 => n4276, B2 => n3341
                           , ZN => n3342);
   U619 : OAI211_X1 port map( C1 => n3446, C2 => n4461, A => n3343, B => n3342,
                           ZN => n3490);
   U620 : INV_X1 port map( A => n3490, ZN => n3346);
   U621 : NOR2_X1 port map( A1 => DATA2(3), A2 => n3344, ZN => n3345);
   U622 : NAND2_X1 port map( A1 => n3454, A2 => n3345, ZN => n4169);
   U623 : OAI22_X1 port map( A1 => n4495, A2 => n3346, B1 => n4493, B2 => n4169
                           , ZN => n3351);
   U624 : AOI222_X1 port map( A1 => n3963, A2 => n4161, B1 => n3964, B2 => 
                           n4196, C1 => n3965, C2 => n4147, ZN => n3349);
   U625 : INV_X1 port map( A => DATA2(8), ZN => n4821);
   U626 : INV_X1 port map( A => n3619, ZN => n4655);
   U627 : AOI22_X1 port map( A1 => n3619, A2 => DATA2(8), B1 => n4821, B2 => 
                           n4655, ZN => n4756);
   U628 : AOI22_X1 port map( A1 => dataout_mul_8_port, A2 => n4491, B1 => n4778
                           , B2 => n4756, ZN => n3348);
   U629 : NAND3_X1 port map( A1 => DATA2(8), A2 => n3619, A3 => n4450, ZN => 
                           n3347);
   U630 : OAI211_X1 port map( C1 => n3349, C2 => n4467, A => n3348, B => n3347,
                           ZN => n3350);
   U631 : AOI221_X1 port map( B1 => n3352, B2 => n4506, C1 => n3351, C2 => 
                           n4506, A => n3350, ZN => n3353);
   U632 : OAI221_X1 port map( B1 => n3544, B2 => n4496, C1 => n3354, C2 => 
                           n4499, A => n3353, ZN => OUTALU(8));
   U633 : NAND2_X1 port map( A1 => n4797, A2 => n3356, ZN => n4785);
   U634 : INV_X1 port map( A => n4785, ZN => n4001);
   U635 : INV_X1 port map( A => n4294, ZN => n4245);
   U636 : OAI21_X1 port map( B1 => n4776, B2 => n4245, A => n3357, ZN => n4004)
                           ;
   U637 : AOI21_X1 port map( B1 => n4051, B2 => n4004, A => n3358, ZN => n3535)
                           ;
   U638 : OAI21_X1 port map( B1 => n3535, B2 => n3540, A => n3359, ZN => n3496)
                           ;
   U639 : INV_X1 port map( A => n3355, ZN => n3502);
   U640 : AOI21_X1 port map( B1 => n3496, B2 => n3502, A => n3360, ZN => n3432)
                           ;
   U641 : OAI21_X1 port map( B1 => n3432, B2 => n3463, A => n3361, ZN => n3417)
                           ;
   U642 : INV_X1 port map( A => n3417, ZN => n3419);
   U643 : OAI21_X1 port map( B1 => n3419, B2 => n3425, A => n3362, ZN => n3364)
                           ;
   U644 : NOR2_X1 port map( A1 => n5139, A2 => n3356, ZN => n4779);
   U645 : NAND2_X1 port map( A1 => n3357, A2 => n4292, ZN => n4002);
   U646 : AOI21_X1 port map( B1 => n4051, B2 => n4002, A => n3358, ZN => n3534)
                           ;
   U647 : OAI21_X1 port map( B1 => n3534, B2 => n3540, A => n3359, ZN => n3495)
                           ;
   U648 : AOI21_X1 port map( B1 => n3495, B2 => n3502, A => n3360, ZN => n3431)
                           ;
   U649 : OAI21_X1 port map( B1 => n3431, B2 => n3463, A => n3361, ZN => n3416)
                           ;
   U650 : INV_X1 port map( A => n3416, ZN => n3418);
   U651 : OAI21_X1 port map( B1 => n3418, B2 => n3425, A => n3362, ZN => n3363)
                           ;
   U652 : AOI22_X1 port map( A1 => n4001, A2 => n3364, B1 => n4779, B2 => n3363
                           , ZN => n3396);
   U653 : INV_X1 port map( A => n4779, ZN => n4003);
   U654 : OAI22_X1 port map( A1 => n4785, A2 => n3364, B1 => n4003, B2 => n3363
                           , ZN => n3370);
   U655 : AOI22_X1 port map( A1 => n3837, A2 => n3964, B1 => n4161, B2 => n3965
                           , ZN => n3368);
   U656 : OAI21_X1 port map( B1 => n4471, B2 => n3471, A => n4470, ZN => n3365)
                           ;
   U657 : AOI22_X1 port map( A1 => DATA2(7), A2 => n3365, B1 => n4476, B2 => 
                           dataout_mul_7_port, ZN => n3367);
   U658 : NOR2_X1 port map( A1 => DATA2(7), A2 => n3471, ZN => n4656);
   U659 : INV_X1 port map( A => DATA2(7), ZN => n4824);
   U660 : NOR2_X1 port map( A1 => DATA1(7), A2 => n4824, ZN => n4672);
   U661 : OAI21_X1 port map( B1 => n4656, B2 => n4672, A => n4372, ZN => n3366)
                           ;
   U662 : OAI211_X1 port map( C1 => n3368, C2 => n4467, A => n3367, B => n3366,
                           ZN => n3369);
   U663 : AOI21_X1 port map( B1 => n3397, B2 => n3370, A => n3369, ZN => n3395)
                           ;
   U664 : NAND3_X1 port map( A1 => DATA2(4), A2 => DATA2(0), A3 => DATA2(3), ZN
                           => n3371);
   U665 : OAI211_X1 port map( C1 => DATA2(2), C2 => DATA2(1), A => DATA2(3), B 
                           => DATA2(4), ZN => n3981);
   U666 : NAND2_X1 port map( A1 => n3371, A2 => n3981, ZN => n4145);
   U667 : INV_X1 port map( A => n4145, ZN => n4585);
   U668 : INV_X1 port map( A => n4169, ZN => n4580);
   U669 : INV_X1 port map( A => n4494, ZN => n3391);
   U670 : AOI22_X1 port map( A1 => DATA1(7), A2 => n4258, B1 => DATA1(11), B2 
                           => n3809, ZN => n3373);
   U671 : NAND2_X1 port map( A1 => n3810, A2 => n5137, ZN => n3612);
   U672 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(9), ZN => n3609);
   U673 : AND4_X1 port map( A1 => n3373, A2 => n3612, A3 => n3609, A4 => n3372,
                           ZN => n3436);
   U674 : OAI222_X1 port map( A1 => n3374, A2 => n3900, B1 => n3436, B2 => 
                           n4113, C1 => n3402, C2 => n3768, ZN => n3477);
   U675 : INV_X1 port map( A => n3477, ZN => n3518);
   U676 : OAI22_X1 port map( A1 => n4534, A2 => n3518, B1 => n3375, B2 => n4531
                           , ZN => n3379);
   U677 : AOI22_X1 port map( A1 => n4542, A2 => n3376, B1 => n3404, B2 => n3403
                           , ZN => n3377);
   U678 : INV_X1 port map( A => n3377, ZN => n3378);
   U679 : AOI211_X1 port map( C1 => n3837, C2 => n3476, A => n3379, B => n3378,
                           ZN => n3521);
   U680 : OAI22_X1 port map( A1 => n3380, A2 => n4545, B1 => n3521, B2 => n4543
                           , ZN => n3384);
   U681 : OAI22_X1 port map( A1 => n4550, A2 => n3382, B1 => n3381, B2 => n4429
                           , ZN => n3383);
   U682 : AOI211_X1 port map( C1 => n4441, C2 => n3480, A => n3384, B => n3383,
                           ZN => n3398);
   U683 : OAI222_X1 port map( A1 => n4560, A2 => n3386, B1 => n4558, B2 => 
                           n3398, C1 => n3385, C2 => n4555, ZN => n3488);
   U684 : INV_X1 port map( A => n3488, ZN => n3526);
   U685 : OAI22_X1 port map( A1 => n3446, A2 => n4455, B1 => n3526, B2 => n4419
                           , ZN => n3390);
   U686 : OAI22_X1 port map( A1 => n3388, A2 => n4459, B1 => n4572, B2 => n3387
                           , ZN => n3389);
   U687 : AOI211_X1 port map( C1 => n4566, C2 => n3449, A => n3390, B => n3389,
                           ZN => n3493);
   U688 : INV_X1 port map( A => n3493, ZN => n3530);
   U689 : INV_X1 port map( A => n4472, ZN => n4574);
   U690 : AOI22_X1 port map( A1 => n4580, A2 => n3391, B1 => n3530, B2 => n4574
                           , ZN => n3393);
   U691 : INV_X1 port map( A => n4492, ZN => n4578);
   U692 : INV_X1 port map( A => n4199, ZN => n4576);
   U693 : AOI22_X1 port map( A1 => n4578, A2 => n3490, B1 => n4576, B2 => n3450
                           , ZN => n3392);
   U694 : OAI211_X1 port map( C1 => n4493, C2 => n4583, A => n3393, B => n3392,
                           ZN => n3453);
   U695 : NAND3_X1 port map( A1 => n4506, A2 => n4585, A3 => n3453, ZN => n3394
                           );
   U696 : OAI211_X1 port map( C1 => n3397, C2 => n3396, A => n3395, B => n3394,
                           ZN => OUTALU(7));
   U697 : INV_X1 port map( A => n3398, ZN => n3445);
   U698 : NAND2_X1 port map( A1 => n4520, A2 => DATA1(8), ZN => n3661);
   U699 : OAI211_X1 port map( C1 => n4255, C2 => n4681, A => n3399, B => n3661,
                           ZN => n3400);
   U700 : AOI211_X1 port map( C1 => DATA1(9), C2 => n3785, A => n3401, B => 
                           n3400, ZN => n3475);
   U701 : OAI222_X1 port map( A1 => n3871, A2 => n3475, B1 => n3768, B2 => 
                           n3436, C1 => n3402, C2 => n3900, ZN => n4017);
   U702 : AOI22_X1 port map( A1 => n4196, A2 => n3476, B1 => n4161, B2 => n4017
                           , ZN => n3406);
   U703 : AOI22_X1 port map( A1 => n3403, A2 => n3437, B1 => n4018, B2 => n3404
                           , ZN => n3405);
   U704 : OAI211_X1 port map( C1 => n3518, C2 => n4535, A => n3406, B => n3405,
                           ZN => n4019);
   U705 : AOI22_X1 port map( A1 => n4440, A2 => n3480, B1 => n4508, B2 => n4019
                           , ZN => n3409);
   U706 : AOI22_X1 port map( A1 => n4554, A2 => n3441, B1 => n3969, B2 => n3407
                           , ZN => n3408);
   U707 : OAI211_X1 port map( C1 => n3521, C2 => n4547, A => n3409, B => n3408,
                           ZN => n3484);
   U708 : AOI222_X1 port map( A1 => n4370, A2 => n3445, B1 => n4407, B2 => 
                           n3484, C1 => n3410, C2 => n4028, ZN => n4031);
   U709 : OAI22_X1 port map( A1 => n4031, A2 => n4457, B1 => n3526, B2 => n4461
                           , ZN => n3412);
   U710 : INV_X1 port map( A => n3449, ZN => n3485);
   U711 : OAI22_X1 port map( A1 => n3485, A2 => n4455, B1 => n3446, B2 => n4459
                           , ZN => n3411);
   U712 : AOI211_X1 port map( C1 => n4276, C2 => n3413, A => n3412, B => n3411,
                           ZN => n4035);
   U713 : INV_X1 port map( A => n4035, ZN => n3489);
   U714 : AOI22_X1 port map( A1 => n4578, A2 => n3530, B1 => n3489, B2 => n4574
                           , ZN => n3415);
   U715 : AOI22_X1 port map( A1 => n4580, A2 => n3450, B1 => n4576, B2 => n3490
                           , ZN => n3414);
   U716 : OAI211_X1 port map( C1 => n4494, C2 => n4583, A => n3415, B => n3414,
                           ZN => n3494);
   U717 : NAND2_X1 port map( A1 => n3981, A2 => n4145, ZN => n4131);
   U718 : INV_X1 port map( A => n4131, ZN => n4587);
   U719 : AOI22_X1 port map( A1 => n4585, A2 => n3494, B1 => n4587, B2 => n3453
                           , ZN => n3429);
   U720 : INV_X1 port map( A => n3425, ZN => n3427);
   U721 : OAI22_X1 port map( A1 => n4785, A2 => n3417, B1 => n4003, B2 => n3416
                           , ZN => n3426);
   U722 : OAI22_X1 port map( A1 => n3419, A2 => n4785, B1 => n3418, B2 => n4003
                           , ZN => n3424);
   U723 : INV_X1 port map( A => DATA2(6), ZN => n4825);
   U724 : INV_X1 port map( A => DATA1(6), ZN => n4604);
   U725 : AOI22_X1 port map( A1 => DATA1(6), A2 => n4825, B1 => DATA2(6), B2 =>
                           n4604, ZN => n4669);
   U726 : OAI21_X1 port map( B1 => n4471, B2 => n4604, A => n4470, ZN => n3420)
                           ;
   U727 : AOI22_X1 port map( A1 => DATA2(6), A2 => n3420, B1 => n4476, B2 => 
                           dataout_mul_6_port, ZN => n3422);
   U728 : INV_X1 port map( A => n4467, ZN => n4509);
   U729 : NAND3_X1 port map( A1 => n4509, A2 => n4161, A3 => n3964, ZN => n3421
                           );
   U730 : OAI211_X1 port map( C1 => n4669, C2 => n4479, A => n3422, B => n3421,
                           ZN => n3423);
   U731 : AOI221_X1 port map( B1 => n3427, B2 => n3426, C1 => n3425, C2 => 
                           n3424, A => n3423, ZN => n3428);
   U732 : OAI21_X1 port map( B1 => n3429, B2 => n4794, A => n3428, ZN => 
                           OUTALU(6));
   U733 : OAI22_X1 port map( A1 => n4785, A2 => n3432, B1 => n4003, B2 => n3431
                           , ZN => n3430);
   U734 : INV_X1 port map( A => n3430, ZN => n3464);
   U735 : AOI22_X1 port map( A1 => n4001, A2 => n3432, B1 => n4779, B2 => n3431
                           , ZN => n3462);
   U736 : OAI21_X1 port map( B1 => n4471, B2 => n4254, A => n4470, ZN => n3460)
                           ;
   U737 : INV_X1 port map( A => n3981, ZN => n4589);
   U738 : INV_X1 port map( A => n4019, ZN => n3444);
   U739 : INV_X1 port map( A => n3521, ZN => n3481);
   U740 : INV_X1 port map( A => n4017, ZN => n3440);
   U741 : NAND2_X1 port map( A1 => n3785, A2 => DATA1(8), ZN => n3608);
   U742 : OAI211_X1 port map( C1 => n3658, C2 => n3617, A => n3608, B => n3433,
                           ZN => n3434);
   U743 : AOI211_X1 port map( C1 => n4258, C2 => DATA1(5), A => n3435, B => 
                           n3434, ZN => n3511);
   U744 : OAI222_X1 port map( A1 => n3871, A2 => n3511, B1 => n4115, B2 => 
                           n3475, C1 => n3436, C2 => n3852, ZN => n3470);
   U745 : AOI22_X1 port map( A1 => n4160, A2 => n3477, B1 => n4161, B2 => n3470
                           , ZN => n3439);
   U746 : AOI22_X1 port map( A1 => n3403, A2 => n3476, B1 => n4542, B2 => n3437
                           , ZN => n3438);
   U747 : OAI211_X1 port map( C1 => n3440, C2 => n4535, A => n3439, B => n3438,
                           ZN => n4021);
   U748 : AOI22_X1 port map( A1 => n4440, A2 => n3481, B1 => n4508, B2 => n4021
                           , ZN => n3443);
   U749 : AOI22_X1 port map( A1 => n4022, A2 => n3480, B1 => n4020, B2 => n3441
                           , ZN => n3442);
   U750 : OAI211_X1 port map( C1 => n3444, C2 => n4547, A => n3443, B => n3442,
                           ZN => n3524);
   U751 : AOI222_X1 port map( A1 => n4357, A2 => n3484, B1 => n4026, B2 => 
                           n3524, C1 => n3445, C2 => n4028, ZN => n4030);
   U752 : OAI22_X1 port map( A1 => n3526, A2 => n4455, B1 => n4030, B2 => n4457
                           , ZN => n3448);
   U753 : OAI22_X1 port map( A1 => n4031, A2 => n4461, B1 => n4572, B2 => n3446
                           , ZN => n3447);
   U754 : AOI211_X1 port map( C1 => n3826, C2 => n3449, A => n3448, B => n3447,
                           ZN => n4034);
   U755 : INV_X1 port map( A => n4034, ZN => n4280);
   U756 : AOI22_X1 port map( A1 => n4578, A2 => n3489, B1 => n4574, B2 => n4280
                           , ZN => n3452);
   U757 : AOI22_X1 port map( A1 => n4580, A2 => n3490, B1 => n4279, B2 => n3450
                           , ZN => n3451);
   U758 : OAI211_X1 port map( C1 => n3493, C2 => n4199, A => n3452, B => n3451,
                           ZN => n3533);
   U759 : AOI222_X1 port map( A1 => n3453, A2 => n4589, B1 => n3494, B2 => 
                           n4587, C1 => n3533, C2 => n4585, ZN => n4250);
   U760 : OAI211_X1 port map( C1 => DATA2(2), C2 => n3454, A => DATA2(3), B => 
                           DATA2(4), ZN => n4126);
   U761 : INV_X1 port map( A => n4126, ZN => n4591);
   U762 : NOR3_X1 port map( A1 => n4250, A2 => n4794, A3 => n4591, ZN => n3459)
                           ;
   U763 : INV_X1 port map( A => DATA2(5), ZN => n4826);
   U764 : NAND2_X1 port map( A1 => DATA1(5), A2 => n4826, ZN => n4666);
   U765 : NAND2_X1 port map( A1 => DATA2(5), A2 => n4254, ZN => n4668);
   U766 : AND2_X1 port map( A1 => n4666, A2 => n4668, ZN => n4759);
   U767 : OAI22_X1 port map( A1 => n3455, A2 => n3871, B1 => n3466, B2 => n3768
                           , ZN => n3456);
   U768 : INV_X1 port map( A => n4403, ZN => n4789);
   U769 : AOI22_X1 port map( A1 => n4509, A2 => n3456, B1 => n4789, B2 => 
                           dataout_mul_5_port, ZN => n3457);
   U770 : OAI21_X1 port map( B1 => n4759, B2 => n4479, A => n3457, ZN => n3458)
                           ;
   U771 : AOI211_X1 port map( C1 => DATA2(5), C2 => n3460, A => n3459, B => 
                           n3458, ZN => n3461);
   U772 : OAI221_X1 port map( B1 => n3465, B2 => n3464, C1 => n3463, C2 => 
                           n3462, A => n3461, ZN => OUTALU(5));
   U773 : AOI22_X1 port map( A1 => n4001, A2 => n3496, B1 => n4779, B2 => n3495
                           , ZN => n3501);
   U774 : NOR3_X1 port map( A1 => n3466, A2 => n4467, A3 => n3871, ZN => n3469)
                           ;
   U775 : INV_X1 port map( A => DATA2(4), ZN => n4827);
   U776 : NOR2_X1 port map( A1 => n4827, A2 => n5136, ZN => n4663);
   U777 : INV_X1 port map( A => n4663, ZN => n4609);
   U778 : NAND2_X1 port map( A1 => n5136, A2 => n4827, ZN => n4667);
   U779 : AND2_X1 port map( A1 => n4609, A2 => n4667, ZN => n4767);
   U780 : INV_X1 port map( A => n4470, ZN => n4511);
   U781 : AOI21_X1 port map( B1 => n4510, B2 => DATA1(4), A => n4511, ZN => 
                           n3467);
   U782 : OAI22_X1 port map( A1 => n4767, A2 => n4479, B1 => n3467, B2 => n4827
                           , ZN => n3468);
   U783 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n4789, A => n3469
                           , B => n3468, ZN => n3500);
   U784 : INV_X1 port map( A => n4021, ZN => n4269);
   U785 : INV_X1 port map( A => n3470, ZN => n4262);
   U786 : NOR2_X1 port map( A1 => n4077, A2 => n3471, ZN => n3660);
   U787 : OAI211_X1 port map( C1 => n4255, C2 => n4655, A => n3473, B => n3472,
                           ZN => n3474);
   U788 : AOI211_X1 port map( C1 => n4258, C2 => DATA1(4), A => n3660, B => 
                           n3474, ZN => n3516);
   U789 : OAI222_X1 port map( A1 => n3871, A2 => n3516, B1 => n4115, B2 => 
                           n3511, C1 => n3475, C2 => n3900, ZN => n4541);
   U790 : AOI22_X1 port map( A1 => n4196, A2 => n4017, B1 => n4193, B2 => n4541
                           , ZN => n3479);
   U791 : AOI22_X1 port map( A1 => n3403, A2 => n3477, B1 => n4018, B2 => n3476
                           , ZN => n3478);
   U792 : OAI211_X1 port map( C1 => n4262, C2 => n4535, A => n3479, B => n3478,
                           ZN => n4023);
   U793 : AOI22_X1 port map( A1 => n4440, A2 => n4019, B1 => n4426, B2 => n4023
                           , ZN => n3483);
   U794 : AOI22_X1 port map( A1 => n4554, A2 => n3481, B1 => n3969, B2 => n3480
                           , ZN => n3482);
   U795 : OAI211_X1 port map( C1 => n4269, C2 => n4547, A => n3483, B => n3482,
                           ZN => n4029);
   U796 : AOI222_X1 port map( A1 => n3484, A2 => n4028, B1 => n3524, B2 => 
                           n4370, C1 => n4029, C2 => n4407, ZN => n4571);
   U797 : OAI22_X1 port map( A1 => n4031, A2 => n4455, B1 => n4571, B2 => n4419
                           , ZN => n3487);
   U798 : OAI22_X1 port map( A1 => n4572, A2 => n3485, B1 => n4030, B2 => n4461
                           , ZN => n3486);
   U799 : AOI211_X1 port map( C1 => n3826, C2 => n3488, A => n3487, B => n3486,
                           ZN => n4584);
   U800 : INV_X1 port map( A => n4584, ZN => n4281);
   U801 : AOI22_X1 port map( A1 => n4578, A2 => n4280, B1 => n4281, B2 => n4574
                           , ZN => n3492);
   U802 : AOI22_X1 port map( A1 => n4279, A2 => n3490, B1 => n4576, B2 => n3489
                           , ZN => n3491);
   U803 : OAI211_X1 port map( C1 => n3493, C2 => n4169, A => n3492, B => n3491,
                           ZN => n4039);
   U804 : AOI222_X1 port map( A1 => n3494, A2 => n4589, B1 => n3533, B2 => 
                           n4587, C1 => n4039, C2 => n4585, ZN => n4598);
   U805 : NOR2_X1 port map( A1 => n3950, A2 => n4126, ZN => n4602);
   U806 : INV_X1 port map( A => n4602, ZN => n4285);
   U807 : OAI22_X1 port map( A1 => n4598, A2 => n4591, B1 => n4250, B2 => n4285
                           , ZN => n3498);
   U808 : OAI22_X1 port map( A1 => n4785, A2 => n3496, B1 => n4003, B2 => n3495
                           , ZN => n3497);
   U809 : AOI22_X1 port map( A1 => n4506, A2 => n3498, B1 => n3502, B2 => n3497
                           , ZN => n3499);
   U810 : OAI211_X1 port map( C1 => n3502, C2 => n3501, A => n3500, B => n3499,
                           ZN => OUTALU(4));
   U811 : AOI22_X1 port map( A1 => n4001, A2 => n3535, B1 => n4779, B2 => n3534
                           , ZN => n3541);
   U812 : OAI211_X1 port map( C1 => n4510, C2 => n4511, A => n5135, B => 
                           DATA2(3), ZN => n3503);
   U813 : INV_X1 port map( A => n3503, ZN => n3509);
   U814 : NAND2_X1 port map( A1 => DATA1(3), A2 => n4828, ZN => n4664);
   U815 : INV_X1 port map( A => n4664, ZN => n3504);
   U816 : NOR2_X1 port map( A1 => DATA1(3), A2 => n4828, ZN => n4662);
   U817 : NOR2_X1 port map( A1 => n3504, A2 => n4662, ZN => n4761);
   U818 : NOR2_X1 port map( A1 => n4242, A2 => n4008, ZN => n4257);
   U819 : AOI22_X1 port map( A1 => n3810, A2 => DATA1(0), B1 => n4073, B2 => 
                           DATA1(1), ZN => n3505);
   U820 : INV_X1 port map( A => n3505, ZN => n3506);
   U821 : AOI211_X1 port map( C1 => n5135, C2 => n4258, A => n4257, B => n3506,
                           ZN => n3507);
   U822 : OAI22_X1 port map( A1 => n4761, A2 => n4479, B1 => n3507, B2 => n4467
                           , ZN => n3508);
   U823 : AOI211_X1 port map( C1 => dataout_mul_3_port, C2 => n4789, A => n3509
                           , B => n3508, ZN => n3539);
   U824 : NAND2_X1 port map( A1 => n3950, A2 => n3510, ZN => n4593);
   U825 : INV_X1 port map( A => n4030, ZN => n4275);
   U826 : INV_X1 port map( A => n4023, ZN => n4549);
   U827 : INV_X1 port map( A => n3511, ZN => n3517);
   U828 : AOI22_X1 port map( A1 => DATA1(3), A2 => n4519, B1 => DATA1(7), B2 =>
                           n3809, ZN => n3515);
   U829 : NAND4_X1 port map( A1 => n3515, A2 => n3514, A3 => n3513, A4 => n3512
                           , ZN => n4261);
   U830 : INV_X1 port map( A => n3516, ZN => n4014);
   U831 : AOI222_X1 port map( A1 => n3517, A2 => n4260, B1 => n4261, B2 => 
                           n4527, C1 => n4014, C2 => n4525, ZN => n4538);
   U832 : INV_X1 port map( A => n4541, ZN => n4264);
   U833 : OAI22_X1 port map( A1 => n4534, A2 => n4538, B1 => n4264, B2 => n4535
                           , ZN => n3520);
   U834 : OAI22_X1 port map( A1 => n3792, A2 => n3518, B1 => n4262, B2 => n4531
                           , ZN => n3519);
   U835 : AOI211_X1 port map( C1 => n3403, C2 => n4017, A => n3520, B => n3519,
                           ZN => n4268);
   U836 : OAI22_X1 port map( A1 => n4549, A2 => n4547, B1 => n4268, B2 => n4543
                           , ZN => n3523);
   U837 : OAI22_X1 port map( A1 => n4550, A2 => n3521, B1 => n4269, B2 => n4545
                           , ZN => n3522);
   U838 : AOI211_X1 port map( C1 => n4554, C2 => n4019, A => n3523, B => n3522,
                           ZN => n4273);
   U839 : INV_X1 port map( A => n4273, ZN => n4027);
   U840 : AOI222_X1 port map( A1 => n4370, A2 => n4029, B1 => n4026, B2 => 
                           n4027, C1 => n3524, C2 => n4028, ZN => n3525);
   U841 : INV_X1 port map( A => n3525, ZN => n4567);
   U842 : AOI22_X1 port map( A1 => n4564, A2 => n4275, B1 => n4562, B2 => n4567
                           , ZN => n3529);
   U843 : OAI22_X1 port map( A1 => n4459, A2 => n4031, B1 => n4572, B2 => n3526
                           , ZN => n3527);
   U844 : INV_X1 port map( A => n3527, ZN => n3528);
   U845 : OAI211_X1 port map( C1 => n4571, C2 => n4461, A => n3529, B => n3528,
                           ZN => n4579);
   U846 : AOI22_X1 port map( A1 => n4280, A2 => n4576, B1 => n4574, B2 => n4579
                           , ZN => n3532);
   U847 : AOI22_X1 port map( A1 => n4281, A2 => n4578, B1 => n3530, B2 => n4279
                           , ZN => n3531);
   U848 : OAI211_X1 port map( C1 => n4169, C2 => n4035, A => n3532, B => n3531,
                           ZN => n4284);
   U849 : AOI222_X1 port map( A1 => n3533, A2 => n4589, B1 => n4284, B2 => 
                           n4585, C1 => n4039, C2 => n4587, ZN => n4596);
   U850 : OAI222_X1 port map( A1 => n4285, A2 => n4598, B1 => n4593, B2 => 
                           n4250, C1 => n4591, C2 => n4596, ZN => n3537);
   U851 : OAI22_X1 port map( A1 => n3535, A2 => n4785, B1 => n3534, B2 => n4003
                           , ZN => n3536);
   U852 : AOI22_X1 port map( A1 => n4506, A2 => n3537, B1 => n3540, B2 => n3536
                           , ZN => n3538);
   U853 : OAI211_X1 port map( C1 => n3541, C2 => n3540, A => n3539, B => n3538,
                           ZN => OUTALU(3));
   U854 : INV_X1 port map( A => DATA1(31), ZN => n4723);
   U855 : OAI211_X1 port map( C1 => n4723, C2 => n4796, A => DATA2(31), B => 
                           n4372, ZN => n3988);
   U856 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n3557);
   U857 : AND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => n3996
                           );
   U858 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n3551);
   U859 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => n3551
                           , ZN => n4186);
   U860 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n4187);
   U861 : XOR2_X1 port map( A => DATA2_I_15_port, B => n4621, Z => n4391);
   U862 : INV_X1 port map( A => n4391, ZN => n4393);
   U863 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n4402);
   U864 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => n4402
                           , ZN => n4421);
   U865 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n4422);
   U866 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => n4422
                           , ZN => n4444);
   U867 : NOR2_X1 port map( A1 => n4421, A2 => n4444, ZN => n4381);
   U868 : NAND2_X1 port map( A1 => n5137, A2 => DATA2_I_10_port, ZN => n4373);
   U869 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => n4373
                           , ZN => n4501);
   U870 : NAND2_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, ZN => 
                           n4382);
   U871 : OAI21_X1 port map( B1 => DATA1(14), B2 => DATA2_I_14_port, A => n4382
                           , ZN => n4415);
   U872 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n4378);
   U873 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => n4378
                           , ZN => n4486);
   U874 : NOR4_X1 port map( A1 => n3542, A2 => n4501, A3 => n4415, A4 => n4486,
                           ZN => n3543);
   U875 : NAND3_X1 port map( A1 => n4381, A2 => n3544, A3 => n3543, ZN => n3546
                           );
   U876 : INV_X1 port map( A => n4415, ZN => n4417);
   U877 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => n4379
                           );
   U878 : AOI21_X1 port map( B1 => DATA2_I_9_port, B2 => DATA1(9), A => n3545, 
                           ZN => n4502);
   U879 : NOR2_X1 port map( A1 => n4502, A2 => n4501, ZN => n4500);
   U880 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => n5137, A => n4500, ZN
                           => n4487);
   U881 : OAI21_X1 port map( B1 => n4379, B2 => n4487, A => n4378, ZN => n4443)
                           ;
   U882 : NOR2_X1 port map( A1 => n4422, A2 => n4421, ZN => n4380);
   U883 : AOI21_X1 port map( B1 => n4381, B2 => n4443, A => n4380, ZN => n4400)
                           ;
   U884 : NAND2_X1 port map( A1 => n4400, A2 => n4402, ZN => n4397);
   U885 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n4417, B2 => n4397, ZN => n4390);
   U886 : OAI21_X1 port map( B1 => n3547, B2 => n3546, A => n4390, ZN => n3548)
                           ;
   U887 : AOI22_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, B1 => 
                           n4393, B2 => n3548, ZN => n4180);
   U888 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n4178);
   U889 : OAI21_X1 port map( B1 => DATA1(21), B2 => DATA2_I_21_port, A => n4178
                           , ZN => n4224);
   U890 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n4176);
   U891 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => n4176
                           , ZN => n4235);
   U892 : INV_X1 port map( A => DATA1(17), ZN => n4342);
   U893 : XOR2_X1 port map( A => DATA2_I_17_port, B => n4342, Z => n4350);
   U894 : INV_X1 port map( A => n4350, ZN => n4352);
   U895 : XOR2_X1 port map( A => DATA2_I_18_port, B => n4324, Z => n4333);
   U896 : INV_X1 port map( A => n4333, ZN => n4336);
   U897 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => n4349
                           );
   U898 : AOI21_X1 port map( B1 => DATA2_I_16_port, B2 => DATA1(16), A => n4349
                           , ZN => n4365);
   U899 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => n4175
                           );
   U900 : AOI21_X1 port map( B1 => DATA2_I_19_port, B2 => DATA1(19), A => n4175
                           , ZN => n4312);
   U901 : NAND4_X1 port map( A1 => n4352, A2 => n4336, A3 => n4365, A4 => n4312
                           , ZN => n3549);
   U902 : NOR4_X1 port map( A1 => n4180, A2 => n4224, A3 => n4235, A4 => n3549,
                           ZN => n3550);
   U903 : INV_X1 port map( A => n4235, ZN => n4237);
   U904 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n4172);
   U905 : NAND3_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, A3 => 
                           n4352, ZN => n4343);
   U906 : NAND2_X1 port map( A1 => n4172, A2 => n4343, ZN => n4331);
   U907 : AOI22_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, B1 => 
                           n4336, B2 => n4331, ZN => n4303);
   U908 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n4174);
   U909 : OAI21_X1 port map( B1 => n4303, B2 => n4175, A => n4174, ZN => n4230)
                           ;
   U910 : AOI22_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, B1 => 
                           n4237, B2 => n4230, ZN => n4214);
   U911 : OAI21_X1 port map( B1 => n4214, B2 => n4224, A => n4178, ZN => n4182)
                           ;
   U912 : XNOR2_X1 port map( A => DATA2_I_22_port, B => n4202, ZN => n4201);
   U913 : OAI21_X1 port map( B1 => n3550, B2 => n4182, A => n4201, ZN => n3552)
                           ;
   U914 : OAI221_X1 port map( B1 => n4186, B2 => n4187, C1 => n4186, C2 => 
                           n3552, A => n3551, ZN => n3555);
   U915 : NOR2_X1 port map( A1 => n5139, A2 => n3555, ZN => n4150);
   U916 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n3554);
   U917 : INV_X1 port map( A => n3554, ZN => n4065);
   U918 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n4082);
   U919 : XNOR2_X1 port map( A => DATA2_I_27_port, B => n4097, ZN => n4107);
   U920 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n3556);
   U921 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n3553);
   U922 : INV_X1 port map( A => n3553, ZN => n4120);
   U923 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n4149);
   U924 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => n3553
                           , ZN => n4137);
   U925 : NOR2_X1 port map( A1 => n4149, A2 => n4137, ZN => n4134);
   U926 : INV_X1 port map( A => DATA1(26), ZN => n4712);
   U927 : XNOR2_X1 port map( A => DATA2_I_26_port, B => n4712, ZN => n4121);
   U928 : OAI21_X1 port map( B1 => n4120, B2 => n4134, A => n4121, ZN => n4123)
                           ;
   U929 : NAND2_X1 port map( A1 => n3556, A2 => n4123, ZN => n4106);
   U930 : NAND2_X1 port map( A1 => n4107, A2 => n4106, ZN => n4105);
   U931 : OAI21_X1 port map( B1 => DATA1(28), B2 => DATA2_I_28_port, A => n3554
                           , ZN => n4090);
   U932 : AOI21_X1 port map( B1 => n4082, B2 => n4105, A => n4090, ZN => n4078)
                           ;
   U933 : INV_X1 port map( A => DATA1(29), ZN => n4052);
   U934 : XNOR2_X1 port map( A => DATA2_I_29_port, B => n4052, ZN => n4069);
   U935 : OAI21_X1 port map( B1 => n4065, B2 => n4078, A => n4069, ZN => n3560)
                           ;
   U936 : NAND2_X1 port map( A1 => n3555, A2 => n4797, ZN => n4135);
   U937 : INV_X1 port map( A => n4135, ZN => n4156);
   U938 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => n4157
                           );
   U939 : NOR2_X1 port map( A1 => n4157, A2 => n4137, ZN => n4136);
   U940 : OAI21_X1 port map( B1 => n4120, B2 => n4136, A => n4121, ZN => n4122)
                           ;
   U941 : NAND2_X1 port map( A1 => n3556, A2 => n4122, ZN => n4104);
   U942 : NAND2_X1 port map( A1 => n4107, A2 => n4104, ZN => n4103);
   U943 : AOI21_X1 port map( B1 => n4082, B2 => n4103, A => n4090, ZN => n4079)
                           ;
   U944 : OAI21_X1 port map( B1 => n4065, B2 => n4079, A => n4069, ZN => n3559)
                           ;
   U945 : AOI22_X1 port map( A1 => n4150, A2 => n3560, B1 => n4156, B2 => n3559
                           , ZN => n4058);
   U946 : XNOR2_X1 port map( A => DATA2_I_30_port, B => n4721, ZN => n4000);
   U947 : OAI22_X1 port map( A1 => n3996, A2 => n4058, B1 => n4000, B2 => n5139
                           , ZN => n3995);
   U948 : NAND2_X1 port map( A1 => n3557, A2 => n3995, ZN => n3955);
   U949 : INV_X1 port map( A => DATA2(31), ZN => n4798);
   U950 : AOI22_X1 port map( A1 => DATA2(31), A2 => n4510, B1 => n4372, B2 => 
                           n4798, ZN => n3564);
   U951 : AOI22_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, B1 => 
                           n3996, B2 => n4000, ZN => n3558);
   U952 : INV_X1 port map( A => n3558, ZN => n3561);
   U953 : INV_X1 port map( A => n4150, ZN => n4133);
   U954 : OAI22_X1 port map( A1 => n4133, A2 => n3560, B1 => n4135, B2 => n3559
                           , ZN => n3989);
   U955 : AOI22_X1 port map( A1 => n3561, A2 => n4797, B1 => n3989, B2 => n4000
                           , ZN => n3957);
   U956 : INV_X1 port map( A => n3957, ZN => n3562);
   U957 : AOI22_X1 port map( A1 => n4519, A2 => n4506, B1 => DATA2_I_31_port, 
                           B2 => n3562, ZN => n3563);
   U958 : OAI211_X1 port map( C1 => DATA2_I_31_port, C2 => n3955, A => n3564, B
                           => n3563, ZN => n3565);
   U959 : AOI22_X1 port map( A1 => DATA1(31), A2 => n3565, B1 => n4789, B2 => 
                           dataout_mul_31_port, ZN => n3987);
   U960 : AOI22_X1 port map( A1 => DATA1(15), A2 => n3785, B1 => n5138, B2 => 
                           n3809, ZN => n3569);
   U961 : NAND4_X1 port map( A1 => n3569, A2 => n3568, A3 => n3567, A4 => n3566
                           , ZN => n3604);
   U962 : INV_X1 port map( A => DATA1(16), ZN => n4603);
   U963 : NOR2_X1 port map( A1 => n3658, A2 => n4603, ZN => n3570);
   U964 : AOI211_X1 port map( C1 => n3785, C2 => DATA1(17), A => n3571, B => 
                           n3570, ZN => n3574);
   U965 : NAND3_X1 port map( A1 => n3574, A2 => n3573, A3 => n3572, ZN => n3651
                           );
   U966 : NOR2_X1 port map( A1 => n3658, A2 => n4621, ZN => n3575);
   U967 : AOI211_X1 port map( C1 => n3810, C2 => DATA1(16), A => n3576, B => 
                           n3575, ZN => n3579);
   U968 : NAND3_X1 port map( A1 => n3579, A2 => n3578, A3 => n3577, ZN => n3636
                           );
   U969 : AOI222_X1 port map( A1 => n3604, A2 => n4529, B1 => n3651, B2 => 
                           n4527, C1 => n3636, C2 => n4525, ZN => n3755);
   U970 : NOR2_X1 port map( A1 => n3658, A2 => n4423, ZN => n3584);
   U971 : NAND3_X1 port map( A1 => n3582, A2 => n3581, A3 => n3580, ZN => n3583
                           );
   U972 : AOI211_X1 port map( C1 => n5138, C2 => n3810, A => n3584, B => n3583,
                           ZN => n3600);
   U973 : INV_X1 port map( A => n3600, ZN => n3603);
   U974 : AOI222_X1 port map( A1 => n4527, A2 => n3636, B1 => n4525, B2 => 
                           n3604, C1 => n3603, C2 => n4529, ZN => n3734);
   U975 : INV_X1 port map( A => n3734, ZN => n3598);
   U976 : OAI211_X1 port map( C1 => n3658, C2 => n4686, A => n3586, B => n3585,
                           ZN => n3587);
   U977 : AOI211_X1 port map( C1 => DATA1(16), C2 => n4258, A => n3588, B => 
                           n3587, ZN => n3601);
   U978 : AND3_X1 port map( A1 => n3591, A2 => n3590, A3 => n3589, ZN => n3592)
                           ;
   U979 : OAI211_X1 port map( C1 => n4473, C2 => n4255, A => n3593, B => n3592,
                           ZN => n3626);
   U980 : INV_X1 port map( A => n3626, ZN => n3599);
   U981 : OAI211_X1 port map( C1 => n4255, C2 => n4681, A => n3595, B => n3594,
                           ZN => n3596);
   U982 : AOI211_X1 port map( C1 => n5138, C2 => n4258, A => n3597, B => n3596,
                           ZN => n3624);
   U983 : OAI222_X1 port map( A1 => n4113, A2 => n3601, B1 => n4115, B2 => 
                           n3599, C1 => n3624, C2 => n3852, ZN => n3667);
   U984 : AOI22_X1 port map( A1 => n4147, A2 => n3598, B1 => n4542, B2 => n3667
                           , ZN => n3606);
   U985 : OAI222_X1 port map( A1 => n3871, A2 => n3600, B1 => n4115, B2 => 
                           n3601, C1 => n3599, C2 => n3900, ZN => n3639);
   U986 : INV_X1 port map( A => n3601, ZN => n3602);
   U987 : AOI222_X1 port map( A1 => n4527, A2 => n3604, B1 => n4525, B2 => 
                           n3603, C1 => n3602, C2 => n4260, ZN => n3640);
   U988 : INV_X1 port map( A => n3640, ZN => n3654);
   U989 : AOI22_X1 port map( A1 => n3403, A2 => n3639, B1 => n4196, B2 => n3654
                           , ZN => n3605);
   U990 : OAI211_X1 port map( C1 => n4534, C2 => n3755, A => n3606, B => n3605,
                           ZN => n3668);
   U991 : AOI21_X1 port map( B1 => DATA1(7), B2 => n4009, A => n3607, ZN => 
                           n3611);
   U992 : NAND4_X1 port map( A1 => n3611, A2 => n3610, A3 => n3609, A4 => n3608
                           , ZN => n3672);
   U993 : AND3_X1 port map( A1 => n3614, A2 => n3613, A3 => n3612, ZN => n3616)
                           ;
   U994 : OAI211_X1 port map( C1 => n3658, C2 => n3617, A => n3616, B => n3615,
                           ZN => n3627);
   U995 : AOI21_X1 port map( B1 => n3619, B2 => n4009, A => n3618, ZN => n3623)
                           ;
   U996 : NAND2_X1 port map( A1 => n3785, A2 => DATA1(9), ZN => n3620);
   U997 : NAND4_X1 port map( A1 => n3623, A2 => n3622, A3 => n3621, A4 => n3620
                           , ZN => n3664);
   U998 : AOI222_X1 port map( A1 => n3672, A2 => n4529, B1 => n3627, B2 => 
                           n4527, C1 => n3664, C2 => n4525, ZN => n3682);
   U999 : INV_X1 port map( A => n3624, ZN => n3625);
   U1000 : AOI222_X1 port map( A1 => n3664, A2 => n4529, B1 => n3625, B2 => 
                           n4527, C1 => n3627, C2 => n4525, ZN => n3671);
   U1001 : OAI22_X1 port map( A1 => n3792, A2 => n3682, B1 => n3671, B2 => 
                           n4537, ZN => n3629);
   U1002 : INV_X1 port map( A => n3639, ZN => n3641);
   U1003 : AOI222_X1 port map( A1 => n3627, A2 => n4529, B1 => n3626, B2 => 
                           n4527, C1 => n3625, C2 => n4525, ZN => n3674);
   U1004 : OAI22_X1 port map( A1 => n4534, A2 => n3641, B1 => n3674, B2 => 
                           n4531, ZN => n3628);
   U1005 : AOI211_X1 port map( C1 => n3837, C2 => n3667, A => n3629, B => n3628
                           , ZN => n3657);
   U1006 : OAI22_X1 port map( A1 => n3792, A2 => n3671, B1 => n3674, B2 => 
                           n4537, ZN => n3631);
   U1007 : OAI22_X1 port map( A1 => n4534, A2 => n3640, B1 => n3641, B2 => 
                           n4535, ZN => n3630);
   U1008 : AOI211_X1 port map( C1 => n4160, C2 => n3667, A => n3631, B => n3630
                           , ZN => n3698);
   U1009 : OAI22_X1 port map( A1 => n4550, A2 => n3657, B1 => n3698, B2 => 
                           n4429, ZN => n3645);
   U1010 : OAI22_X1 port map( A1 => n3734, A2 => n4531, B1 => n3640, B2 => 
                           n4537, ZN => n3638);
   U1011 : NOR2_X1 port map( A1 => n4255, A2 => n4342, ZN => n3632);
   U1012 : AOI211_X1 port map( C1 => n3810, C2 => DATA1(18), A => n3633, B => 
                           n3632, ZN => n3635);
   U1013 : OAI211_X1 port map( C1 => n4248, C2 => n4218, A => n3635, B => n3634
                           , ZN => n3732);
   U1014 : AOI222_X1 port map( A1 => n3636, A2 => n4260, B1 => n3732, B2 => 
                           n4527, C1 => n3651, C2 => n4525, ZN => n3771);
   U1015 : OAI22_X1 port map( A1 => n4534, A2 => n3771, B1 => n3755, B2 => 
                           n4535, ZN => n3637);
   U1016 : AOI211_X1 port map( C1 => n4018, C2 => n3639, A => n3638, B => n3637
                           , ZN => n3774);
   U1017 : OAI22_X1 port map( A1 => n4263, A2 => n3674, B1 => n4534, B2 => 
                           n3734, ZN => n3643);
   U1018 : OAI22_X1 port map( A1 => n3641, A2 => n4531, B1 => n3640, B2 => 
                           n4535, ZN => n3642);
   U1019 : AOI211_X1 port map( C1 => n3403, C2 => n3667, A => n3643, B => n3642
                           , ZN => n3737);
   U1020 : OAI22_X1 port map( A1 => n3774, A2 => n4543, B1 => n3737, B2 => 
                           n4545, ZN => n3644);
   U1021 : AOI211_X1 port map( C1 => n4425, C2 => n3668, A => n3645, B => n3644
                           , ZN => n3741);
   U1022 : OAI22_X1 port map( A1 => n4550, A2 => n3698, B1 => n3737, B2 => 
                           n4429, ZN => n3656);
   U1023 : AND4_X1 port map( A1 => n3649, A2 => n3648, A3 => n3647, A4 => n3646
                           , ZN => n3650);
   U1024 : OAI21_X1 port map( B1 => n4202, B2 => n4248, A => n3650, ZN => n3731
                           );
   U1025 : AOI222_X1 port map( A1 => n3651, A2 => n4260, B1 => n3731, B2 => 
                           n4527, C1 => n3732, C2 => n4525, ZN => n3791);
   U1026 : OAI22_X1 port map( A1 => n4534, A2 => n3791, B1 => n3771, B2 => 
                           n4535, ZN => n3653);
   U1027 : OAI22_X1 port map( A1 => n3755, A2 => n4531, B1 => n3734, B2 => 
                           n4537, ZN => n3652);
   U1028 : AOI211_X1 port map( C1 => n4542, C2 => n3654, A => n3653, B => n3652
                           , ZN => n3797);
   U1029 : OAI22_X1 port map( A1 => n3774, A2 => n4547, B1 => n3797, B2 => 
                           n4543, ZN => n3655);
   U1030 : AOI211_X1 port map( C1 => n4440, C2 => n3668, A => n3656, B => n3655
                           , ZN => n3759);
   U1031 : INV_X1 port map( A => n3657, ZN => n3702);
   U1032 : NOR2_X1 port map( A1 => n3658, A2 => n4604, ZN => n3659);
   U1033 : AOI211_X1 port map( C1 => n5137, C2 => n4519, A => n3660, B => n3659
                           , ZN => n3663);
   U1034 : NAND3_X1 port map( A1 => n3663, A2 => n3662, A3 => n3661, ZN => 
                           n3678);
   U1035 : AOI222_X1 port map( A1 => n3678, A2 => n4260, B1 => n3664, B2 => 
                           n4527, C1 => n3672, C2 => n4525, ZN => n3677);
   U1036 : OAI22_X1 port map( A1 => n4263, A2 => n3677, B1 => n3671, B2 => 
                           n4531, ZN => n3666);
   U1037 : OAI22_X1 port map( A1 => n3674, A2 => n4535, B1 => n3682, B2 => 
                           n4537, ZN => n3665);
   U1038 : AOI211_X1 port map( C1 => n4161, C2 => n3667, A => n3666, B => n3665
                           , ZN => n3692);
   U1039 : OAI22_X1 port map( A1 => n4550, A2 => n3692, B1 => n3698, B2 => 
                           n4545, ZN => n3670);
   U1040 : INV_X1 port map( A => n3668, ZN => n3756);
   U1041 : OAI22_X1 port map( A1 => n3756, A2 => n4543, B1 => n3737, B2 => 
                           n4547, ZN => n3669);
   U1042 : AOI211_X1 port map( C1 => n4022, C2 => n3702, A => n3670, B => n3669
                           , ZN => n3709);
   U1043 : OAI222_X1 port map( A1 => n4560, A2 => n3741, B1 => n4558, B2 => 
                           n3759, C1 => n3709, C2 => n4555, ZN => n3784);
   U1044 : INV_X1 port map( A => n3671, ZN => n3683);
   U1045 : AOI222_X1 port map( A1 => n3673, A2 => n4529, B1 => n3672, B2 => 
                           n4527, C1 => n3678, C2 => n4525, ZN => n3716);
   U1046 : OAI22_X1 port map( A1 => n4263, A2 => n3716, B1 => n3682, B2 => 
                           n4531, ZN => n3676);
   U1047 : OAI22_X1 port map( A1 => n4534, A2 => n3674, B1 => n3677, B2 => 
                           n4537, ZN => n3675);
   U1048 : AOI211_X1 port map( C1 => n4147, C2 => n3683, A => n3676, B => n3675
                           , ZN => n3701);
   U1049 : INV_X1 port map( A => n3677, ZN => n3688);
   U1050 : INV_X1 port map( A => n3678, ZN => n3681);
   U1051 : OAI222_X1 port map( A1 => n3871, A2 => n3681, B1 => n3768, B2 => 
                           n3680, C1 => n3679, C2 => n3852, ZN => n3962);
   U1052 : AOI22_X1 port map( A1 => n4160, A2 => n3688, B1 => n4018, B2 => 
                           n3962, ZN => n3685);
   U1053 : INV_X1 port map( A => n3682, ZN => n3689);
   U1054 : AOI22_X1 port map( A1 => n3837, A2 => n3689, B1 => n4193, B2 => 
                           n3683, ZN => n3684);
   U1055 : OAI211_X1 port map( C1 => n3716, C2 => n4537, A => n3685, B => n3684
                           , ZN => n3970);
   U1056 : AOI22_X1 port map( A1 => n4196, A2 => n3962, B1 => n4193, B2 => 
                           n3688, ZN => n3687);
   U1057 : AOI22_X1 port map( A1 => n3403, A2 => n3715, B1 => n4018, B2 => 
                           n3963, ZN => n3686);
   U1058 : OAI211_X1 port map( C1 => n3716, C2 => n4535, A => n3687, B => n3686
                           , ZN => n4439);
   U1059 : AOI22_X1 port map( A1 => n4440, A2 => n3970, B1 => n4020, B2 => 
                           n4439, ZN => n3694);
   U1060 : AOI22_X1 port map( A1 => n3837, A2 => n3688, B1 => n3403, B2 => 
                           n3962, ZN => n3691);
   U1061 : AOI22_X1 port map( A1 => n4018, A2 => n3715, B1 => n4193, B2 => 
                           n3689, ZN => n3690);
   U1062 : OAI211_X1 port map( C1 => n3716, C2 => n4531, A => n3691, B => n3690
                           , ZN => n4427);
   U1063 : INV_X1 port map( A => n3692, ZN => n3703);
   U1064 : AOI22_X1 port map( A1 => n4022, A2 => n4427, B1 => n4508, B2 => 
                           n3703, ZN => n3693);
   U1065 : OAI211_X1 port map( C1 => n3701, C2 => n4547, A => n3694, B => n3693
                           , ZN => n3973);
   U1066 : INV_X1 port map( A => n3970, ZN => n3697);
   U1067 : INV_X1 port map( A => n3701, ZN => n3719);
   U1068 : AOI22_X1 port map( A1 => n4440, A2 => n3719, B1 => n3969, B2 => 
                           n4427, ZN => n3696);
   U1069 : AOI22_X1 port map( A1 => n4441, A2 => n3703, B1 => n4508, B2 => 
                           n3702, ZN => n3695);
   U1070 : OAI211_X1 port map( C1 => n3697, C2 => n4429, A => n3696, B => n3695
                           , ZN => n3723);
   U1071 : AOI22_X1 port map( A1 => n4440, A2 => n3703, B1 => n4020, B2 => 
                           n3970, ZN => n3700);
   U1072 : INV_X1 port map( A => n3698, ZN => n3704);
   U1073 : AOI22_X1 port map( A1 => n4441, A2 => n3702, B1 => n4508, B2 => 
                           n3704, ZN => n3699);
   U1074 : OAI211_X1 port map( C1 => n3701, C2 => n4429, A => n3700, B => n3699
                           , ZN => n3708);
   U1075 : AOI222_X1 port map( A1 => n3973, A2 => n4028, B1 => n3723, B2 => 
                           n4357, C1 => n3708, C2 => n4407, ZN => n4304);
   U1076 : AOI22_X1 port map( A1 => n4440, A2 => n3702, B1 => n3969, B2 => 
                           n3719, ZN => n3706);
   U1077 : AOI22_X1 port map( A1 => n4425, A2 => n3704, B1 => n4022, B2 => 
                           n3703, ZN => n3705);
   U1078 : OAI211_X1 port map( C1 => n3737, C2 => n4543, A => n3706, B => n3705
                           , ZN => n3707);
   U1079 : AOI222_X1 port map( A1 => n3723, A2 => n4028, B1 => n3708, B2 => 
                           n4370, C1 => n3707, C2 => n4026, ZN => n3975);
   U1080 : OAI22_X1 port map( A1 => n4572, A2 => n4304, B1 => n3975, B2 => 
                           n4459, ZN => n3713);
   U1081 : INV_X1 port map( A => n3707, ZN => n3710);
   U1082 : OAI222_X1 port map( A1 => n3710, A2 => n4555, B1 => n3709, B2 => 
                           n4560, C1 => n3741, C2 => n4558, ZN => n3763);
   U1083 : INV_X1 port map( A => n3763, ZN => n3744);
   U1084 : INV_X1 port map( A => n3708, ZN => n3711);
   U1085 : OAI222_X1 port map( A1 => n3711, A2 => n4555, B1 => n3710, B2 => 
                           n4560, C1 => n3709, C2 => n4558, ZN => n3745);
   U1086 : INV_X1 port map( A => n3745, ZN => n3974);
   U1087 : OAI22_X1 port map( A1 => n3744, A2 => n4461, B1 => n3974, B2 => 
                           n4455, ZN => n3712);
   U1088 : AOI211_X1 port map( C1 => n4562, C2 => n3784, A => n3713, B => n3712
                           , ZN => n4198);
   U1089 : INV_X1 port map( A => n3975, ZN => n4305);
   U1090 : INV_X1 port map( A => n4439, ZN => n3722);
   U1091 : AOI22_X1 port map( A1 => n3962, A2 => n4147, B1 => n3963, B2 => 
                           n3403, ZN => n3714);
   U1092 : INV_X1 port map( A => n3714, ZN => n3718);
   U1093 : INV_X1 port map( A => n3715, ZN => n3968);
   U1094 : OAI22_X1 port map( A1 => n4534, A2 => n3716, B1 => n3968, B2 => 
                           n4531, ZN => n3717);
   U1095 : AOI211_X1 port map( C1 => n4542, C2 => n3965, A => n3718, B => n3717
                           , ZN => n4475);
   U1096 : INV_X1 port map( A => n4475, ZN => n4442);
   U1097 : AOI22_X1 port map( A1 => n3969, A2 => n4442, B1 => n4427, B2 => 
                           n4440, ZN => n3721);
   U1098 : AOI22_X1 port map( A1 => n3719, A2 => n4426, B1 => n3970, B2 => 
                           n4425, ZN => n3720);
   U1099 : OAI211_X1 port map( C1 => n4429, C2 => n3722, A => n3721, B => n3720
                           , ZN => n4371);
   U1100 : AOI222_X1 port map( A1 => n4357, A2 => n3973, B1 => n4026, B2 => 
                           n3723, C1 => n4371, C2 => n4028, ZN => n3724);
   U1101 : INV_X1 port map( A => n3724, ZN => n4341);
   U1102 : AOI22_X1 port map( A1 => n4564, A2 => n4305, B1 => n4276, B2 => 
                           n4341, ZN => n3726);
   U1103 : AOI22_X1 port map( A1 => n4562, A2 => n3763, B1 => n4566, B2 => 
                           n3745, ZN => n3725);
   U1104 : OAI211_X1 port map( C1 => n4304, C2 => n4459, A => n3726, B => n3725
                           , ZN => n4168);
   U1105 : AOI22_X1 port map( A1 => n3826, A2 => n3745, B1 => n4276, B2 => 
                           n4305, ZN => n3743);
   U1106 : INV_X1 port map( A => n3774, ZN => n3740);
   U1107 : NOR2_X1 port map( A1 => n4255, A2 => n4315, ZN => n3730);
   U1108 : OAI211_X1 port map( C1 => n4248, C2 => n4163, A => n3728, B => n3727
                           , ZN => n3729);
   U1109 : AOI211_X1 port map( C1 => DATA1(20), C2 => n3785, A => n3730, B => 
                           n3729, ZN => n3769);
   U1110 : INV_X1 port map( A => n3731, ZN => n3751);
   U1111 : INV_X1 port map( A => n3732, ZN => n3733);
   U1112 : OAI222_X1 port map( A1 => n4113, A2 => n3769, B1 => n4115, B2 => 
                           n3751, C1 => n3733, C2 => n3900, ZN => n3818);
   U1113 : OAI22_X1 port map( A1 => n3792, A2 => n3734, B1 => n3791, B2 => 
                           n4535, ZN => n3736);
   U1114 : OAI22_X1 port map( A1 => n3771, A2 => n4531, B1 => n3755, B2 => 
                           n4537, ZN => n3735);
   U1115 : AOI211_X1 port map( C1 => n4161, C2 => n3818, A => n3736, B => n3735
                           , ZN => n3823);
   U1116 : OAI22_X1 port map( A1 => n3823, A2 => n4543, B1 => n3756, B2 => 
                           n4429, ZN => n3739);
   U1117 : OAI22_X1 port map( A1 => n4550, A2 => n3737, B1 => n3797, B2 => 
                           n4547, ZN => n3738);
   U1118 : AOI211_X1 port map( C1 => n4440, C2 => n3740, A => n3739, B => n3738
                           , ZN => n3777);
   U1119 : OAI222_X1 port map( A1 => n4560, A2 => n3759, B1 => n4558, B2 => 
                           n3777, C1 => n3741, C2 => n4555, ZN => n3825);
   U1120 : AOI22_X1 port map( A1 => n4562, A2 => n3825, B1 => n4566, B2 => 
                           n3784, ZN => n3742);
   U1121 : OAI211_X1 port map( C1 => n3744, C2 => n4455, A => n3743, B => n3742
                           , ZN => n3806);
   U1122 : AOI22_X1 port map( A1 => n4279, A2 => n4168, B1 => n4576, B2 => 
                           n3806, ZN => n3782);
   U1123 : INV_X1 port map( A => n3825, ZN => n3762);
   U1124 : AOI22_X1 port map( A1 => n3826, A2 => n3763, B1 => n4276, B2 => 
                           n3745, ZN => n3761);
   U1125 : NAND2_X1 port map( A1 => DATA1(20), A2 => n3809, ZN => n3747);
   U1126 : OAI211_X1 port map( C1 => n4218, C2 => n4077, A => n3747, B => n3746
                           , ZN => n3748);
   U1127 : NOR3_X1 port map( A1 => n3750, A2 => n3749, A3 => n3748, ZN => n3790
                           );
   U1128 : OAI222_X1 port map( A1 => n4113, A2 => n3790, B1 => n4115, B2 => 
                           n3769, C1 => n3751, C2 => n3852, ZN => n3838);
   U1129 : AOI22_X1 port map( A1 => n3837, A2 => n3818, B1 => n4193, B2 => 
                           n3838, ZN => n3754);
   U1130 : OAI22_X1 port map( A1 => n4537, A2 => n3771, B1 => n4531, B2 => 
                           n3791, ZN => n3752);
   U1131 : INV_X1 port map( A => n3752, ZN => n3753);
   U1132 : OAI211_X1 port map( C1 => n4263, C2 => n3755, A => n3754, B => n3753
                           , ZN => n3841);
   U1133 : OAI22_X1 port map( A1 => n4550, A2 => n3756, B1 => n3797, B2 => 
                           n4545, ZN => n3758);
   U1134 : OAI22_X1 port map( A1 => n3774, A2 => n4429, B1 => n3823, B2 => 
                           n4547, ZN => n3757);
   U1135 : AOI211_X1 port map( C1 => n4426, C2 => n3841, A => n3758, B => n3757
                           , ZN => n3800);
   U1136 : OAI222_X1 port map( A1 => n4560, A2 => n3777, B1 => n4558, B2 => 
                           n3800, C1 => n3759, C2 => n4555, ZN => n3889);
   U1137 : AOI22_X1 port map( A1 => n4564, A2 => n3784, B1 => n4562, B2 => 
                           n3889, ZN => n3760);
   U1138 : OAI211_X1 port map( C1 => n3762, C2 => n4461, A => n3761, B => n3760
                           , ZN => n3939);
   U1139 : INV_X1 port map( A => n3889, ZN => n3780);
   U1140 : AOI22_X1 port map( A1 => n4568, A2 => n3784, B1 => n4276, B2 => 
                           n3763, ZN => n3779);
   U1141 : OAI22_X1 port map( A1 => n3823, A2 => n4545, B1 => n3797, B2 => 
                           n4429, ZN => n3776);
   U1142 : AOI22_X1 port map( A1 => DATA1(22), A2 => n3810, B1 => DATA1(21), B2
                           => n3809, ZN => n3767);
   U1143 : AND4_X1 port map( A1 => n3767, A2 => n3766, A3 => n3765, A4 => n3764
                           , ZN => n3817);
   U1144 : OAI222_X1 port map( A1 => n3769, A2 => n3852, B1 => n3817, B2 => 
                           n4113, C1 => n3790, C2 => n3768, ZN => n3854);
   U1145 : AOI22_X1 port map( A1 => n4161, A2 => n3854, B1 => n3838, B2 => 
                           n3837, ZN => n3770);
   U1146 : INV_X1 port map( A => n3770, ZN => n3773);
   U1147 : OAI22_X1 port map( A1 => n4263, A2 => n3771, B1 => n3791, B2 => 
                           n4537, ZN => n3772);
   U1148 : AOI211_X1 port map( C1 => n4160, C2 => n3818, A => n3773, B => n3772
                           , ZN => n3860);
   U1149 : OAI22_X1 port map( A1 => n4550, A2 => n3774, B1 => n3860, B2 => 
                           n4543, ZN => n3775);
   U1150 : AOI211_X1 port map( C1 => n4441, C2 => n3841, A => n3776, B => n3775
                           , ZN => n3807);
   U1151 : OAI222_X1 port map( A1 => n4560, A2 => n3800, B1 => n4558, B2 => 
                           n3807, C1 => n3777, C2 => n4555, ZN => n3862);
   U1152 : AOI22_X1 port map( A1 => n4564, A2 => n3825, B1 => n4562, B2 => 
                           n3862, ZN => n3778);
   U1153 : OAI211_X1 port map( C1 => n3780, C2 => n4461, A => n3779, B => n3778
                           , ZN => n3803);
   U1154 : AOI22_X1 port map( A1 => n4578, A2 => n3939, B1 => n4574, B2 => 
                           n3803, ZN => n3781);
   U1155 : OAI211_X1 port map( C1 => n4198, C2 => n4169, A => n3782, B => n3781
                           , ZN => n3783);
   U1156 : INV_X1 port map( A => n3783, ZN => n4132);
   U1157 : INV_X1 port map( A => n3862, ZN => n3885);
   U1158 : AOI22_X1 port map( A1 => n3826, A2 => n3825, B1 => n4276, B2 => 
                           n3784, ZN => n3802);
   U1159 : INV_X1 port map( A => n3860, ZN => n3842);
   U1160 : INV_X1 port map( A => n3841, ZN => n3796);
   U1161 : AOI22_X1 port map( A1 => DATA1(23), A2 => n3785, B1 => DATA1(22), B2
                           => n3809, ZN => n3789);
   U1162 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(25), ZN => n3787);
   U1163 : AND4_X1 port map( A1 => n3789, A2 => n3788, A3 => n3787, A4 => n3786
                           , ZN => n3836);
   U1164 : OAI222_X1 port map( A1 => n3790, A2 => n3900, B1 => n3836, B2 => 
                           n4113, C1 => n3817, C2 => n4115, ZN => n3872);
   U1165 : INV_X1 port map( A => n3872, ZN => n3857);
   U1166 : OAI22_X1 port map( A1 => n3792, A2 => n3791, B1 => n4534, B2 => 
                           n3857, ZN => n3795);
   U1167 : AOI22_X1 port map( A1 => n3818, A2 => n3403, B1 => n3854, B2 => 
                           n3837, ZN => n3793);
   U1168 : INV_X1 port map( A => n3793, ZN => n3794);
   U1169 : AOI211_X1 port map( C1 => n4196, C2 => n3838, A => n3795, B => n3794
                           , ZN => n3845);
   U1170 : OAI22_X1 port map( A1 => n3796, A2 => n4545, B1 => n3845, B2 => 
                           n4543, ZN => n3799);
   U1171 : OAI22_X1 port map( A1 => n4550, A2 => n3797, B1 => n3823, B2 => 
                           n4429, ZN => n3798);
   U1172 : AOI211_X1 port map( C1 => n4441, C2 => n3842, A => n3799, B => n3798
                           , ZN => n3808);
   U1173 : OAI222_X1 port map( A1 => n4560, A2 => n3807, B1 => n4558, B2 => 
                           n3808, C1 => n3800, C2 => n4555, ZN => n3881);
   U1174 : AOI22_X1 port map( A1 => n4564, A2 => n3889, B1 => n4562, B2 => 
                           n3881, ZN => n3801);
   U1175 : OAI211_X1 port map( C1 => n3885, C2 => n4461, A => n3802, B => n3801
                           , ZN => n3945);
   U1176 : INV_X1 port map( A => n3945, ZN => n3933);
   U1177 : OAI22_X1 port map( A1 => n4583, A2 => n4198, B1 => n4495, B2 => 
                           n3933, ZN => n3805);
   U1178 : INV_X1 port map( A => n3806, ZN => n4167);
   U1179 : INV_X1 port map( A => n3803, ZN => n3942);
   U1180 : OAI22_X1 port map( A1 => n4169, A2 => n4167, B1 => n4492, B2 => 
                           n3942, ZN => n3804);
   U1181 : AOI211_X1 port map( C1 => n3939, C2 => n4576, A => n3805, B => n3804
                           , ZN => n3982);
   U1182 : AOI22_X1 port map( A1 => n4580, A2 => n3939, B1 => n4279, B2 => 
                           n3806, ZN => n3830);
   U1183 : INV_X1 port map( A => n3807, ZN => n3824);
   U1184 : INV_X1 port map( A => n3808, ZN => n3846);
   U1185 : NAND2_X1 port map( A1 => DATA1(23), A2 => n3809, ZN => n3814);
   U1186 : NAND2_X1 port map( A1 => n3810, A2 => DATA1(24), ZN => n3813);
   U1187 : NAND4_X1 port map( A1 => n3814, A2 => n3813, A3 => n3812, A4 => 
                           n3811, ZN => n3815);
   U1188 : NOR2_X1 port map( A1 => n3816, A2 => n3815, ZN => n3853);
   U1189 : OAI222_X1 port map( A1 => n4113, A2 => n3853, B1 => n4115, B2 => 
                           n3836, C1 => n3817, C2 => n3900, ZN => n3906);
   U1190 : AOI22_X1 port map( A1 => n3403, A2 => n3838, B1 => n4193, B2 => 
                           n3906, ZN => n3820);
   U1191 : AOI22_X1 port map( A1 => n4196, A2 => n3854, B1 => n4542, B2 => 
                           n3818, ZN => n3819);
   U1192 : OAI211_X1 port map( C1 => n3857, C2 => n4535, A => n3820, B => n3819
                           , ZN => n3913);
   U1193 : AOI22_X1 port map( A1 => n4554, A2 => n3841, B1 => n4426, B2 => 
                           n3913, ZN => n3822);
   U1194 : INV_X1 port map( A => n3845, ZN => n3876);
   U1195 : AOI22_X1 port map( A1 => n4425, A2 => n3876, B1 => n4440, B2 => 
                           n3842, ZN => n3821);
   U1196 : OAI211_X1 port map( C1 => n4550, C2 => n3823, A => n3822, B => n3821
                           , ZN => n3861);
   U1197 : AOI222_X1 port map( A1 => n3824, A2 => n4028, B1 => n3846, B2 => 
                           n4357, C1 => n3861, C2 => n4026, ZN => n3924);
   U1198 : AOI22_X1 port map( A1 => n4564, A2 => n3862, B1 => n4276, B2 => 
                           n3825, ZN => n3828);
   U1199 : AOI22_X1 port map( A1 => n3826, A2 => n3889, B1 => n4566, B2 => 
                           n3881, ZN => n3827);
   U1200 : OAI211_X1 port map( C1 => n3924, C2 => n4419, A => n3828, B => n3827
                           , ZN => n3890);
   U1201 : AOI22_X1 port map( A1 => n4578, A2 => n3945, B1 => n4574, B2 => 
                           n3890, ZN => n3829);
   U1202 : OAI211_X1 port map( C1 => n3942, C2 => n4199, A => n3830, B => n3829
                           , ZN => n3831);
   U1203 : INV_X1 port map( A => n3831, ZN => n3952);
   U1204 : OAI222_X1 port map( A1 => n4132, A2 => n3981, B1 => n3982, B2 => 
                           n4131, C1 => n3952, C2 => n4145, ZN => n4071);
   U1205 : INV_X1 port map( A => n4071, ZN => n4096);
   U1206 : NOR2_X1 port map( A1 => n4077, A2 => n4708, ZN => n3835);
   U1207 : OAI211_X1 port map( C1 => n4248, C2 => n4642, A => n3833, B => n3832
                           , ZN => n3834);
   U1208 : AOI211_X1 port map( C1 => DATA1(24), C2 => n4009, A => n3835, B => 
                           n3834, ZN => n3870);
   U1209 : OAI222_X1 port map( A1 => n3871, A2 => n3870, B1 => n4115, B2 => 
                           n3853, C1 => n3836, C2 => n3852, ZN => n3896);
   U1210 : AOI22_X1 port map( A1 => n3837, A2 => n3906, B1 => n4193, B2 => 
                           n3896, ZN => n3840);
   U1211 : AOI22_X1 port map( A1 => n3403, A2 => n3854, B1 => n4542, B2 => 
                           n3838, ZN => n3839);
   U1212 : OAI211_X1 port map( C1 => n3857, C2 => n4531, A => n3840, B => n3839
                           , ZN => n3895);
   U1213 : AOI22_X1 port map( A1 => n4508, A2 => n3895, B1 => n4020, B2 => 
                           n3841, ZN => n3844);
   U1214 : AOI22_X1 port map( A1 => n4441, A2 => n3913, B1 => n4554, B2 => 
                           n3842, ZN => n3843);
   U1215 : OAI211_X1 port map( C1 => n3845, C2 => n4545, A => n3844, B => n3843
                           , ZN => n3880);
   U1216 : AOI222_X1 port map( A1 => n3846, A2 => n4028, B1 => n3861, B2 => 
                           n4370, C1 => n3880, C2 => n4026, ZN => n3923);
   U1217 : AOI22_X1 port map( A1 => n3913, A2 => n4440, B1 => n3895, B2 => 
                           n4425, ZN => n3859);
   U1218 : NAND4_X1 port map( A1 => n3850, A2 => n3849, A3 => n3848, A4 => 
                           n3847, ZN => n3851);
   U1219 : AOI21_X1 port map( B1 => n4519, B2 => DATA1(29), A => n3851, ZN => 
                           n3901);
   U1220 : OAI222_X1 port map( A1 => n3853, A2 => n3852, B1 => n3901, B2 => 
                           n4113, C1 => n3870, C2 => n3768, ZN => n3905);
   U1221 : AOI22_X1 port map( A1 => n4161, A2 => n3905, B1 => n3906, B2 => 
                           n4196, ZN => n3856);
   U1222 : AOI22_X1 port map( A1 => n4018, A2 => n3854, B1 => n3896, B2 => 
                           n4147, ZN => n3855);
   U1223 : OAI211_X1 port map( C1 => n4537, C2 => n3857, A => n3856, B => n3855
                           , ZN => n3912);
   U1224 : AOI22_X1 port map( A1 => n3876, A2 => n4554, B1 => n3912, B2 => 
                           n4508, ZN => n3858);
   U1225 : OAI211_X1 port map( C1 => n4550, C2 => n3860, A => n3859, B => n3858
                           , ZN => n3920);
   U1226 : AOI222_X1 port map( A1 => n4370, A2 => n3880, B1 => n4026, B2 => 
                           n3920, C1 => n3861, C2 => n4028, ZN => n3922);
   U1227 : INV_X1 port map( A => n3922, ZN => n3884);
   U1228 : AOI22_X1 port map( A1 => n4562, A2 => n3884, B1 => n4276, B2 => 
                           n3862, ZN => n3865);
   U1229 : INV_X1 port map( A => n3924, ZN => n3863);
   U1230 : AOI22_X1 port map( A1 => n4564, A2 => n3863, B1 => n4568, B2 => 
                           n3881, ZN => n3864);
   U1231 : OAI211_X1 port map( C1 => n3923, C2 => n4461, A => n3865, B => n3864
                           , ZN => n3928);
   U1232 : INV_X1 port map( A => n3912, ZN => n3879);
   U1233 : INV_X1 port map( A => n3906, ZN => n3875);
   U1234 : OAI211_X1 port map( C1 => n4248, C2 => n4721, A => n3867, B => n3866
                           , ZN => n3868);
   U1235 : AOI211_X1 port map( C1 => DATA1(29), C2 => n4074, A => n3869, B => 
                           n3868, ZN => n3902);
   U1236 : OAI222_X1 port map( A1 => n3871, A2 => n3902, B1 => n4115, B2 => 
                           n3901, C1 => n3870, C2 => n3900, ZN => n3907);
   U1237 : AOI22_X1 port map( A1 => n4196, A2 => n3896, B1 => n4193, B2 => 
                           n3907, ZN => n3874);
   U1238 : AOI22_X1 port map( A1 => n4147, A2 => n3905, B1 => n4018, B2 => 
                           n3872, ZN => n3873);
   U1239 : OAI211_X1 port map( C1 => n3875, C2 => n4537, A => n3874, B => n3873
                           , ZN => n3914);
   U1240 : AOI22_X1 port map( A1 => n4440, A2 => n3895, B1 => n4508, B2 => 
                           n3914, ZN => n3878);
   U1241 : AOI22_X1 port map( A1 => n4022, A2 => n3913, B1 => n3969, B2 => 
                           n3876, ZN => n3877);
   U1242 : OAI211_X1 port map( C1 => n3879, C2 => n4547, A => n3878, B => n3877
                           , ZN => n3919);
   U1243 : AOI222_X1 port map( A1 => n3880, A2 => n4028, B1 => n3920, B2 => 
                           n4357, C1 => n3919, C2 => n4026, ZN => n3894);
   U1244 : OAI22_X1 port map( A1 => n3923, A2 => n4455, B1 => n3894, B2 => 
                           n4457, ZN => n3883);
   U1245 : INV_X1 port map( A => n3881, ZN => n3886);
   U1246 : OAI22_X1 port map( A1 => n4572, A2 => n3886, B1 => n3924, B2 => 
                           n4459, ZN => n3882);
   U1247 : AOI211_X1 port map( C1 => n4566, C2 => n3884, A => n3883, B => n3882
                           , ZN => n3893);
   U1248 : OAI22_X1 port map( A1 => n3885, A2 => n4459, B1 => n3923, B2 => 
                           n4419, ZN => n3888);
   U1249 : OAI22_X1 port map( A1 => n3886, A2 => n4455, B1 => n3924, B2 => 
                           n4461, ZN => n3887);
   U1250 : AOI211_X1 port map( C1 => n4276, C2 => n3889, A => n3888, B => n3887
                           , ZN => n3940);
   U1251 : OAI22_X1 port map( A1 => n4472, A2 => n3893, B1 => n3940, B2 => 
                           n4199, ZN => n3892);
   U1252 : INV_X1 port map( A => n3890, ZN => n3941);
   U1253 : OAI22_X1 port map( A1 => n3933, A2 => n4583, B1 => n3941, B2 => 
                           n4169, ZN => n3891);
   U1254 : AOI211_X1 port map( C1 => n4578, C2 => n3928, A => n3892, B => n3891
                           , ZN => n3947);
   U1255 : INV_X1 port map( A => n3893, ZN => n3932);
   U1256 : INV_X1 port map( A => n3894, ZN => n3927);
   U1257 : INV_X1 port map( A => n3895, ZN => n3917);
   U1258 : INV_X1 port map( A => n3896, ZN => n3910);
   U1259 : NOR2_X1 port map( A1 => n4242, A2 => n4721, ZN => n4053);
   U1260 : NAND2_X1 port map( A1 => DATA1(27), A2 => n4009, ZN => n3898);
   U1261 : OAI211_X1 port map( C1 => n4077, C2 => n4642, A => n3898, B => n3897
                           , ZN => n3899);
   U1262 : AOI211_X1 port map( C1 => DATA1(31), C2 => n4519, A => n4053, B => 
                           n3899, ZN => n3903);
   U1263 : OAI222_X1 port map( A1 => n4113, A2 => n3903, B1 => n4115, B2 => 
                           n3902, C1 => n3901, C2 => n3900, ZN => n3904);
   U1264 : AOI22_X1 port map( A1 => n4160, A2 => n3905, B1 => n4193, B2 => 
                           n3904, ZN => n3909);
   U1265 : AOI22_X1 port map( A1 => n4147, A2 => n3907, B1 => n4018, B2 => 
                           n3906, ZN => n3908);
   U1266 : OAI211_X1 port map( C1 => n3910, C2 => n4537, A => n3909, B => n3908
                           , ZN => n3911);
   U1267 : AOI22_X1 port map( A1 => n4440, A2 => n3912, B1 => n4426, B2 => 
                           n3911, ZN => n3916);
   U1268 : AOI22_X1 port map( A1 => n4425, A2 => n3914, B1 => n4020, B2 => 
                           n3913, ZN => n3915);
   U1269 : OAI211_X1 port map( C1 => n3917, C2 => n4429, A => n3916, B => n3915
                           , ZN => n3918);
   U1270 : AOI222_X1 port map( A1 => n3920, A2 => n4028, B1 => n3919, B2 => 
                           n4370, C1 => n3918, C2 => n4026, ZN => n3921);
   U1271 : OAI22_X1 port map( A1 => n3922, A2 => n4455, B1 => n3921, B2 => 
                           n4457, ZN => n3926);
   U1272 : OAI22_X1 port map( A1 => n4572, A2 => n3924, B1 => n3923, B2 => 
                           n4459, ZN => n3925);
   U1273 : AOI211_X1 port map( C1 => n4566, C2 => n3927, A => n3926, B => n3925
                           , ZN => n3929);
   U1274 : INV_X1 port map( A => n3928, ZN => n3934);
   U1275 : OAI22_X1 port map( A1 => n4472, A2 => n3929, B1 => n3934, B2 => 
                           n4199, ZN => n3931);
   U1276 : OAI22_X1 port map( A1 => n3941, A2 => n4583, B1 => n3940, B2 => 
                           n4169, ZN => n3930);
   U1277 : AOI211_X1 port map( C1 => n4578, C2 => n3932, A => n3931, B => n3930
                           , ZN => n3938);
   U1278 : INV_X1 port map( A => n3940, ZN => n3937);
   U1279 : OAI22_X1 port map( A1 => n4495, A2 => n3934, B1 => n3933, B2 => 
                           n4169, ZN => n3936);
   U1280 : OAI22_X1 port map( A1 => n3942, A2 => n4583, B1 => n3941, B2 => 
                           n4199, ZN => n3935);
   U1281 : AOI211_X1 port map( C1 => n4578, C2 => n3937, A => n3936, B => n3935
                           , ZN => n3948);
   U1282 : OAI222_X1 port map( A1 => n4131, A2 => n3947, B1 => n4145, B2 => 
                           n3938, C1 => n3948, C2 => n3981, ZN => n3946);
   U1283 : INV_X1 port map( A => n4593, ZN => n4070);
   U1284 : INV_X1 port map( A => n3939, ZN => n3978);
   U1285 : OAI22_X1 port map( A1 => n4495, A2 => n3940, B1 => n3978, B2 => 
                           n4583, ZN => n3944);
   U1286 : OAI22_X1 port map( A1 => n3942, A2 => n4169, B1 => n3941, B2 => 
                           n4492, ZN => n3943);
   U1287 : AOI211_X1 port map( C1 => n4576, C2 => n3945, A => n3944, B => n3943
                           , ZN => n3951);
   U1288 : OAI222_X1 port map( A1 => n4131, A2 => n3951, B1 => n4145, B2 => 
                           n3948, C1 => n3952, C2 => n3981, ZN => n4060);
   U1289 : AOI22_X1 port map( A1 => n4126, A2 => n3946, B1 => n4070, B2 => 
                           n4060, ZN => n3954);
   U1290 : OAI222_X1 port map( A1 => n4131, A2 => n3948, B1 => n4145, B2 => 
                           n3947, C1 => n3951, C2 => n3981, ZN => n3961);
   U1291 : NAND2_X1 port map( A1 => n3950, A2 => n3949, ZN => n4595);
   U1292 : INV_X1 port map( A => n4595, ZN => n4059);
   U1293 : OAI222_X1 port map( A1 => n4131, A2 => n3952, B1 => n4145, B2 => 
                           n3951, C1 => n3982, C2 => n3981, ZN => n4072);
   U1294 : AOI22_X1 port map( A1 => n4602, A2 => n3961, B1 => n4059, B2 => 
                           n4072, ZN => n3953);
   U1295 : OAI211_X1 port map( C1 => n4096, C2 => n4597, A => n3954, B => n3953
                           , ZN => n3959);
   U1296 : INV_X1 port map( A => DATA2_I_31_port, ZN => n3956);
   U1297 : AOI221_X1 port map( B1 => n3957, B2 => n3956, C1 => n3955, C2 => 
                           DATA2_I_31_port, A => DATA1(31), ZN => n3958);
   U1298 : AOI21_X1 port map( B1 => n4509, B2 => n3959, A => n3958, ZN => n3986
                           );
   U1299 : NOR3_X1 port map( A1 => n4831, A2 => n4597, A3 => n3960, ZN => n4791
                           );
   U1300 : AOI22_X1 port map( A1 => n4126, A2 => n3961, B1 => n4070, B2 => 
                           n4072, ZN => n3984);
   U1301 : AOI22_X1 port map( A1 => n4160, A2 => n3963, B1 => n4161, B2 => 
                           n3962, ZN => n3967);
   U1302 : AOI22_X1 port map( A1 => n3403, A2 => n3965, B1 => n4542, B2 => 
                           n3964, ZN => n3966);
   U1303 : OAI211_X1 port map( C1 => n3968, C2 => n4535, A => n3967, B => n3966
                           , ZN => n4507);
   U1304 : AOI22_X1 port map( A1 => n4440, A2 => n4439, B1 => n3969, B2 => 
                           n4507, ZN => n3972);
   U1305 : AOI22_X1 port map( A1 => n4441, A2 => n4427, B1 => n4508, B2 => 
                           n3970, ZN => n3971);
   U1306 : OAI211_X1 port map( C1 => n4475, C2 => n4429, A => n3972, B => n3971
                           , ZN => n4406);
   U1307 : AOI222_X1 port map( A1 => n4406, A2 => n4028, B1 => n4371, B2 => 
                           n4357, C1 => n3973, C2 => n4026, ZN => n4361);
   U1308 : OAI22_X1 port map( A1 => n4572, A2 => n4361, B1 => n4304, B2 => 
                           n4455, ZN => n3977);
   U1309 : OAI22_X1 port map( A1 => n3975, A2 => n4461, B1 => n3974, B2 => 
                           n4419, ZN => n3976);
   U1310 : AOI211_X1 port map( C1 => n4568, C2 => n4341, A => n3977, B => n3976
                           , ZN => n4232);
   U1311 : OAI22_X1 port map( A1 => n4198, A2 => n4199, B1 => n4232, B2 => 
                           n4583, ZN => n3980);
   U1312 : OAI22_X1 port map( A1 => n4495, A2 => n3978, B1 => n4167, B2 => 
                           n4492, ZN => n3979);
   U1313 : AOI211_X1 port map( C1 => n4580, C2 => n4168, A => n3980, B => n3979
                           , ZN => n4146);
   U1314 : OAI222_X1 port map( A1 => n4131, A2 => n4132, B1 => n4145, B2 => 
                           n3982, C1 => n4146, C2 => n3981, ZN => n4125);
   U1315 : AOI22_X1 port map( A1 => n4602, A2 => n4060, B1 => n4288, B2 => 
                           n4125, ZN => n3983);
   U1316 : OAI211_X1 port map( C1 => n4096, C2 => n4595, A => n3984, B => n3983
                           , ZN => n3994);
   U1317 : NAND3_X1 port map( A1 => n4770, A2 => n4791, A3 => n3994, ZN => 
                           n3985);
   U1318 : NAND4_X1 port map( A1 => n3988, A2 => n3987, A3 => n3986, A4 => 
                           n3985, ZN => OUTALU(31));
   U1319 : INV_X1 port map( A => n3989, ZN => n3999);
   U1320 : AOI22_X1 port map( A1 => n4074, A2 => DATA1(31), B1 => n4519, B2 => 
                           DATA1(30), ZN => n3992);
   U1321 : INV_X1 port map( A => DATA2(30), ZN => n4799);
   U1322 : AOI22_X1 port map( A1 => DATA1(30), A2 => DATA2(30), B1 => n4799, B2
                           => n4721, ZN => n4716);
   U1323 : AOI22_X1 port map( A1 => dataout_mul_30_port, A2 => n4491, B1 => 
                           n4778, B2 => n4716, ZN => n3991);
   U1324 : OAI211_X1 port map( C1 => n4511, C2 => n4510, A => DATA1(30), B => 
                           DATA2(30), ZN => n3990);
   U1325 : OAI211_X1 port map( C1 => n3992, C2 => n4794, A => n3991, B => n3990
                           , ZN => n3993);
   U1326 : AOI21_X1 port map( B1 => n4509, B2 => n3994, A => n3993, ZN => n3998
                           );
   U1327 : OAI21_X1 port map( B1 => n3996, B2 => n4000, A => n3995, ZN => n3997
                           );
   U1328 : OAI211_X1 port map( C1 => n4000, C2 => n3999, A => n3998, B => n3997
                           , ZN => OUTALU(30));
   U1329 : AOI22_X1 port map( A1 => n4001, A2 => n4004, B1 => n4779, B2 => 
                           n4002, ZN => n4050);
   U1330 : OAI22_X1 port map( A1 => n4785, A2 => n4004, B1 => n4003, B2 => 
                           n4002, ZN => n4005);
   U1331 : INV_X1 port map( A => n4005, ZN => n4048);
   U1332 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(2), ZN => n4006);
   U1333 : NAND2_X1 port map( A1 => n4074, A2 => DATA1(1), ZN => n4523);
   U1334 : OAI211_X1 port map( C1 => n4007, C2 => n4750, A => n4006, B => n4523
                           , ZN => n4046);
   U1335 : AOI21_X1 port map( B1 => n4781, B2 => DATA1(2), A => n4511, ZN => 
                           n4044);
   U1336 : AOI22_X1 port map( A1 => DATA2(2), A2 => DATA1(2), B1 => n4008, B2 
                           => n4829, ZN => n4753);
   U1337 : AOI22_X1 port map( A1 => dataout_mul_2_port, A2 => n4491, B1 => 
                           n4778, B2 => n4753, ZN => n4043);
   U1338 : OAI22_X1 port map( A1 => n4596, A2 => n4285, B1 => n4598, B2 => 
                           n4593, ZN => n4041);
   U1339 : AOI22_X1 port map( A1 => DATA1(2), A2 => n4519, B1 => DATA1(6), B2 
                           => n4009, ZN => n4013);
   U1340 : NAND4_X1 port map( A1 => n4013, A2 => n4012, A3 => n4011, A4 => 
                           n4010, ZN => n4530);
   U1341 : AOI222_X1 port map( A1 => n4014, A2 => n4260, B1 => n4530, B2 => 
                           n4527, C1 => n4261, C2 => n4525, ZN => n4532);
   U1342 : OAI22_X1 port map( A1 => n4534, A2 => n4532, B1 => n4262, B2 => 
                           n4537, ZN => n4016);
   U1343 : OAI22_X1 port map( A1 => n4264, A2 => n4531, B1 => n4538, B2 => 
                           n4535, ZN => n4015);
   U1344 : AOI211_X1 port map( C1 => n4018, C2 => n4017, A => n4016, B => n4015
                           , ZN => n4546);
   U1345 : INV_X1 port map( A => n4268, ZN => n4553);
   U1346 : AOI22_X1 port map( A1 => n4425, A2 => n4553, B1 => n4020, B2 => 
                           n4019, ZN => n4025);
   U1347 : AOI22_X1 port map( A1 => n4440, A2 => n4023, B1 => n4022, B2 => 
                           n4021, ZN => n4024);
   U1348 : OAI211_X1 port map( C1 => n4546, C2 => n4543, A => n4025, B => n4024
                           , ZN => n4251);
   U1349 : AOI222_X1 port map( A1 => n4029, A2 => n4028, B1 => n4027, B2 => 
                           n4370, C1 => n4251, C2 => n4026, ZN => n4518);
   U1350 : OAI22_X1 port map( A1 => n4571, A2 => n4455, B1 => n4518, B2 => 
                           n4457, ZN => n4033);
   U1351 : OAI22_X1 port map( A1 => n4572, A2 => n4031, B1 => n4030, B2 => 
                           n4459, ZN => n4032);
   U1352 : AOI211_X1 port map( C1 => n4566, C2 => n4567, A => n4033, B => n4032
                           , ZN => n4517);
   U1353 : OAI22_X1 port map( A1 => n4472, A2 => n4517, B1 => n4584, B2 => 
                           n4199, ZN => n4037);
   U1354 : OAI22_X1 port map( A1 => n4035, A2 => n4583, B1 => n4034, B2 => 
                           n4169, ZN => n4036);
   U1355 : AOI211_X1 port map( C1 => n4578, C2 => n4579, A => n4037, B => n4036
                           , ZN => n4038);
   U1356 : INV_X1 port map( A => n4038, ZN => n4590);
   U1357 : AOI222_X1 port map( A1 => n4039, A2 => n4589, B1 => n4284, B2 => 
                           n4587, C1 => n4590, C2 => n4585, ZN => n4594);
   U1358 : OAI22_X1 port map( A1 => n4594, A2 => n4591, B1 => n4250, B2 => 
                           n4595, ZN => n4040);
   U1359 : OAI21_X1 port map( B1 => n4041, B2 => n4040, A => n4506, ZN => n4042
                           );
   U1360 : OAI211_X1 port map( C1 => n4044, C2 => n4829, A => n4043, B => n4042
                           , ZN => n4045);
   U1361 : AOI21_X1 port map( B1 => n4509, B2 => n4046, A => n4045, ZN => n4047
                           );
   U1362 : OAI221_X1 port map( B1 => n4051, B2 => n4050, C1 => n4049, C2 => 
                           n4048, A => n4047, ZN => OUTALU(2));
   U1363 : AOI22_X1 port map( A1 => n4150, A2 => n4078, B1 => n4156, B2 => 
                           n4079, ZN => n4068);
   U1364 : INV_X1 port map( A => DATA2(29), ZN => n4800);
   U1365 : AOI211_X1 port map( C1 => n4470, C2 => n4471, A => n4052, B => n4800
                           , ZN => n4057);
   U1366 : NOR2_X1 port map( A1 => DATA2(29), A2 => n4052, ZN => n4646);
   U1367 : NAND2_X1 port map( A1 => DATA2(29), A2 => n4052, ZN => n4643);
   U1368 : INV_X1 port map( A => n4643, ZN => n4717);
   U1369 : NOR2_X1 port map( A1 => n4646, A2 => n4717, ZN => n4760);
   U1370 : NOR2_X1 port map( A1 => n4248, A2 => n4052, ZN => n4054);
   U1371 : AOI211_X1 port map( C1 => DATA1(31), C2 => n4520, A => n4054, B => 
                           n4053, ZN => n4055);
   U1372 : OAI22_X1 port map( A1 => n4760, A2 => n4479, B1 => n4055, B2 => 
                           n4794, ZN => n4056);
   U1373 : AOI211_X1 port map( C1 => dataout_mul_29_port, C2 => n4491, A => 
                           n4057, B => n4056, ZN => n4067);
   U1374 : INV_X1 port map( A => n4058, ZN => n4064);
   U1375 : AOI22_X1 port map( A1 => n4602, A2 => n4072, B1 => n4070, B2 => 
                           n4071, ZN => n4062);
   U1376 : AOI22_X1 port map( A1 => n4126, A2 => n4060, B1 => n4059, B2 => 
                           n4125, ZN => n4061);
   U1377 : AOI21_X1 port map( B1 => n4062, B2 => n4061, A => n4467, ZN => n4063
                           );
   U1378 : AOI221_X1 port map( B1 => n4065, B2 => n4064, C1 => n4069, C2 => 
                           n4064, A => n4063, ZN => n4066);
   U1379 : OAI211_X1 port map( C1 => n4069, C2 => n4068, A => n4067, B => n4066
                           , ZN => OUTALU(29));
   U1380 : AOI222_X1 port map( A1 => n4072, A2 => n4126, B1 => n4071, B2 => 
                           n4602, C1 => n4125, C2 => n4070, ZN => n4094);
   U1381 : AOI22_X1 port map( A1 => n4074, A2 => DATA1(29), B1 => n4073, B2 => 
                           DATA1(30), ZN => n4076);
   U1382 : NAND2_X1 port map( A1 => n4258, A2 => DATA1(28), ZN => n4075);
   U1383 : OAI211_X1 port map( C1 => n4723, C2 => n4077, A => n4076, B => n4075
                           , ZN => n4089);
   U1384 : OR2_X1 port map( A1 => n4133, A2 => n4078, ZN => n4081);
   U1385 : NOR2_X1 port map( A1 => n4135, A2 => n4079, ZN => n4083);
   U1386 : INV_X1 port map( A => n4083, ZN => n4080);
   U1387 : AOI22_X1 port map( A1 => n4082, A2 => n4090, B1 => n4081, B2 => 
                           n4080, ZN => n4088);
   U1388 : INV_X1 port map( A => DATA2(28), ZN => n4801);
   U1389 : AOI22_X1 port map( A1 => DATA1(28), A2 => DATA2(28), B1 => n4801, B2
                           => n4642, ZN => n4730);
   U1390 : INV_X1 port map( A => n4730, ZN => n4714);
   U1391 : INV_X1 port map( A => n4103, ZN => n4084);
   U1392 : AOI22_X1 port map( A1 => n4491, A2 => dataout_mul_28_port, B1 => 
                           n4084, B2 => n4083, ZN => n4086);
   U1393 : NAND3_X1 port map( A1 => DATA2(28), A2 => DATA1(28), A3 => n4450, ZN
                           => n4085);
   U1394 : OAI211_X1 port map( C1 => n4714, C2 => n4479, A => n4086, B => n4085
                           , ZN => n4087);
   U1395 : AOI211_X1 port map( C1 => n4506, C2 => n4089, A => n4088, B => n4087
                           , ZN => n4093);
   U1396 : INV_X1 port map( A => n4105, ZN => n4091);
   U1397 : NAND3_X1 port map( A1 => n4091, A2 => n4150, A3 => n4090, ZN => 
                           n4092);
   U1398 : OAI211_X1 port map( C1 => n4094, C2 => n4467, A => n4093, B => n4092
                           , ZN => OUTALU(28));
   U1399 : INV_X1 port map( A => n4125, ZN => n4095);
   U1400 : OAI22_X1 port map( A1 => n4096, A2 => n4591, B1 => n4095, B2 => 
                           n4285, ZN => n4102);
   U1401 : NOR3_X1 port map( A1 => n4114, A2 => n4794, A3 => n4113, ZN => n4101
                           );
   U1402 : INV_X1 port map( A => DATA2(27), ZN => n4802);
   U1403 : NAND2_X1 port map( A1 => n4802, A2 => DATA1(27), ZN => n4711);
   U1404 : NAND2_X1 port map( A1 => n4097, A2 => DATA2(27), ZN => n4713);
   U1405 : OAI21_X1 port map( B1 => n4471, B2 => n4802, A => n4470, ZN => n4098
                           );
   U1406 : AOI22_X1 port map( A1 => DATA1(27), A2 => n4098, B1 => n4476, B2 => 
                           dataout_mul_27_port, ZN => n4099);
   U1407 : OAI221_X1 port map( B1 => n4479, B2 => n4711, C1 => n4479, C2 => 
                           n4713, A => n4099, ZN => n4100);
   U1408 : AOI211_X1 port map( C1 => n4509, C2 => n4102, A => n4101, B => n4100
                           , ZN => n4110);
   U1409 : OAI211_X1 port map( C1 => n4107, C2 => n4104, A => n4156, B => n4103
                           , ZN => n4109);
   U1410 : OAI211_X1 port map( C1 => n4107, C2 => n4106, A => n4150, B => n4105
                           , ZN => n4108);
   U1411 : NAND3_X1 port map( A1 => n4110, A2 => n4109, A3 => n4108, ZN => 
                           OUTALU(27));
   U1412 : INV_X1 port map( A => DATA2(26), ZN => n4803);
   U1413 : NOR3_X1 port map( A1 => n4111, A2 => n4803, A3 => n4712, ZN => n4119
                           );
   U1414 : OAI22_X1 port map( A1 => n4712, A2 => DATA2(26), B1 => n4803, B2 => 
                           DATA1(26), ZN => n4707);
   U1415 : OAI22_X1 port map( A1 => n4115, A2 => n4114, B1 => n4113, B2 => 
                           n4112, ZN => n4116);
   U1416 : AOI22_X1 port map( A1 => n4707, A2 => n4372, B1 => n4116, B2 => 
                           n4506, ZN => n4117);
   U1417 : INV_X1 port map( A => n4117, ZN => n4118);
   U1418 : AOI211_X1 port map( C1 => n4789, C2 => dataout_mul_26_port, A => 
                           n4119, B => n4118, ZN => n4130);
   U1419 : OR2_X1 port map( A1 => n4121, A2 => n4120, ZN => n4124);
   U1420 : OAI211_X1 port map( C1 => n4136, C2 => n4124, A => n4156, B => n4122
                           , ZN => n4129);
   U1421 : OAI211_X1 port map( C1 => n4134, C2 => n4124, A => n4150, B => n4123
                           , ZN => n4128);
   U1422 : NAND3_X1 port map( A1 => n4509, A2 => n4126, A3 => n4125, ZN => 
                           n4127);
   U1423 : NAND4_X1 port map( A1 => n4130, A2 => n4129, A3 => n4128, A4 => 
                           n4127, ZN => OUTALU(26));
   U1424 : INV_X1 port map( A => DATA2(25), ZN => n4804);
   U1425 : AOI22_X1 port map( A1 => DATA1(25), A2 => DATA2(25), B1 => n4804, B2
                           => n4708, ZN => n4740);
   U1426 : AOI22_X1 port map( A1 => n4740, A2 => n4372, B1 => n4491, B2 => 
                           dataout_mul_25_port, ZN => n4144);
   U1427 : OAI22_X1 port map( A1 => n4132, A2 => n4145, B1 => n4146, B2 => 
                           n4131, ZN => n4140);
   U1428 : AOI211_X1 port map( C1 => n4149, C2 => n4137, A => n4134, B => n4133
                           , ZN => n4139);
   U1429 : AOI211_X1 port map( C1 => n4157, C2 => n4137, A => n4136, B => n4135
                           , ZN => n4138);
   U1430 : AOI211_X1 port map( C1 => n4509, C2 => n4140, A => n4139, B => n4138
                           , ZN => n4143);
   U1431 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n4450, ZN
                           => n4142);
   U1432 : NAND3_X1 port map( A1 => n4506, A2 => n4161, A3 => n4197, ZN => 
                           n4141);
   U1433 : NAND4_X1 port map( A1 => n4144, A2 => n4143, A3 => n4142, A4 => 
                           n4141, ZN => OUTALU(25));
   U1434 : AOI22_X1 port map( A1 => DATA2(24), A2 => n4510, B1 => 
                           DATA2_I_24_port, B2 => n4156, ZN => n4159);
   U1435 : NOR3_X1 port map( A1 => n4146, A2 => n4467, A3 => n4145, ZN => n4155
                           );
   U1436 : AOI22_X1 port map( A1 => n4147, A2 => n4197, B1 => n4161, B2 => 
                           n4195, ZN => n4153);
   U1437 : INV_X1 port map( A => DATA2(24), ZN => n4805);
   U1438 : OAI22_X1 port map( A1 => n4636, A2 => DATA2(24), B1 => n4805, B2 => 
                           DATA1(24), ZN => n4732);
   U1439 : AOI22_X1 port map( A1 => dataout_mul_24_port, A2 => n4491, B1 => 
                           n4778, B2 => n4732, ZN => n4152);
   U1440 : INV_X1 port map( A => n4157, ZN => n4148);
   U1441 : NAND3_X1 port map( A1 => n4150, A2 => n4149, A3 => n4148, ZN => 
                           n4151);
   U1442 : OAI211_X1 port map( C1 => n4153, C2 => n4794, A => n4152, B => n4151
                           , ZN => n4154);
   U1443 : AOI211_X1 port map( C1 => n4157, C2 => n4156, A => n4155, B => n4154
                           , ZN => n4158);
   U1444 : OAI221_X1 port map( B1 => n4636, B2 => n4159, C1 => n4636, C2 => 
                           n4470, A => n4158, ZN => OUTALU(24));
   U1445 : INV_X1 port map( A => DATA2(23), ZN => n4806);
   U1446 : NAND2_X1 port map( A1 => DATA1(23), A2 => n4806, ZN => n4632);
   U1447 : NAND2_X1 port map( A1 => DATA2(23), A2 => n4163, ZN => n4705);
   U1448 : AOI21_X1 port map( B1 => n4632, B2 => n4705, A => n4479, ZN => n4166
                           );
   U1449 : AOI21_X1 port map( B1 => n4510, B2 => DATA2(23), A => n4511, ZN => 
                           n4164);
   U1450 : AOI222_X1 port map( A1 => n4194, A2 => n4161, B1 => n4197, B2 => 
                           n4160, C1 => n4195, C2 => n3837, ZN => n4162);
   U1451 : OAI22_X1 port map( A1 => n4164, A2 => n4163, B1 => n4162, B2 => 
                           n4794, ZN => n4165);
   U1452 : AOI211_X1 port map( C1 => n4789, C2 => dataout_mul_23_port, A => 
                           n4166, B => n4165, ZN => n4191);
   U1453 : OAI22_X1 port map( A1 => n4495, A2 => n4167, B1 => n4198, B2 => 
                           n4492, ZN => n4171);
   U1454 : INV_X1 port map( A => n4168, ZN => n4215);
   U1455 : OAI22_X1 port map( A1 => n4215, A2 => n4199, B1 => n4232, B2 => 
                           n4169, ZN => n4170);
   U1456 : OAI21_X1 port map( B1 => n4171, B2 => n4170, A => n4509, ZN => n4190
                           );
   U1457 : INV_X1 port map( A => n4182, ZN => n4181);
   U1458 : NAND2_X1 port map( A1 => n4797, A2 => n4180, ZN => n4329);
   U1459 : OAI21_X1 port map( B1 => n4350, B2 => n4349, A => n4172, ZN => n4330
                           );
   U1460 : AND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n4173);
   U1461 : AOI21_X1 port map( B1 => n4330, B2 => n4336, A => n4173, ZN => n4302
                           );
   U1462 : OAI21_X1 port map( B1 => n4175, B2 => n4302, A => n4174, ZN => n4229
                           );
   U1463 : INV_X1 port map( A => n4176, ZN => n4177);
   U1464 : AOI21_X1 port map( B1 => n4229, B2 => n4237, A => n4177, ZN => n4213
                           );
   U1465 : OAI21_X1 port map( B1 => n4224, B2 => n4213, A => n4178, ZN => n4179
                           );
   U1466 : INV_X1 port map( A => n4179, ZN => n4184);
   U1467 : NOR2_X1 port map( A1 => n5139, A2 => n4180, ZN => n4364);
   U1468 : INV_X1 port map( A => n4364, ZN => n4328);
   U1469 : OAI22_X1 port map( A1 => n4181, A2 => n4329, B1 => n4184, B2 => 
                           n4328, ZN => n4200);
   U1470 : NAND3_X1 port map( A1 => n4201, A2 => n4186, A3 => n4200, ZN => 
                           n4189);
   U1471 : OAI21_X1 port map( B1 => n4182, B2 => n4329, A => n4201, ZN => n4183
                           );
   U1472 : AOI21_X1 port map( B1 => n4364, B2 => n4184, A => n4183, ZN => n4206
                           );
   U1473 : OAI21_X1 port map( B1 => n4206, B2 => n4186, A => n4187, ZN => n4185
                           );
   U1474 : OAI211_X1 port map( C1 => n4187, C2 => n4186, A => n4797, B => n4185
                           , ZN => n4188);
   U1475 : NAND4_X1 port map( A1 => n4191, A2 => n4190, A3 => n4189, A4 => 
                           n4188, ZN => OUTALU(23));
   U1476 : AOI22_X1 port map( A1 => n4147, A2 => n4194, B1 => n4193, B2 => 
                           n4192, ZN => n4211);
   U1477 : AOI22_X1 port map( A1 => n3403, A2 => n4197, B1 => n4196, B2 => 
                           n4195, ZN => n4210);
   U1478 : OAI222_X1 port map( A1 => n4199, A2 => n4232, B1 => n4492, B2 => 
                           n4215, C1 => n4198, C2 => n4472, ZN => n4208);
   U1479 : NOR2_X1 port map( A1 => n4201, A2 => n4200, ZN => n4205);
   U1480 : INV_X1 port map( A => DATA2(22), ZN => n4807);
   U1481 : AOI22_X1 port map( A1 => DATA1(22), A2 => DATA2(22), B1 => n4807, B2
                           => n4202, ZN => n4629);
   U1482 : AOI22_X1 port map( A1 => dataout_mul_22_port, A2 => n4491, B1 => 
                           n4778, B2 => n4629, ZN => n4204);
   U1483 : NAND3_X1 port map( A1 => DATA2(22), A2 => DATA1(22), A3 => n4450, ZN
                           => n4203);
   U1484 : OAI211_X1 port map( C1 => n4206, C2 => n4205, A => n4204, B => n4203
                           , ZN => n4207);
   U1485 : AOI21_X1 port map( B1 => n4509, B2 => n4208, A => n4207, ZN => n4209
                           );
   U1486 : OAI221_X1 port map( B1 => n4794, B2 => n4211, C1 => n4794, C2 => 
                           n4210, A => n4209, ZN => OUTALU(22));
   U1487 : INV_X1 port map( A => n4224, ZN => n4226);
   U1488 : OAI22_X1 port map( A1 => n4328, A2 => n4213, B1 => n4329, B2 => 
                           n4214, ZN => n4212);
   U1489 : INV_X1 port map( A => n4212, ZN => n4225);
   U1490 : INV_X1 port map( A => n4329, ZN => n4366);
   U1491 : AOI22_X1 port map( A1 => n4214, A2 => n4366, B1 => n4364, B2 => 
                           n4213, ZN => n4223);
   U1492 : OAI22_X1 port map( A1 => n4472, A2 => n4215, B1 => n4232, B2 => 
                           n4492, ZN => n4221);
   U1493 : AOI21_X1 port map( B1 => n4781, B2 => DATA2(21), A => n4511, ZN => 
                           n4219);
   U1494 : INV_X1 port map( A => DATA2(21), ZN => n4808);
   U1495 : NAND2_X1 port map( A1 => n4808, A2 => DATA1(21), ZN => n4698);
   U1496 : NAND2_X1 port map( A1 => n4218, A2 => DATA2(21), ZN => n4700);
   U1497 : NAND2_X1 port map( A1 => n4698, A2 => n4700, ZN => n4739);
   U1498 : AOI22_X1 port map( A1 => dataout_mul_21_port, A2 => n4491, B1 => 
                           n4778, B2 => n4739, ZN => n4217);
   U1499 : NAND3_X1 port map( A1 => n4506, A2 => n4426, A3 => n4320, ZN => 
                           n4216);
   U1500 : OAI211_X1 port map( C1 => n4219, C2 => n4218, A => n4217, B => n4216
                           , ZN => n4220);
   U1501 : AOI21_X1 port map( B1 => n4509, B2 => n4221, A => n4220, ZN => n4222
                           );
   U1502 : OAI221_X1 port map( B1 => n4226, B2 => n4225, C1 => n4224, C2 => 
                           n4223, A => n4222, ZN => OUTALU(21));
   U1503 : AOI21_X1 port map( B1 => n4781, B2 => DATA2(20), A => n4511, ZN => 
                           n4241);
   U1504 : NOR2_X1 port map( A1 => n4240, A2 => DATA2(20), ZN => n4703);
   U1505 : AOI21_X1 port map( B1 => DATA2(20), B2 => n4240, A => n4703, ZN => 
                           n4649);
   U1506 : AOI22_X1 port map( A1 => n4441, A2 => n4320, B1 => n4508, B2 => 
                           n4321, ZN => n4227);
   U1507 : OAI22_X1 port map( A1 => n4649, A2 => n4479, B1 => n4227, B2 => 
                           n4794, ZN => n4228);
   U1508 : AOI21_X1 port map( B1 => n4789, B2 => dataout_mul_20_port, A => 
                           n4228, ZN => n4239);
   U1509 : OAI22_X1 port map( A1 => n4230, A2 => n4329, B1 => n4328, B2 => 
                           n4229, ZN => n4236);
   U1510 : AOI22_X1 port map( A1 => n4230, A2 => n4366, B1 => n4229, B2 => 
                           n4364, ZN => n4231);
   U1511 : INV_X1 port map( A => n4231, ZN => n4234);
   U1512 : NOR3_X1 port map( A1 => n4472, A2 => n4232, A3 => n4467, ZN => n4233
                           );
   U1513 : AOI221_X1 port map( B1 => n4237, B2 => n4236, C1 => n4235, C2 => 
                           n4234, A => n4233, ZN => n4238);
   U1514 : OAI211_X1 port map( C1 => n4241, C2 => n4240, A => n4239, B => n4238
                           , ZN => OUTALU(20));
   U1515 : NOR3_X1 port map( A1 => n4242, A2 => n4750, A3 => n4467, ZN => n4243
                           );
   U1516 : AOI21_X1 port map( B1 => n4789, B2 => dataout_mul_1_port, A => n4243
                           , ZN => n4298);
   U1517 : NAND2_X1 port map( A1 => DATA1(1), A2 => n4830, ZN => n4657);
   U1518 : NOR2_X1 port map( A1 => DATA1(1), A2 => n4830, ZN => n4659);
   U1519 : INV_X1 port map( A => n4659, ZN => n4244);
   U1520 : NAND2_X1 port map( A1 => n4657, A2 => n4244, ZN => n4737);
   U1521 : INV_X1 port map( A => n4776, ZN => n4246);
   U1522 : AOI221_X1 port map( B1 => n4246, B2 => n4294, C1 => n4776, C2 => 
                           n4245, A => n4785, ZN => n4247);
   U1523 : AOI21_X1 port map( B1 => n4372, B2 => n4737, A => n4247, ZN => n4297
                           );
   U1524 : OAI21_X1 port map( B1 => n4467, B2 => n4248, A => n4470, ZN => n4782
                           );
   U1525 : AOI21_X1 port map( B1 => DATA2(1), B2 => n4510, A => n4782, ZN => 
                           n4249);
   U1526 : INV_X1 port map( A => n4249, ZN => n4291);
   U1527 : INV_X1 port map( A => n4250, ZN => n4289);
   U1528 : INV_X1 port map( A => n4251, ZN => n4556);
   U1529 : INV_X1 port map( A => n4546, ZN => n4272);
   U1530 : INV_X1 port map( A => n4532, ZN => n4267);
   U1531 : OAI211_X1 port map( C1 => n4255, C2 => n4254, A => n4253, B => n4252
                           , ZN => n4256);
   U1532 : AOI211_X1 port map( C1 => DATA1(1), C2 => n4258, A => n4257, B => 
                           n4256, ZN => n4259);
   U1533 : INV_X1 port map( A => n4259, ZN => n4526);
   U1534 : AOI222_X1 port map( A1 => n4527, A2 => n4526, B1 => n4525, B2 => 
                           n4530, C1 => n4261, C2 => n4260, ZN => n4536);
   U1535 : OAI22_X1 port map( A1 => n4531, A2 => n4538, B1 => n4534, B2 => 
                           n4536, ZN => n4266);
   U1536 : OAI22_X1 port map( A1 => n4537, A2 => n4264, B1 => n4263, B2 => 
                           n4262, ZN => n4265);
   U1537 : AOI211_X1 port map( C1 => n4267, C2 => n4147, A => n4266, B => n4265
                           , ZN => n4548);
   U1538 : OAI22_X1 port map( A1 => n4545, A2 => n4268, B1 => n4543, B2 => 
                           n4548, ZN => n4271);
   U1539 : OAI22_X1 port map( A1 => n4429, A2 => n4549, B1 => n4550, B2 => 
                           n4269, ZN => n4270);
   U1540 : AOI211_X1 port map( C1 => n4272, C2 => n4425, A => n4271, B => n4270
                           , ZN => n4559);
   U1541 : OAI222_X1 port map( A1 => n4273, A2 => n4555, B1 => n4556, B2 => 
                           n4560, C1 => n4559, C2 => n4558, ZN => n4565);
   U1542 : AOI22_X1 port map( A1 => n4567, A2 => n4564, B1 => n4565, B2 => 
                           n4562, ZN => n4278);
   U1543 : INV_X1 port map( A => n4571, ZN => n4274);
   U1544 : AOI22_X1 port map( A1 => n4276, A2 => n4275, B1 => n4274, B2 => 
                           n4568, ZN => n4277);
   U1545 : OAI211_X1 port map( C1 => n4461, C2 => n4518, A => n4278, B => n4277
                           , ZN => n4577);
   U1546 : AOI22_X1 port map( A1 => n4579, A2 => n4576, B1 => n4574, B2 => 
                           n4577, ZN => n4283);
   U1547 : AOI22_X1 port map( A1 => n4281, A2 => n4580, B1 => n4280, B2 => 
                           n4279, ZN => n4282);
   U1548 : OAI211_X1 port map( C1 => n4492, C2 => n4517, A => n4283, B => n4282
                           , ZN => n4588);
   U1549 : AOI222_X1 port map( A1 => n4587, A2 => n4590, B1 => n4585, B2 => 
                           n4588, C1 => n4284, C2 => n4589, ZN => n4516);
   U1550 : OAI22_X1 port map( A1 => n4595, A2 => n4598, B1 => n4591, B2 => 
                           n4516, ZN => n4287);
   U1551 : OAI22_X1 port map( A1 => n4285, A2 => n4594, B1 => n4593, B2 => 
                           n4596, ZN => n4286);
   U1552 : AOI211_X1 port map( C1 => n4289, C2 => n4288, A => n4287, B => n4286
                           , ZN => n4290);
   U1553 : INV_X1 port map( A => n4290, ZN => n4790);
   U1554 : AOI22_X1 port map( A1 => DATA1(1), A2 => n4291, B1 => n4506, B2 => 
                           n4790, ZN => n4296);
   U1555 : OR2_X1 port map( A1 => n4780, A2 => DATA2_I_0_port, ZN => n4293);
   U1556 : OAI211_X1 port map( C1 => n4294, C2 => n4293, A => n4779, B => n4292
                           , ZN => n4295);
   U1557 : NAND4_X1 port map( A1 => n4298, A2 => n4297, A3 => n4296, A4 => 
                           n4295, ZN => OUTALU(1));
   U1558 : INV_X1 port map( A => DATA2(19), ZN => n4810);
   U1559 : AOI221_X1 port map( B1 => n4510, B2 => DATA2(19), C1 => n4372, C2 =>
                           n4810, A => n4511, ZN => n4316);
   U1560 : AOI222_X1 port map( A1 => n4321, A2 => n4441, B1 => n4320, B2 => 
                           n4440, C1 => n4319, C2 => n4426, ZN => n4299);
   U1561 : NOR2_X1 port map( A1 => n4810, A2 => DATA1(19), ZN => n4625);
   U1562 : INV_X1 port map( A => n4625, ZN => n4648);
   U1563 : OAI22_X1 port map( A1 => n4299, A2 => n4794, B1 => n4648, B2 => 
                           n4479, ZN => n4300);
   U1564 : AOI21_X1 port map( B1 => n4789, B2 => dataout_mul_19_port, A => 
                           n4300, ZN => n4314);
   U1565 : AOI22_X1 port map( A1 => n4303, A2 => n4366, B1 => n4364, B2 => 
                           n4302, ZN => n4301);
   U1566 : INV_X1 port map( A => n4301, ZN => n4311);
   U1567 : INV_X1 port map( A => n4312, ZN => n4310);
   U1568 : OAI22_X1 port map( A1 => n4303, A2 => n4329, B1 => n4302, B2 => 
                           n4328, ZN => n4309);
   U1569 : INV_X1 port map( A => n4304, ZN => n4317);
   U1570 : AOI22_X1 port map( A1 => n4562, A2 => n4305, B1 => n4566, B2 => 
                           n4317, ZN => n4307);
   U1571 : INV_X1 port map( A => n4361, ZN => n4340);
   U1572 : AOI22_X1 port map( A1 => n4564, A2 => n4341, B1 => n4568, B2 => 
                           n4340, ZN => n4306);
   U1573 : AOI21_X1 port map( B1 => n4307, B2 => n4306, A => n4467, ZN => n4308
                           );
   U1574 : AOI221_X1 port map( B1 => n4312, B2 => n4311, C1 => n4310, C2 => 
                           n4309, A => n4308, ZN => n4313);
   U1575 : OAI211_X1 port map( C1 => n4316, C2 => n4315, A => n4314, B => n4313
                           , ZN => OUTALU(19));
   U1576 : AOI222_X1 port map( A1 => n4340, A2 => n4564, B1 => n4317, B2 => 
                           n4562, C1 => n4341, C2 => n4566, ZN => n4339);
   U1577 : AOI22_X1 port map( A1 => n4425, A2 => n4319, B1 => n4508, B2 => 
                           n4318, ZN => n4323);
   U1578 : AOI22_X1 port map( A1 => n4440, A2 => n4321, B1 => n4554, B2 => 
                           n4320, ZN => n4322);
   U1579 : AOI21_X1 port map( B1 => n4323, B2 => n4322, A => n4794, ZN => n4327
                           );
   U1580 : NOR2_X1 port map( A1 => n4324, A2 => DATA2(18), ZN => n4650);
   U1581 : INV_X1 port map( A => DATA2(18), ZN => n4811);
   U1582 : NOR2_X1 port map( A1 => n4811, A2 => DATA1(18), ZN => n4764);
   U1583 : NOR2_X1 port map( A1 => n4650, A2 => n4764, ZN => n4695);
   U1584 : AOI21_X1 port map( B1 => n4781, B2 => DATA2(18), A => n4511, ZN => 
                           n4325);
   U1585 : OAI22_X1 port map( A1 => n4695, A2 => n4479, B1 => n4325, B2 => 
                           n4324, ZN => n4326);
   U1586 : AOI211_X1 port map( C1 => dataout_mul_18_port, C2 => n4491, A => 
                           n4327, B => n4326, ZN => n4338);
   U1587 : OAI22_X1 port map( A1 => n4331, A2 => n4329, B1 => n4328, B2 => 
                           n4330, ZN => n4335);
   U1588 : AOI22_X1 port map( A1 => n4331, A2 => n4366, B1 => n4330, B2 => 
                           n4364, ZN => n4332);
   U1589 : INV_X1 port map( A => n4332, ZN => n4334);
   U1590 : AOI22_X1 port map( A1 => n4336, A2 => n4335, B1 => n4334, B2 => 
                           n4333, ZN => n4337);
   U1591 : OAI211_X1 port map( C1 => n4339, C2 => n4467, A => n4338, B => n4337
                           , ZN => OUTALU(18));
   U1592 : AOI22_X1 port map( A1 => n4562, A2 => n4341, B1 => n4566, B2 => 
                           n4340, ZN => n4355);
   U1593 : NOR2_X1 port map( A1 => DATA2(17), A2 => n4342, ZN => n4697);
   U1594 : INV_X1 port map( A => n4697, ZN => n4627);
   U1595 : NAND2_X1 port map( A1 => DATA2(17), A2 => n4342, ZN => n4694);
   U1596 : NAND2_X1 port map( A1 => n4627, A2 => n4694, ZN => n4738);
   U1597 : AOI22_X1 port map( A1 => dataout_mul_17_port, A2 => n4491, B1 => 
                           n4778, B2 => n4738, ZN => n4348);
   U1598 : AND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n4344);
   U1599 : OAI211_X1 port map( C1 => n4344, C2 => n4352, A => n4366, B => n4343
                           , ZN => n4347);
   U1600 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n4450, ZN
                           => n4346);
   U1601 : NAND3_X1 port map( A1 => n4506, A2 => n4407, A3 => n4356, ZN => 
                           n4345);
   U1602 : AND4_X1 port map( A1 => n4348, A2 => n4347, A3 => n4346, A4 => n4345
                           , ZN => n4354);
   U1603 : INV_X1 port map( A => n4349, ZN => n4351);
   U1604 : OAI221_X1 port map( B1 => n4352, B2 => n4351, C1 => n4350, C2 => 
                           n4349, A => n4364, ZN => n4353);
   U1605 : OAI211_X1 port map( C1 => n4355, C2 => n4467, A => n4354, B => n4353
                           , ZN => OUTALU(17));
   U1606 : INV_X1 port map( A => DATA2(16), ZN => n4813);
   U1607 : AOI221_X1 port map( B1 => n4781, B2 => DATA2(16), C1 => n4372, C2 =>
                           n4813, A => n4511, ZN => n4369);
   U1608 : AOI22_X1 port map( A1 => n4407, A2 => n4358, B1 => n4357, B2 => 
                           n4356, ZN => n4359);
   U1609 : NAND2_X1 port map( A1 => DATA2(16), A2 => n4603, ZN => n4652);
   U1610 : OAI22_X1 port map( A1 => n4359, A2 => n4794, B1 => n4652, B2 => 
                           n4479, ZN => n4360);
   U1611 : AOI21_X1 port map( B1 => n4789, B2 => dataout_mul_16_port, A => 
                           n4360, ZN => n4368);
   U1612 : INV_X1 port map( A => n4365, ZN => n4363);
   U1613 : NOR3_X1 port map( A1 => n4361, A2 => n4467, A3 => n4419, ZN => n4362
                           );
   U1614 : AOI221_X1 port map( B1 => n4366, B2 => n4365, C1 => n4364, C2 => 
                           n4363, A => n4362, ZN => n4367);
   U1615 : OAI211_X1 port map( C1 => n4369, C2 => n4603, A => n4368, B => n4367
                           , ZN => OUTALU(16));
   U1616 : AOI22_X1 port map( A1 => n4407, A2 => n4371, B1 => n4370, B2 => 
                           n4406, ZN => n4396);
   U1617 : NOR3_X1 port map( A1 => n4460, A2 => n4794, A3 => n4457, ZN => n4389
                           );
   U1618 : NAND2_X1 port map( A1 => DATA2(15), A2 => n4621, ZN => n4653);
   U1619 : INV_X1 port map( A => DATA2(15), ZN => n4814);
   U1620 : OAI221_X1 port map( B1 => DATA2(15), B2 => n4372, C1 => n4814, C2 =>
                           n4450, A => DATA1(15), ZN => n4387);
   U1621 : INV_X1 port map( A => n4373, ZN => n4377);
   U1622 : INV_X1 port map( A => n4374, ZN => n4376);
   U1623 : NOR2_X1 port map( A1 => n4376, A2 => n4375, ZN => n4498);
   U1624 : NOR2_X1 port map( A1 => n4498, A2 => n4501, ZN => n4497);
   U1625 : NOR2_X1 port map( A1 => n4377, A2 => n4497, ZN => n4469);
   U1626 : OAI21_X1 port map( B1 => n4379, B2 => n4469, A => n4378, ZN => n4448
                           );
   U1627 : AOI21_X1 port map( B1 => n4381, B2 => n4448, A => n4380, ZN => n4399
                           );
   U1628 : NAND2_X1 port map( A1 => n4399, A2 => n4402, ZN => n4398);
   U1629 : INV_X1 port map( A => n4398, ZN => n4383);
   U1630 : OAI21_X1 port map( B1 => n4383, B2 => n4415, A => n4382, ZN => n4385
                           );
   U1631 : AOI21_X1 port map( B1 => n4393, B2 => n4385, A => n4496, ZN => n4384
                           );
   U1632 : OAI21_X1 port map( B1 => n4393, B2 => n4385, A => n4384, ZN => n4386
                           );
   U1633 : OAI211_X1 port map( C1 => n4479, C2 => n4653, A => n4387, B => n4386
                           , ZN => n4388);
   U1634 : AOI211_X1 port map( C1 => n4789, C2 => dataout_mul_15_port, A => 
                           n4389, B => n4388, ZN => n4395);
   U1635 : INV_X1 port map( A => n4390, ZN => n4392);
   U1636 : INV_X1 port map( A => n4499, ZN => n4483);
   U1637 : OAI221_X1 port map( B1 => n4393, B2 => n4392, C1 => n4391, C2 => 
                           n4390, A => n4483, ZN => n4394);
   U1638 : OAI211_X1 port map( C1 => n4396, C2 => n4467, A => n4395, B => n4394
                           , ZN => OUTALU(15));
   U1639 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           ZN => n5063);
   U1640 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A => n5063, ZN => n5064);
   U1641 : NAND2_X1 port map( A1 => n5064, A2 => 
                           boothmul_pipelined_i_muxes_in_7_233_port, ZN => 
                           n4404);
   U1642 : NOR2_X1 port map( A1 => n4404, A2 => n5126, ZN => n3087);
   U1643 : INV_X1 port map( A => n4496, ZN => n4447);
   U1644 : AOI22_X1 port map( A1 => n4447, A2 => n4398, B1 => n4483, B2 => 
                           n4397, ZN => n4416);
   U1645 : AOI22_X1 port map( A1 => n4400, A2 => n4483, B1 => n4447, B2 => 
                           n4399, ZN => n4420);
   U1646 : INV_X1 port map( A => n4420, ZN => n4401);
   U1647 : NAND2_X1 port map( A1 => n4402, A2 => n4401, ZN => n4414);
   U1648 : OAI22_X1 port map( A1 => n4456, A2 => n4419, B1 => n4460, B2 => 
                           n4461, ZN => n4412);
   U1649 : AOI211_X1 port map( C1 => n4404, C2 => n5126, A => n3087, B => n4403
                           , ZN => n4411);
   U1650 : NOR2_X1 port map( A1 => DATA2(14), A2 => n4405, ZN => n4654);
   U1651 : NAND2_X1 port map( A1 => DATA2(14), A2 => n4405, ZN => n4618);
   U1652 : INV_X1 port map( A => n4618, ZN => n4765);
   U1653 : NOR2_X1 port map( A1 => n4654, A2 => n4765, ZN => n4689);
   U1654 : OAI211_X1 port map( C1 => n4511, C2 => n4510, A => n5138, B => 
                           DATA2(14), ZN => n4409);
   U1655 : NAND3_X1 port map( A1 => n4509, A2 => n4407, A3 => n4406, ZN => 
                           n4408);
   U1656 : OAI211_X1 port map( C1 => n4689, C2 => n4479, A => n4409, B => n4408
                           , ZN => n4410);
   U1657 : AOI211_X1 port map( C1 => n4506, C2 => n4412, A => n4411, B => n4410
                           , ZN => n4413);
   U1658 : OAI221_X1 port map( B1 => n4417, B2 => n4416, C1 => n4415, C2 => 
                           n4414, A => n4413, ZN => OUTALU(14));
   U1659 : INV_X1 port map( A => n4444, ZN => n4449);
   U1660 : NAND2_X1 port map( A1 => n4449, A2 => n4448, ZN => n4446);
   U1661 : OAI211_X1 port map( C1 => n4443, C2 => n4418, A => n4797, B => n4421
                           , ZN => n4438);
   U1662 : OAI222_X1 port map( A1 => n4419, A2 => n4462, B1 => n4461, B2 => 
                           n4456, C1 => n4455, C2 => n4460, ZN => n4436);
   U1663 : AOI21_X1 port map( B1 => n4422, B2 => n4421, A => n4420, ZN => n4435
                           );
   U1664 : NOR2_X1 port map( A1 => DATA2(13), A2 => n4423, ZN => n4691);
   U1665 : NOR2_X1 port map( A1 => DATA1(13), A2 => n4816, ZN => n4687);
   U1666 : NOR2_X1 port map( A1 => n4691, A2 => n4687, ZN => n4758);
   U1667 : OAI21_X1 port map( B1 => n4471, B2 => n4816, A => n4470, ZN => n4424
                           );
   U1668 : AOI22_X1 port map( A1 => DATA1(13), A2 => n4424, B1 => n4476, B2 => 
                           dataout_mul_13_port, ZN => n4433);
   U1669 : AOI22_X1 port map( A1 => n4427, A2 => n4426, B1 => n4439, B2 => 
                           n4425, ZN => n4428);
   U1670 : INV_X1 port map( A => n4428, ZN => n4431);
   U1671 : INV_X1 port map( A => n4507, ZN => n4474);
   U1672 : OAI22_X1 port map( A1 => n4475, A2 => n4545, B1 => n4474, B2 => 
                           n4429, ZN => n4430);
   U1673 : OAI21_X1 port map( B1 => n4431, B2 => n4430, A => n4509, ZN => n4432
                           );
   U1674 : OAI211_X1 port map( C1 => n4758, C2 => n4479, A => n4433, B => n4432
                           , ZN => n4434);
   U1675 : AOI211_X1 port map( C1 => n4506, C2 => n4436, A => n4435, B => n4434
                           , ZN => n4437);
   U1676 : OAI21_X1 port map( B1 => n4446, B2 => n4438, A => n4437, ZN => 
                           OUTALU(13));
   U1677 : AOI222_X1 port map( A1 => n4442, A2 => n4441, B1 => n4507, B2 => 
                           n4440, C1 => n4439, C2 => n4508, ZN => n4468);
   U1678 : INV_X1 port map( A => n4443, ZN => n4445);
   U1679 : AOI221_X1 port map( B1 => n4445, B2 => n4444, C1 => n4443, C2 => 
                           n4449, A => n4499, ZN => n4454);
   U1680 : OAI22_X1 port map( A1 => n4686, A2 => DATA2(12), B1 => n4817, B2 => 
                           DATA1(12), ZN => n4751);
   U1681 : INV_X1 port map( A => n4751, ZN => n4683);
   U1682 : OAI211_X1 port map( C1 => n4449, C2 => n4448, A => n4447, B => n4446
                           , ZN => n4452);
   U1683 : NAND3_X1 port map( A1 => DATA2(12), A2 => DATA1(12), A3 => n4450, ZN
                           => n4451);
   U1684 : OAI211_X1 port map( C1 => n4683, C2 => n4479, A => n4452, B => n4451
                           , ZN => n4453);
   U1685 : AOI211_X1 port map( C1 => n4789, C2 => dataout_mul_12_port, A => 
                           n4454, B => n4453, ZN => n4466);
   U1686 : OAI22_X1 port map( A1 => n4458, A2 => n4457, B1 => n4456, B2 => 
                           n4455, ZN => n4464);
   U1687 : OAI22_X1 port map( A1 => n4462, A2 => n4461, B1 => n4460, B2 => 
                           n4459, ZN => n4463);
   U1688 : OAI21_X1 port map( B1 => n4464, B2 => n4463, A => n4506, ZN => n4465
                           );
   U1689 : OAI211_X1 port map( C1 => n4468, C2 => n4467, A => n4466, B => n4465
                           , ZN => OUTALU(12));
   U1690 : XNOR2_X1 port map( A => n4469, B => n4486, ZN => n4490);
   U1691 : OAI21_X1 port map( B1 => n4471, B2 => n4473, A => n4470, ZN => n4482
                           );
   U1692 : NOR3_X1 port map( A1 => n4472, A2 => n4493, A3 => n4794, ZN => n4481
                           );
   U1693 : NAND2_X1 port map( A1 => DATA1(11), A2 => n4818, ZN => n4680);
   U1694 : NAND2_X1 port map( A1 => DATA2(11), A2 => n4473, ZN => n4682);
   U1695 : OAI22_X1 port map( A1 => n4475, A2 => n4543, B1 => n4474, B2 => 
                           n4547, ZN => n4477);
   U1696 : AOI22_X1 port map( A1 => n4509, A2 => n4477, B1 => n4476, B2 => 
                           dataout_mul_11_port, ZN => n4478);
   U1697 : OAI221_X1 port map( B1 => n4479, B2 => n4680, C1 => n4479, C2 => 
                           n4682, A => n4478, ZN => n4480);
   U1698 : AOI211_X1 port map( C1 => DATA2(11), C2 => n4482, A => n4481, B => 
                           n4480, ZN => n4489);
   U1699 : INV_X1 port map( A => n4487, ZN => n4485);
   U1700 : INV_X1 port map( A => n4486, ZN => n4484);
   U1701 : OAI221_X1 port map( B1 => n4487, B2 => n4486, C1 => n4485, C2 => 
                           n4484, A => n4483, ZN => n4488);
   U1702 : OAI211_X1 port map( C1 => n4490, C2 => n4496, A => n4489, B => n4488
                           , ZN => OUTALU(11));
   U1703 : AOI22_X1 port map( A1 => DATA1(10), A2 => DATA2(10), B1 => n4819, B2
                           => n4681, ZN => n4677);
   U1704 : AOI22_X1 port map( A1 => dataout_mul_10_port, A2 => n4491, B1 => 
                           n4778, B2 => n4677, ZN => n4515);
   U1705 : OAI22_X1 port map( A1 => n4495, A2 => n4494, B1 => n4493, B2 => 
                           n4492, ZN => n4505);
   U1706 : AOI211_X1 port map( C1 => n4498, C2 => n4501, A => n4497, B => n4496
                           , ZN => n4504);
   U1707 : AOI211_X1 port map( C1 => n4502, C2 => n4501, A => n4500, B => n4499
                           , ZN => n4503);
   U1708 : AOI211_X1 port map( C1 => n4506, C2 => n4505, A => n4504, B => n4503
                           , ZN => n4514);
   U1709 : NAND3_X1 port map( A1 => n4509, A2 => n4508, A3 => n4507, ZN => 
                           n4513);
   U1710 : OAI211_X1 port map( C1 => n4511, C2 => n4510, A => DATA2(10), B => 
                           n5137, ZN => n4512);
   U1711 : NAND4_X1 port map( A1 => n4515, A2 => n4514, A3 => n4513, A4 => 
                           n4512, ZN => OUTALU(10));
   U1712 : INV_X1 port map( A => n4516, ZN => n4601);
   U1713 : INV_X1 port map( A => n4517, ZN => n4575);
   U1714 : INV_X1 port map( A => n4518, ZN => n4563);
   U1715 : AOI22_X1 port map( A1 => n4520, A2 => DATA1(2), B1 => n4519, B2 => 
                           n4780, ZN => n4524);
   U1716 : NAND4_X1 port map( A1 => n4524, A2 => n4523, A3 => n4522, A4 => 
                           n4521, ZN => n4528);
   U1717 : AOI222_X1 port map( A1 => n4530, A2 => n4529, B1 => n4528, B2 => 
                           n4527, C1 => n4526, C2 => n4525, ZN => n4533);
   U1718 : OAI22_X1 port map( A1 => n4534, A2 => n4533, B1 => n4532, B2 => 
                           n4531, ZN => n4540);
   U1719 : OAI22_X1 port map( A1 => n4538, A2 => n4537, B1 => n4536, B2 => 
                           n4535, ZN => n4539);
   U1720 : AOI211_X1 port map( C1 => n4542, C2 => n4541, A => n4540, B => n4539
                           , ZN => n4544);
   U1721 : OAI22_X1 port map( A1 => n4546, A2 => n4545, B1 => n4544, B2 => 
                           n4543, ZN => n4552);
   U1722 : OAI22_X1 port map( A1 => n4550, A2 => n4549, B1 => n4548, B2 => 
                           n4547, ZN => n4551);
   U1723 : AOI211_X1 port map( C1 => n4554, C2 => n4553, A => n4552, B => n4551
                           , ZN => n4557);
   U1724 : OAI222_X1 port map( A1 => n4560, A2 => n4559, B1 => n4558, B2 => 
                           n4557, C1 => n4556, C2 => n4555, ZN => n4561);
   U1725 : AOI22_X1 port map( A1 => n4564, A2 => n4563, B1 => n4562, B2 => 
                           n4561, ZN => n4570);
   U1726 : AOI22_X1 port map( A1 => n4568, A2 => n4567, B1 => n4566, B2 => 
                           n4565, ZN => n4569);
   U1727 : OAI211_X1 port map( C1 => n4572, C2 => n4571, A => n4570, B => n4569
                           , ZN => n4573);
   U1728 : AOI22_X1 port map( A1 => n4576, A2 => n4575, B1 => n4574, B2 => 
                           n4573, ZN => n4582);
   U1729 : AOI22_X1 port map( A1 => n4580, A2 => n4579, B1 => n4578, B2 => 
                           n4577, ZN => n4581);
   U1730 : OAI211_X1 port map( C1 => n4584, C2 => n4583, A => n4582, B => n4581
                           , ZN => n4586);
   U1731 : AOI222_X1 port map( A1 => n4590, A2 => n4589, B1 => n4588, B2 => 
                           n4587, C1 => n4586, C2 => n4585, ZN => n4592);
   U1732 : OAI22_X1 port map( A1 => n4594, A2 => n4593, B1 => n4592, B2 => 
                           n4591, ZN => n4600);
   U1733 : OAI22_X1 port map( A1 => n4598, A2 => n4597, B1 => n4596, B2 => 
                           n4595, ZN => n4599);
   U1734 : AOI211_X1 port map( C1 => n4602, C2 => n4601, A => n4600, B => n4599
                           , ZN => n4795);
   U1735 : OAI21_X1 port map( B1 => n4803, B2 => DATA1(26), A => n4713, ZN => 
                           n4742);
   U1736 : INV_X1 port map( A => DATA2(20), ZN => n4809);
   U1737 : OAI21_X1 port map( B1 => n4809, B2 => DATA1(20), A => n4700, ZN => 
                           n4631);
   U1738 : NOR2_X1 port map( A1 => DATA2(16), A2 => n4603, ZN => n4651);
   U1739 : AOI21_X1 port map( B1 => DATA2(12), B2 => n4686, A => n4687, ZN => 
                           n4617);
   U1740 : AOI21_X1 port map( B1 => DATA2(6), B2 => n4604, A => n4672, ZN => 
                           n4727);
   U1741 : NOR2_X1 port map( A1 => DATA1(0), A2 => n4831, ZN => n4605);
   U1742 : AOI21_X1 port map( B1 => n4605, B2 => n4657, A => n4659, ZN => n4606
                           );
   U1743 : OAI22_X1 port map( A1 => DATA1(2), A2 => n4829, B1 => n4606, B2 => 
                           n4753, ZN => n4607);
   U1744 : OAI211_X1 port map( C1 => n4662, C2 => n4607, A => n4664, B => n4667
                           , ZN => n4608);
   U1745 : NAND3_X1 port map( A1 => n4609, A2 => n4668, A3 => n4608, ZN => 
                           n4610);
   U1746 : NAND3_X1 port map( A1 => n4669, A2 => n4666, A3 => n4610, ZN => 
                           n4611);
   U1747 : AOI211_X1 port map( C1 => n4727, C2 => n4611, A => n4656, B => n4756
                           , ZN => n4612);
   U1748 : AOI21_X1 port map( B1 => DATA2(8), B2 => n4655, A => n4612, ZN => 
                           n4614);
   U1749 : AOI211_X1 port map( C1 => n4614, C2 => n4674, A => n4613, B => n4677
                           , ZN => n4615);
   U1750 : OAI21_X1 port map( B1 => n5137, B2 => n4819, A => n4682, ZN => n4744
                           );
   U1751 : OAI211_X1 port map( C1 => n4615, C2 => n4744, A => n4683, B => n4680
                           , ZN => n4616);
   U1752 : AOI211_X1 port map( C1 => n4617, C2 => n4616, A => n4691, B => n4654
                           , ZN => n4620);
   U1753 : NAND2_X1 port map( A1 => n4618, A2 => n4653, ZN => n4619);
   U1754 : OAI22_X1 port map( A1 => DATA2(15), A2 => n4621, B1 => n4620, B2 => 
                           n4619, ZN => n4622);
   U1755 : OAI211_X1 port map( C1 => n4651, C2 => n4622, A => n4694, B => n4652
                           , ZN => n4623);
   U1756 : INV_X1 port map( A => n4623, ZN => n4624);
   U1757 : NOR2_X1 port map( A1 => n4650, A2 => n4624, ZN => n4626);
   U1758 : AOI211_X1 port map( C1 => n4627, C2 => n4626, A => n4625, B => n4764
                           , ZN => n4628);
   U1759 : AOI211_X1 port map( C1 => n4810, C2 => DATA1(19), A => n4703, B => 
                           n4628, ZN => n4630);
   U1760 : INV_X1 port map( A => n4629, ZN => n4701);
   U1761 : OAI211_X1 port map( C1 => n4631, C2 => n4630, A => n4698, B => n4701
                           , ZN => n4634);
   U1762 : OAI21_X1 port map( B1 => DATA1(22), B2 => n4807, A => n4705, ZN => 
                           n4743);
   U1763 : INV_X1 port map( A => n4743, ZN => n4633);
   U1764 : INV_X1 port map( A => n4632, ZN => n4647);
   U1765 : AOI211_X1 port map( C1 => n4634, C2 => n4633, A => n4732, B => n4647
                           , ZN => n4635);
   U1766 : AOI21_X1 port map( B1 => n4636, B2 => DATA2(24), A => n4635, ZN => 
                           n4638);
   U1767 : OR2_X1 port map( A1 => n4638, A2 => DATA1(25), ZN => n4637);
   U1768 : AOI221_X1 port map( B1 => n4638, B2 => DATA1(25), C1 => n4804, C2 =>
                           n4637, A => n4707, ZN => n4639);
   U1769 : OAI211_X1 port map( C1 => n4742, C2 => n4639, A => n4711, B => n4714
                           , ZN => n4640);
   U1770 : INV_X1 port map( A => n4640, ZN => n4641);
   U1771 : AOI21_X1 port map( B1 => DATA2(28), B2 => n4642, A => n4641, ZN => 
                           n4644);
   U1772 : AOI211_X1 port map( C1 => n4644, C2 => n4643, A => n4646, B => n4716
                           , ZN => n4645);
   U1773 : OAI22_X1 port map( A1 => DATA1(30), A2 => n4799, B1 => DATA2(31), B2
                           => n4723, ZN => n4741);
   U1774 : NAND2_X1 port map( A1 => DATA2(31), A2 => n4723, ZN => n4720);
   U1775 : OAI21_X1 port map( B1 => n4645, B2 => n4741, A => n4720, ZN => n4726
                           );
   U1776 : AOI21_X1 port map( B1 => DATA1(28), B2 => n4801, A => n4646, ZN => 
                           n4719);
   U1777 : AOI21_X1 port map( B1 => DATA1(22), B2 => n4807, A => n4647, ZN => 
                           n4734);
   U1778 : NAND2_X1 port map( A1 => n4649, A2 => n4648, ZN => n4755);
   U1779 : AOI21_X1 port map( B1 => DATA1(19), B2 => n4810, A => n4650, ZN => 
                           n4735);
   U1780 : INV_X1 port map( A => n4651, ZN => n4692);
   U1781 : NAND3_X1 port map( A1 => n4692, A2 => n4653, A3 => n4652, ZN => 
                           n4763);
   U1782 : AOI21_X1 port map( B1 => DATA1(15), B2 => n4814, A => n4654, ZN => 
                           n4736);
   U1783 : NOR2_X1 port map( A1 => DATA2(8), A2 => n4655, ZN => n4676);
   U1784 : AOI21_X1 port map( B1 => DATA1(6), B2 => n4825, A => n4656, ZN => 
                           n4749);
   U1785 : INV_X1 port map( A => n4753, ZN => n4661);
   U1786 : NAND2_X1 port map( A1 => n4780, A2 => n4831, ZN => n4658);
   U1787 : OAI21_X1 port map( B1 => n4659, B2 => n4658, A => n4657, ZN => n4660
                           );
   U1788 : AOI22_X1 port map( A1 => n4661, A2 => n4660, B1 => DATA1(2), B2 => 
                           n4829, ZN => n4665);
   U1789 : AOI211_X1 port map( C1 => n4665, C2 => n4664, A => n4663, B => n4662
                           , ZN => n4671);
   U1790 : NAND2_X1 port map( A1 => n4667, A2 => n4666, ZN => n4670);
   U1791 : OAI211_X1 port map( C1 => n4671, C2 => n4670, A => n4669, B => n4668
                           , ZN => n4673);
   U1792 : AOI211_X1 port map( C1 => n4749, C2 => n4673, A => n4672, B => n4756
                           , ZN => n4675);
   U1793 : OAI21_X1 port map( B1 => n4676, B2 => n4675, A => n4674, ZN => n4678
                           );
   U1794 : AOI21_X1 port map( B1 => n4679, B2 => n4678, A => n4677, ZN => n4684
                           );
   U1795 : OAI21_X1 port map( B1 => DATA2(10), B2 => n4681, A => n4680, ZN => 
                           n4752);
   U1796 : OAI211_X1 port map( C1 => n4684, C2 => n4752, A => n4683, B => n4682
                           , ZN => n4685);
   U1797 : OAI21_X1 port map( B1 => DATA2(12), B2 => n4686, A => n4685, ZN => 
                           n4690);
   U1798 : INV_X1 port map( A => n4687, ZN => n4688);
   U1799 : OAI211_X1 port map( C1 => n4691, C2 => n4690, A => n4689, B => n4688
                           , ZN => n4693);
   U1800 : OAI221_X1 port map( B1 => n4763, B2 => n4736, C1 => n4763, C2 => 
                           n4693, A => n4692, ZN => n4696);
   U1801 : OAI211_X1 port map( C1 => n4697, C2 => n4696, A => n4695, B => n4694
                           , ZN => n4699);
   U1802 : OAI221_X1 port map( B1 => n4755, B2 => n4735, C1 => n4755, C2 => 
                           n4699, A => n4698, ZN => n4702);
   U1803 : OAI211_X1 port map( C1 => n4703, C2 => n4702, A => n4701, B => n4700
                           , ZN => n4704);
   U1804 : AOI21_X1 port map( B1 => n4734, B2 => n4704, A => n4732, ZN => n4706
                           );
   U1805 : AOI22_X1 port map( A1 => DATA1(24), A2 => n4805, B1 => n4706, B2 => 
                           n4705, ZN => n4709);
   U1806 : OR2_X1 port map( A1 => n4709, A2 => n4708, ZN => n4710);
   U1807 : AOI221_X1 port map( B1 => DATA2(25), B2 => n4710, C1 => n4709, C2 =>
                           n4708, A => n4707, ZN => n4715);
   U1808 : OAI21_X1 port map( B1 => DATA2(26), B2 => n4712, A => n4711, ZN => 
                           n4731);
   U1809 : OAI211_X1 port map( C1 => n4715, C2 => n4731, A => n4714, B => n4713
                           , ZN => n4718);
   U1810 : AOI211_X1 port map( C1 => n4719, C2 => n4718, A => n4717, B => n4716
                           , ZN => n4722);
   U1811 : OAI21_X1 port map( B1 => DATA2(30), B2 => n4721, A => n4720, ZN => 
                           n4729);
   U1812 : OAI22_X1 port map( A1 => DATA2(31), A2 => n4723, B1 => n4722, B2 => 
                           n4729, ZN => n4725);
   U1813 : OAI221_X1 port map( B1 => FUNC(3), B2 => n4726, C1 => n4796, C2 => 
                           n4725, A => n4724, ZN => n4775);
   U1814 : INV_X1 port map( A => n4727, ZN => n4728);
   U1815 : NOR4_X1 port map( A1 => n4731, A2 => n4730, A3 => n4729, A4 => n4728
                           , ZN => n4748);
   U1816 : INV_X1 port map( A => n4732, ZN => n4733);
   U1817 : AND4_X1 port map( A1 => n4736, A2 => n4735, A3 => n4734, A4 => n4733
                           , ZN => n4747);
   U1818 : NOR4_X1 port map( A1 => n4740, A2 => n4739, A3 => n4738, A4 => n4737
                           , ZN => n4746);
   U1819 : NOR4_X1 port map( A1 => n4744, A2 => n4743, A3 => n4742, A4 => n4741
                           , ZN => n4745);
   U1820 : NAND4_X1 port map( A1 => n4748, A2 => n4747, A3 => n4746, A4 => 
                           n4745, ZN => n4772);
   U1821 : INV_X1 port map( A => n4749, ZN => n4757);
   U1822 : OAI22_X1 port map( A1 => n4831, A2 => n4780, B1 => n4750, B2 => 
                           DATA2(0), ZN => n4777);
   U1823 : OR4_X1 port map( A1 => n4753, A2 => n4752, A3 => n4751, A4 => n4777,
                           ZN => n4754);
   U1824 : NOR4_X1 port map( A1 => n4757, A2 => n4756, A3 => n4755, A4 => n4754
                           , ZN => n4769);
   U1825 : NAND4_X1 port map( A1 => n4761, A2 => n4760, A3 => n4759, A4 => 
                           n4758, ZN => n4762);
   U1826 : NOR4_X1 port map( A1 => n4765, A2 => n4764, A3 => n4763, A4 => n4762
                           , ZN => n4766);
   U1827 : NAND4_X1 port map( A1 => n4769, A2 => n4768, A3 => n4767, A4 => 
                           n4766, ZN => n4771);
   U1828 : OAI21_X1 port map( B1 => n4772, B2 => n4771, A => n4770, ZN => n4774
                           );
   U1829 : AOI211_X1 port map( C1 => n4775, C2 => n4774, A => FUNC(1), B => 
                           n4773, ZN => n4788);
   U1830 : OAI21_X1 port map( B1 => DATA1(0), B2 => DATA2_I_0_port, A => n4776,
                           ZN => n4786);
   U1831 : AOI22_X1 port map( A1 => n4779, A2 => n4786, B1 => n4778, B2 => 
                           n4777, ZN => n4784);
   U1832 : OAI221_X1 port map( B1 => n4782, B2 => DATA2(0), C1 => n4782, C2 => 
                           n4781, A => n4780, ZN => n4783);
   U1833 : OAI211_X1 port map( C1 => n4786, C2 => n4785, A => n4784, B => n4783
                           , ZN => n4787);
   U1834 : AOI211_X1 port map( C1 => n4789, C2 => dataout_mul_0_port, A => 
                           n4788, B => n4787, ZN => n4793);
   U1835 : NAND4_X1 port map( A1 => FUNC(2), A2 => FUNC(3), A3 => n4791, A4 => 
                           n4790, ZN => n4792);
   U1836 : OAI211_X1 port map( C1 => n4795, C2 => n4794, A => n4793, B => n4792
                           , ZN => OUTALU(0));
   U1837 : NAND2_X1 port map( A1 => n4797, A2 => n4796, ZN => n4833);
   U1838 : CLKBUF_X1 port map( A => n4833, Z => n4823);
   U1839 : NAND2_X1 port map( A1 => FUNC(3), A2 => n4797, ZN => n4832);
   U1840 : AOI22_X1 port map( A1 => DATA2(31), A2 => n4823, B1 => n4822, B2 => 
                           n4798, ZN => N2548);
   U1841 : AOI22_X1 port map( A1 => DATA2(30), A2 => n4833, B1 => n4832, B2 => 
                           n4799, ZN => N2547);
   U1842 : AOI22_X1 port map( A1 => DATA2(29), A2 => n4823, B1 => n4822, B2 => 
                           n4800, ZN => N2546);
   U1843 : AOI22_X1 port map( A1 => DATA2(28), A2 => n4833, B1 => n4832, B2 => 
                           n4801, ZN => N2545);
   U1844 : AOI22_X1 port map( A1 => DATA2(27), A2 => n4823, B1 => n4822, B2 => 
                           n4802, ZN => N2544);
   U1845 : AOI22_X1 port map( A1 => DATA2(26), A2 => n4833, B1 => n4832, B2 => 
                           n4803, ZN => N2543);
   U1846 : AOI22_X1 port map( A1 => DATA2(25), A2 => n4823, B1 => n4822, B2 => 
                           n4804, ZN => N2542);
   U1847 : AOI22_X1 port map( A1 => DATA2(24), A2 => n4833, B1 => n4832, B2 => 
                           n4805, ZN => N2541);
   U1848 : AOI22_X1 port map( A1 => DATA2(23), A2 => n4823, B1 => n4822, B2 => 
                           n4806, ZN => N2540);
   U1849 : AOI22_X1 port map( A1 => DATA2(22), A2 => n4833, B1 => n4832, B2 => 
                           n4807, ZN => N2539);
   U1850 : AOI22_X1 port map( A1 => DATA2(21), A2 => n4833, B1 => n4832, B2 => 
                           n4808, ZN => N2538);
   U1851 : AOI22_X1 port map( A1 => DATA2(20), A2 => n4833, B1 => n4832, B2 => 
                           n4809, ZN => N2537);
   U1852 : AOI22_X1 port map( A1 => DATA2(19), A2 => n4823, B1 => n4822, B2 => 
                           n4810, ZN => N2536);
   U1853 : AOI22_X1 port map( A1 => DATA2(18), A2 => n4823, B1 => n4822, B2 => 
                           n4811, ZN => N2535);
   U1854 : INV_X1 port map( A => DATA2(17), ZN => n4812);
   U1855 : AOI22_X1 port map( A1 => DATA2(17), A2 => n4823, B1 => n4822, B2 => 
                           n4812, ZN => N2534);
   U1856 : AOI22_X1 port map( A1 => DATA2(16), A2 => n4823, B1 => n4822, B2 => 
                           n4813, ZN => N2533);
   U1857 : AOI22_X1 port map( A1 => DATA2(15), A2 => n4823, B1 => n4822, B2 => 
                           n4814, ZN => N2532);
   U1858 : INV_X1 port map( A => DATA2(14), ZN => n4815);
   U1859 : AOI22_X1 port map( A1 => DATA2(14), A2 => n4823, B1 => n4822, B2 => 
                           n4815, ZN => N2531);
   U1860 : AOI22_X1 port map( A1 => DATA2(13), A2 => n4823, B1 => n4822, B2 => 
                           n4816, ZN => N2530);
   U1861 : AOI22_X1 port map( A1 => DATA2(12), A2 => n4823, B1 => n4822, B2 => 
                           n4817, ZN => N2529);
   U1862 : AOI22_X1 port map( A1 => DATA2(11), A2 => n4823, B1 => n4822, B2 => 
                           n4818, ZN => N2528);
   U1863 : AOI22_X1 port map( A1 => DATA2(10), A2 => n4823, B1 => n4822, B2 => 
                           n4819, ZN => N2527);
   U1864 : AOI22_X1 port map( A1 => DATA2(9), A2 => n4823, B1 => n4822, B2 => 
                           n4820, ZN => N2526);
   U1865 : AOI22_X1 port map( A1 => DATA2(8), A2 => n4823, B1 => n4822, B2 => 
                           n4821, ZN => N2525);
   U1866 : AOI22_X1 port map( A1 => DATA2(7), A2 => n4833, B1 => n4832, B2 => 
                           n4824, ZN => N2524);
   U1867 : AOI22_X1 port map( A1 => DATA2(6), A2 => n4833, B1 => n4832, B2 => 
                           n4825, ZN => N2523);
   U1868 : AOI22_X1 port map( A1 => DATA2(5), A2 => n4833, B1 => n4832, B2 => 
                           n4826, ZN => N2522);
   U1869 : AOI22_X1 port map( A1 => DATA2(4), A2 => n4833, B1 => n4832, B2 => 
                           n4827, ZN => N2521);
   U1870 : AOI22_X1 port map( A1 => DATA2(3), A2 => n4833, B1 => n4832, B2 => 
                           n4828, ZN => N2520);
   U1871 : AOI22_X1 port map( A1 => DATA2(2), A2 => n4833, B1 => n4832, B2 => 
                           n4829, ZN => N2519);
   U1872 : AOI22_X1 port map( A1 => DATA2(1), A2 => n4833, B1 => n4832, B2 => 
                           n4830, ZN => N2518);
   U1873 : AOI22_X1 port map( A1 => DATA2(0), A2 => n4833, B1 => n4832, B2 => 
                           n4831, ZN => N2517);
   U1874 : NOR2_X1 port map( A1 => n4834, A2 => n1994, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1875 : NAND2_X1 port map( A1 => n4875, A2 => data2_mul_3_port, ZN => n4838)
                           ;
   U1876 : INV_X1 port map( A => data2_mul_3_port, ZN => n4871);
   U1877 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n4871, ZN => n4870);
   U1878 : INV_X1 port map( A => n4835, ZN => n4836);
   U1879 : NOR2_X1 port map( A1 => n4836, A2 => n4871, ZN => n4873);
   U1880 : NOR2_X1 port map( A1 => data2_mul_3_port, A2 => n4836, ZN => n4863);
   U1881 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n4873, B1 => data1_mul_1_port, B2 => n4863, ZN
                           => n4837);
   U1882 : OAI221_X1 port map( B1 => n1994, B2 => n4838, C1 => n1994, C2 => 
                           n4870, A => n4837, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1883 : INV_X1 port map( A => n4838, ZN => n4872);
   U1884 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n4863, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n4872, ZN => n4840);
   U1885 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n4873, ZN => n4839);
   U1886 : OAI211_X1 port map( C1 => n1993, C2 => n4870, A => n4840, B => n4839
                           , ZN => boothmul_pipelined_i_mux_out_1_4_port);
   U1887 : CLKBUF_X1 port map( A => n4863, Z => n4867);
   U1888 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n4872, B1 => n4867, B2 => data1_mul_3_port, ZN
                           => n4842);
   U1889 : CLKBUF_X1 port map( A => n4873, Z => n4864);
   U1890 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n4841);
   U1891 : OAI211_X1 port map( C1 => n4870, C2 => n1992, A => n4842, B => n4841
                           , ZN => boothmul_pipelined_i_mux_out_1_5_port);
   U1892 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n4867, B2 => data1_mul_4_port, ZN => n4844);
   U1893 : NAND2_X1 port map( A1 => n4873, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n4843);
   U1894 : OAI211_X1 port map( C1 => n1991, C2 => n4870, A => n4844, B => n4843
                           , ZN => boothmul_pipelined_i_mux_out_1_6_port);
   U1895 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n4867, B2 => data1_mul_5_port, ZN => n4846);
   U1896 : NAND2_X1 port map( A1 => n4873, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n4845);
   U1897 : OAI211_X1 port map( C1 => n1990, C2 => n4870, A => n4846, B => n4845
                           , ZN => boothmul_pipelined_i_mux_out_1_7_port);
   U1898 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n4867, B2 => data1_mul_6_port, ZN => n4848);
   U1899 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n4847);
   U1900 : OAI211_X1 port map( C1 => n1989, C2 => n4870, A => n4848, B => n4847
                           , ZN => boothmul_pipelined_i_mux_out_1_8_port);
   U1901 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n4863, B2 => data1_mul_7_port, ZN => n4850);
   U1902 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n4849);
   U1903 : OAI211_X1 port map( C1 => n1988, C2 => n4870, A => n4850, B => n4849
                           , ZN => boothmul_pipelined_i_mux_out_1_9_port);
   U1904 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n4863, B2 => data1_mul_8_port, ZN => n4852);
   U1905 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n4851);
   U1906 : OAI211_X1 port map( C1 => n1987, C2 => n4870, A => n4852, B => n4851
                           , ZN => boothmul_pipelined_i_mux_out_1_10_port);
   U1907 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n4867, B2 => data1_mul_9_port, ZN => n4854);
   U1908 : NAND2_X1 port map( A1 => n4873, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n4853);
   U1909 : OAI211_X1 port map( C1 => n1986, C2 => n4870, A => n4854, B => n4853
                           , ZN => boothmul_pipelined_i_mux_out_1_11_port);
   U1910 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n4863, B2 => data1_mul_10_port, ZN => n4856);
   U1911 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n4855);
   U1912 : OAI211_X1 port map( C1 => n1985, C2 => n4870, A => n4856, B => n4855
                           , ZN => boothmul_pipelined_i_mux_out_1_12_port);
   U1913 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n4867, B2 => data1_mul_11_port, ZN => n4858);
   U1914 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n4857);
   U1915 : OAI211_X1 port map( C1 => n1984, C2 => n4870, A => n4858, B => n4857
                           , ZN => boothmul_pipelined_i_mux_out_1_13_port);
   U1916 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n4867, B2 => data1_mul_12_port, ZN => n4860);
   U1917 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n4859);
   U1918 : OAI211_X1 port map( C1 => n1983, C2 => n4870, A => n4860, B => n4859
                           , ZN => boothmul_pipelined_i_mux_out_1_14_port);
   U1919 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n4863, B2 => data1_mul_13_port, ZN => n4862);
   U1920 : NAND2_X1 port map( A1 => n4873, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n4861);
   U1921 : OAI211_X1 port map( C1 => n1982, C2 => n4870, A => n4862, B => n4861
                           , ZN => boothmul_pipelined_i_mux_out_1_15_port);
   U1922 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n4863, B2 => data1_mul_14_port, ZN => n4866);
   U1923 : NAND2_X1 port map( A1 => n4864, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n4865);
   U1924 : OAI211_X1 port map( C1 => n1981, C2 => n4870, A => n4866, B => n4865
                           , ZN => boothmul_pipelined_i_mux_out_1_16_port);
   U1925 : AOI22_X1 port map( A1 => n4872, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n4867, B2 => data1_mul_15_port, ZN => n4869);
   U1926 : NAND2_X1 port map( A1 => n4873, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n4868);
   U1927 : OAI211_X1 port map( C1 => n1980, C2 => n4870, A => n4869, B => n4868
                           , ZN => boothmul_pipelined_i_mux_out_1_17_port);
   U1928 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n4871, ZN => n4876
                           );
   U1929 : AOI22_X1 port map( A1 => n4873, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n4872, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n4874);
   U1930 : OAI21_X1 port map( B1 => n4876, B2 => n4875, A => n4874, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1931 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n4915);
   U1932 : NAND2_X1 port map( A1 => n4915, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n4879);
   U1933 : NAND3_X1 port map( A1 => n3076, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n4911);
   U1934 : NOR2_X1 port map( A1 => n3076, A2 => n4877, ZN => n4892);
   U1935 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4877, ZN => n4905);
   U1936 : CLKBUF_X1 port map( A => n4905, Z => n4908);
   U1937 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n4892, B1 => data1_mul_1_port, B2 => n4908, ZN
                           => n4878);
   U1938 : OAI221_X1 port map( B1 => n1994, B2 => n4879, C1 => n1994, C2 => 
                           n4911, A => n4878, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1939 : INV_X1 port map( A => n4879, ZN => n4913);
   U1940 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n4905, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n4913, ZN => n4881);
   U1941 : CLKBUF_X1 port map( A => n4892, Z => n4912);
   U1942 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n4912, ZN => n4880);
   U1943 : OAI211_X1 port map( C1 => n4911, C2 => n1993, A => n4881, B => n4880
                           , ZN => boothmul_pipelined_i_mux_out_2_6_port);
   U1944 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n4913, B1 => data1_mul_3_port, B2 => n4908, ZN
                           => n4883);
   U1945 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n4892, ZN => n4882);
   U1946 : OAI211_X1 port map( C1 => n4911, C2 => n1992, A => n4883, B => n4882
                           , ZN => boothmul_pipelined_i_mux_out_2_7_port);
   U1947 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n4913, B1 => data1_mul_4_port, B2 => n4908, ZN
                           => n4885);
   U1948 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n4892, ZN => n4884);
   U1949 : OAI211_X1 port map( C1 => n4911, C2 => n1991, A => n4885, B => n4884
                           , ZN => boothmul_pipelined_i_mux_out_2_8_port);
   U1950 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n4913, B1 => data1_mul_5_port, B2 => n4905, ZN
                           => n4887);
   U1951 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n4892, ZN => n4886);
   U1952 : OAI211_X1 port map( C1 => n4911, C2 => n1990, A => n4887, B => n4886
                           , ZN => boothmul_pipelined_i_mux_out_2_9_port);
   U1953 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n4913, B1 => data1_mul_6_port, B2 => n4908, ZN
                           => n4889);
   U1954 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n4892, ZN => n4888);
   U1955 : OAI211_X1 port map( C1 => n4911, C2 => n1989, A => n4889, B => n4888
                           , ZN => boothmul_pipelined_i_mux_out_2_10_port);
   U1956 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n4913, B1 => data1_mul_7_port, B2 => n4905, ZN
                           => n4891);
   U1957 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n4892, ZN => n4890);
   U1958 : OAI211_X1 port map( C1 => n4911, C2 => n1988, A => n4891, B => n4890
                           , ZN => boothmul_pipelined_i_mux_out_2_11_port);
   U1959 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n4913, B1 => data1_mul_8_port, B2 => n4908, ZN
                           => n4894);
   U1960 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n4892, ZN => n4893);
   U1961 : OAI211_X1 port map( C1 => n4911, C2 => n1987, A => n4894, B => n4893
                           , ZN => boothmul_pipelined_i_mux_out_2_12_port);
   U1962 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n4913, B1 => data1_mul_9_port, B2 => n4908, ZN
                           => n4896);
   U1963 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n4912, ZN => n4895);
   U1964 : OAI211_X1 port map( C1 => n4911, C2 => n1986, A => n4896, B => n4895
                           , ZN => boothmul_pipelined_i_mux_out_2_13_port);
   U1965 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n4913, B1 => data1_mul_10_port, B2 => n4905, 
                           ZN => n4898);
   U1966 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n4912, ZN => n4897);
   U1967 : OAI211_X1 port map( C1 => n4911, C2 => n1985, A => n4898, B => n4897
                           , ZN => boothmul_pipelined_i_mux_out_2_14_port);
   U1968 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n4913, B1 => data1_mul_11_port, B2 => n4905, 
                           ZN => n4900);
   U1969 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n4912, ZN => n4899);
   U1970 : OAI211_X1 port map( C1 => n4911, C2 => n1984, A => n4900, B => n4899
                           , ZN => boothmul_pipelined_i_mux_out_2_15_port);
   U1971 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n4913, B1 => data1_mul_12_port, B2 => n4908, 
                           ZN => n4902);
   U1972 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n4912, ZN => n4901);
   U1973 : OAI211_X1 port map( C1 => n4911, C2 => n1983, A => n4902, B => n4901
                           , ZN => boothmul_pipelined_i_mux_out_2_16_port);
   U1974 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n4913, B1 => data1_mul_13_port, B2 => n4905, 
                           ZN => n4904);
   U1975 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n4912, ZN => n4903);
   U1976 : OAI211_X1 port map( C1 => n4911, C2 => n1982, A => n4904, B => n4903
                           , ZN => boothmul_pipelined_i_mux_out_2_17_port);
   U1977 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n4913, B1 => data1_mul_14_port, B2 => n4905, 
                           ZN => n4907);
   U1978 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n4912, ZN => n4906);
   U1979 : OAI211_X1 port map( C1 => n4911, C2 => n1981, A => n4907, B => n4906
                           , ZN => boothmul_pipelined_i_mux_out_2_18_port);
   U1980 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n4913, B1 => data1_mul_15_port, B2 => n4908, 
                           ZN => n4910);
   U1981 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n4912, ZN => n4909);
   U1982 : OAI211_X1 port map( C1 => n4911, C2 => n1980, A => n4910, B => n4909
                           , ZN => boothmul_pipelined_i_mux_out_2_19_port);
   U1983 : NAND2_X1 port map( A1 => n3076, A2 => data1_mul_15_port, ZN => n4916
                           );
   U1984 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n4913, B1 => n4912, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n4914);
   U1985 : OAI21_X1 port map( B1 => n4916, B2 => n4915, A => n4914, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1986 : INV_X1 port map( A => n4949, ZN => n4918);
   U1987 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_176_port, ZN
                           => n4917);
   U1988 : OAI221_X1 port map( B1 => n3077, B2 => n4919, C1 => n3077, C2 => 
                           n4918, A => n4917, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1989 : CLKBUF_X1 port map( A => n4949, Z => n4945);
   U1990 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_3_60_port, A2
                           => n4950, B1 => n4945, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n4921);
   U1991 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n4920);
   U1992 : NAND2_X1 port map( A1 => n4921, A2 => n4920, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1993 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n4949
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n4923);
   U1994 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n4922);
   U1995 : NAND2_X1 port map( A1 => n4923, A2 => n4922, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1996 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n4949
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n4925);
   U1997 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n4924);
   U1998 : NAND2_X1 port map( A1 => n4925, A2 => n4924, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1999 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n4927);
   U2000 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n4926);
   U2001 : NAND2_X1 port map( A1 => n4927, A2 => n4926, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U2002 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n4929);
   U2003 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n4928);
   U2004 : NAND2_X1 port map( A1 => n4929, A2 => n4928, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U2005 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n4931);
   U2006 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n4930);
   U2007 : NAND2_X1 port map( A1 => n4931, A2 => n4930, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U2008 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n4934);
   U2009 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n4932
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n4933);
   U2010 : NAND2_X1 port map( A1 => n4934, A2 => n4933, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U2011 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n4936);
   U2012 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n4935);
   U2013 : NAND2_X1 port map( A1 => n4936, A2 => n4935, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U2014 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n4938);
   U2015 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n4937);
   U2016 : NAND2_X1 port map( A1 => n4938, A2 => n4937, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U2017 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n4940);
   U2018 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n4939);
   U2019 : NAND2_X1 port map( A1 => n4940, A2 => n4939, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U2020 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n4942);
   U2021 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n4941);
   U2022 : NAND2_X1 port map( A1 => n4942, A2 => n4941, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U2023 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n4949
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n4944);
   U2024 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n4943);
   U2025 : NAND2_X1 port map( A1 => n4944, A2 => n4943, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U2026 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n4945
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n4948);
   U2027 : AOI22_X1 port map( A1 => n4946, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n4947);
   U2028 : NAND2_X1 port map( A1 => n4948, A2 => n4947, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U2029 : AOI22_X1 port map( A1 => n4950, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n4949
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n4954);
   U2030 : AOI22_X1 port map( A1 => n4952, A2 => 
                           boothmul_pipelined_i_muxes_in_3_46_port, B1 => n4951
                           , B2 => boothmul_pipelined_i_muxes_in_3_162_port, ZN
                           => n4953);
   U2031 : NAND2_X1 port map( A1 => n4954, A2 => n4953, ZN => 
                           boothmul_pipelined_i_mux_out_3_21_port);
   U2032 : NAND3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n5109);
   U2033 : NOR3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n5107);
   U2034 : INV_X1 port map( A => n5107, ZN => n4958);
   U2035 : NAND2_X1 port map( A1 => n3078, A2 => n4955, ZN => n5110);
   U2036 : INV_X1 port map( A => n5110, ZN => n4988);
   U2037 : NOR2_X1 port map( A1 => n3078, A2 => n4956, ZN => n4971);
   U2038 : CLKBUF_X1 port map( A => n4971, Z => n5106);
   U2039 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_190_port, ZN
                           => n4957);
   U2040 : OAI221_X1 port map( B1 => n5121, B2 => n5109, C1 => n5121, C2 => 
                           n4958, A => n4957, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U2041 : INV_X1 port map( A => n5109, ZN => n4987);
   U2042 : CLKBUF_X1 port map( A => n5107, Z => n4984);
   U2043 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_64_port, A2
                           => n4987, B1 => n4984, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n4960);
   U2044 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n4959);
   U2045 : NAND2_X1 port map( A1 => n4960, A2 => n4959, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U2046 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n5107
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n4962);
   U2047 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n4961);
   U2048 : NAND2_X1 port map( A1 => n4962, A2 => n4961, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U2049 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n5107
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n4964);
   U2050 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n4963);
   U2051 : NAND2_X1 port map( A1 => n4964, A2 => n4963, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2052 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n4966);
   U2053 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n4965);
   U2054 : NAND2_X1 port map( A1 => n4966, A2 => n4965, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2055 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n4968);
   U2056 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n4967);
   U2057 : NAND2_X1 port map( A1 => n4968, A2 => n4967, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2058 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n4970);
   U2059 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n4969);
   U2060 : NAND2_X1 port map( A1 => n4970, A2 => n4969, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2061 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n4973);
   U2062 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n4971
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n4972);
   U2063 : NAND2_X1 port map( A1 => n4973, A2 => n4972, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2064 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n4975);
   U2065 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n4974);
   U2066 : NAND2_X1 port map( A1 => n4975, A2 => n4974, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2067 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n4977);
   U2068 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n4976);
   U2069 : NAND2_X1 port map( A1 => n4977, A2 => n4976, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2070 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n4979);
   U2071 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n4978);
   U2072 : NAND2_X1 port map( A1 => n4979, A2 => n4978, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2073 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n4981);
   U2074 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n4980);
   U2075 : NAND2_X1 port map( A1 => n4981, A2 => n4980, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2076 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n5107
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n4983);
   U2077 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n4982);
   U2078 : NAND2_X1 port map( A1 => n4983, A2 => n4982, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2079 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n4984
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n4986);
   U2080 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n4985);
   U2081 : NAND2_X1 port map( A1 => n4986, A2 => n4985, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2082 : AOI22_X1 port map( A1 => n4987, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n5107
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n4990);
   U2083 : AOI22_X1 port map( A1 => n4988, A2 => 
                           boothmul_pipelined_i_muxes_in_4_50_port, B1 => n5106
                           , B2 => boothmul_pipelined_i_muxes_in_4_176_port, ZN
                           => n4989);
   U2084 : NAND2_X1 port map( A1 => n4990, A2 => n4989, ZN => 
                           boothmul_pipelined_i_mux_out_4_23_port);
   U2085 : NAND3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n5114);
   U2086 : NOR3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n5112);
   U2087 : INV_X1 port map( A => n5112, ZN => n4994);
   U2088 : NAND2_X1 port map( A1 => n3079, A2 => n4991, ZN => n5115);
   U2089 : INV_X1 port map( A => n5115, ZN => n5024);
   U2090 : NOR2_X1 port map( A1 => n3079, A2 => n4992, ZN => n5007);
   U2091 : CLKBUF_X1 port map( A => n5007, Z => n5111);
   U2092 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_204_port, ZN
                           => n4993);
   U2093 : OAI221_X1 port map( B1 => n5122, B2 => n5114, C1 => n5122, C2 => 
                           n4994, A => n4993, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2094 : INV_X1 port map( A => n5114, ZN => n5023);
   U2095 : CLKBUF_X1 port map( A => n5112, Z => n5020);
   U2096 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_5_68_port, A2
                           => n5023, B1 => n5020, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n4996);
   U2097 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n4995);
   U2098 : NAND2_X1 port map( A1 => n4996, A2 => n4995, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2099 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n5112
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n4998);
   U2100 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n4997);
   U2101 : NAND2_X1 port map( A1 => n4998, A2 => n4997, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2102 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n5112
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n5000);
   U2103 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n4999);
   U2104 : NAND2_X1 port map( A1 => n5000, A2 => n4999, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2105 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n5002);
   U2106 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n5001);
   U2107 : NAND2_X1 port map( A1 => n5002, A2 => n5001, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2108 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n5004);
   U2109 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n5003);
   U2110 : NAND2_X1 port map( A1 => n5004, A2 => n5003, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2111 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n5006);
   U2112 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n5005);
   U2113 : NAND2_X1 port map( A1 => n5006, A2 => n5005, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2114 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n5009);
   U2115 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n5007
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n5008);
   U2116 : NAND2_X1 port map( A1 => n5009, A2 => n5008, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2117 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n5011);
   U2118 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n5010);
   U2119 : NAND2_X1 port map( A1 => n5011, A2 => n5010, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2120 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n5013);
   U2121 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n5012);
   U2122 : NAND2_X1 port map( A1 => n5013, A2 => n5012, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2123 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n5015);
   U2124 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n5014);
   U2125 : NAND2_X1 port map( A1 => n5015, A2 => n5014, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2126 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n5017);
   U2127 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n5016);
   U2128 : NAND2_X1 port map( A1 => n5017, A2 => n5016, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2129 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n5112
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n5019);
   U2130 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n5018);
   U2131 : NAND2_X1 port map( A1 => n5019, A2 => n5018, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2132 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n5020
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n5022);
   U2133 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n5021);
   U2134 : NAND2_X1 port map( A1 => n5022, A2 => n5021, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2135 : AOI22_X1 port map( A1 => n5023, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n5112
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n5026);
   U2136 : AOI22_X1 port map( A1 => n5024, A2 => 
                           boothmul_pipelined_i_muxes_in_5_54_port, B1 => n5111
                           , B2 => boothmul_pipelined_i_muxes_in_5_190_port, ZN
                           => n5025);
   U2137 : NAND2_X1 port map( A1 => n5026, A2 => n5025, ZN => 
                           boothmul_pipelined_i_mux_out_5_25_port);
   U2138 : NAND3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n5119);
   U2139 : NOR3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n5117);
   U2140 : INV_X1 port map( A => n5117, ZN => n5030);
   U2141 : NAND2_X1 port map( A1 => n3080, A2 => n5027, ZN => n5120);
   U2142 : INV_X1 port map( A => n5120, ZN => n5060);
   U2143 : NOR2_X1 port map( A1 => n3080, A2 => n5028, ZN => n5043);
   U2144 : CLKBUF_X1 port map( A => n5043, Z => n5116);
   U2145 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_218_port, ZN
                           => n5029);
   U2146 : OAI221_X1 port map( B1 => n5123, B2 => n5119, C1 => n5123, C2 => 
                           n5030, A => n5029, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2147 : INV_X1 port map( A => n5119, ZN => n5059);
   U2148 : CLKBUF_X1 port map( A => n5117, Z => n5056);
   U2149 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_6_72_port, A2
                           => n5059, B1 => n5056, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n5032);
   U2150 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n5031);
   U2151 : NAND2_X1 port map( A1 => n5032, A2 => n5031, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2152 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n5117
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n5034);
   U2153 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n5033);
   U2154 : NAND2_X1 port map( A1 => n5034, A2 => n5033, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2155 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n5117
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n5036);
   U2156 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n5035);
   U2157 : NAND2_X1 port map( A1 => n5036, A2 => n5035, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2158 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n5038);
   U2159 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n5037);
   U2160 : NAND2_X1 port map( A1 => n5038, A2 => n5037, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2161 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n5040);
   U2162 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n5039);
   U2163 : NAND2_X1 port map( A1 => n5040, A2 => n5039, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2164 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n5042);
   U2165 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n5041);
   U2166 : NAND2_X1 port map( A1 => n5042, A2 => n5041, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2167 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n5045);
   U2168 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n5043
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n5044);
   U2169 : NAND2_X1 port map( A1 => n5045, A2 => n5044, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2170 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n5047);
   U2171 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n5046);
   U2172 : NAND2_X1 port map( A1 => n5047, A2 => n5046, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2173 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n5049);
   U2174 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n5048);
   U2175 : NAND2_X1 port map( A1 => n5049, A2 => n5048, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2176 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n5051);
   U2177 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n5050);
   U2178 : NAND2_X1 port map( A1 => n5051, A2 => n5050, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2179 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n5053);
   U2180 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n5052);
   U2181 : NAND2_X1 port map( A1 => n5053, A2 => n5052, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2182 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n5117
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n5055);
   U2183 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n5054);
   U2184 : NAND2_X1 port map( A1 => n5055, A2 => n5054, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2185 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n5056
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n5058);
   U2186 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n5057);
   U2187 : NAND2_X1 port map( A1 => n5058, A2 => n5057, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2188 : AOI22_X1 port map( A1 => n5059, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n5117
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n5062);
   U2189 : AOI22_X1 port map( A1 => n5060, A2 => 
                           boothmul_pipelined_i_muxes_in_6_58_port, B1 => n5116
                           , B2 => boothmul_pipelined_i_muxes_in_6_204_port, ZN
                           => n5061);
   U2190 : NAND2_X1 port map( A1 => n5062, A2 => n5061, ZN => 
                           boothmul_pipelined_i_mux_out_6_27_port);
   U2191 : NAND3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A3 => n5125, ZN => n5066);
   U2192 : NAND2_X1 port map( A1 => n5063, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, ZN 
                           => n5067);
   U2193 : AND2_X1 port map( A1 => n5125, A2 => n5064, ZN => n5097);
   U2194 : AND2_X1 port map( A1 => n5064, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, ZN 
                           => n5098);
   U2195 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_76_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_232_port, ZN
                           => n5065);
   U2196 : OAI221_X1 port map( B1 => n5134, B2 => n5066, C1 => n5134, C2 => 
                           n5067, A => n5065, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2197 : INV_X1 port map( A => n5066, ZN => n5096);
   U2198 : INV_X1 port map( A => n5067, ZN => n5099);
   U2199 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_7_76_port, A2
                           => n5096, B1 => n5099, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n5069);
   U2200 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n5068);
   U2201 : NAND2_X1 port map( A1 => n5069, A2 => n5068, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2202 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n5071);
   U2203 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n5070);
   U2204 : NAND2_X1 port map( A1 => n5071, A2 => n5070, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2205 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n5073);
   U2206 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n5072);
   U2207 : NAND2_X1 port map( A1 => n5073, A2 => n5072, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2208 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n5075);
   U2209 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n5074);
   U2210 : NAND2_X1 port map( A1 => n5075, A2 => n5074, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2211 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n5077);
   U2212 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n5076);
   U2213 : NAND2_X1 port map( A1 => n5077, A2 => n5076, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2214 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n5079);
   U2215 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n5078);
   U2216 : NAND2_X1 port map( A1 => n5079, A2 => n5078, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2217 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n5081);
   U2218 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n5080);
   U2219 : NAND2_X1 port map( A1 => n5081, A2 => n5080, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2220 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n5083);
   U2221 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n5082);
   U2222 : NAND2_X1 port map( A1 => n5083, A2 => n5082, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2223 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n5085);
   U2224 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n5084);
   U2225 : NAND2_X1 port map( A1 => n5085, A2 => n5084, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2226 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n5087);
   U2227 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n5086);
   U2228 : NAND2_X1 port map( A1 => n5087, A2 => n5086, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2229 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n5089);
   U2230 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n5088);
   U2231 : NAND2_X1 port map( A1 => n5089, A2 => n5088, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2232 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n5091);
   U2233 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n5090);
   U2234 : NAND2_X1 port map( A1 => n5091, A2 => n5090, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2235 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n5093);
   U2236 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n5092);
   U2237 : NAND2_X1 port map( A1 => n5093, A2 => n5092, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2238 : AOI22_X1 port map( A1 => n5096, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n5099
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n5095);
   U2239 : AOI22_X1 port map( A1 => n5097, A2 => 
                           boothmul_pipelined_i_muxes_in_7_62_port, B1 => n5098
                           , B2 => boothmul_pipelined_i_muxes_in_7_218_port, ZN
                           => n5094);
   U2240 : NAND2_X1 port map( A1 => n5095, A2 => n5094, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2241 : OAI21_X1 port map( B1 => n5097, B2 => n5096, A => 
                           boothmul_pipelined_i_muxes_in_7_62_port, ZN => n5101
                           );
   U2242 : AOI22_X1 port map( A1 => n5099, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n5098, B2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, ZN => 
                           n5100);
   U2243 : NAND2_X1 port map( A1 => n5101, A2 => n5100, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2244 : AOI22_X1 port map( A1 => n5103, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n5102, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n5104);
   U2245 : OAI21_X1 port map( B1 => n5105, B2 => n1979, A => n5104, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2246 : AOI22_X1 port map( A1 => n5107, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, B1 => 
                           n5106, B2 => 
                           boothmul_pipelined_i_muxes_in_4_175_port, ZN => 
                           n5108);
   U2247 : OAI221_X1 port map( B1 => n5127, B2 => n5110, C1 => n5127, C2 => 
                           n5109, A => n5108, ZN => n1997);
   U2248 : AOI22_X1 port map( A1 => n5112, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, B1 => 
                           n5111, B2 => 
                           boothmul_pipelined_i_muxes_in_5_189_port, ZN => 
                           n5113);
   U2249 : OAI221_X1 port map( B1 => n5128, B2 => n5115, C1 => n5128, C2 => 
                           n5114, A => n5113, ZN => n1996);
   U2250 : AOI22_X1 port map( A1 => n5117, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, B1 => 
                           n5116, B2 => 
                           boothmul_pipelined_i_muxes_in_6_203_port, ZN => 
                           n5118);
   U2251 : OAI221_X1 port map( B1 => n5129, B2 => n5120, C1 => n5129, C2 => 
                           n5119, A => n5118, ZN => n1995);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
      n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, 
      n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
      n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
      n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, 
      n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, 
      n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
      n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, 
      n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
      n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, 
      n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
      n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, 
      n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, 
      n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
      n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, 
      n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, 
      n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, 
      n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
      n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, 
      n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, 
      n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, 
      n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, 
      n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
      n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, 
      n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, 
      n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, 
      n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, 
      n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
      n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, 
      n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
      n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
      n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
      n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
      n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, 
      n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, 
      n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, 
      n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
      n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
      n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
      n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, 
      n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
      n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
      n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, 
      n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
      n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
      n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
      n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
      n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, 
      n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
      n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
      n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
      n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, 
      n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, 
      n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
      n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, 
      n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, 
      n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, 
      n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, 
      n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
      n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, 
      n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
      n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
      n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, 
      n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, 
      n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
      n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
      n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
      n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, 
      n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, 
      n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, 
      n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, 
      n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, 
      n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, 
      n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, 
      n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, 
      n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, 
      n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, 
      n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, 
      n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, 
      n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, 
      n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, 
      n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, 
      n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, 
      n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, 
      n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, 
      n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, 
      n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, 
      n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, 
      n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, 
      n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, 
      n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, 
      n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, 
      n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, 
      n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, 
      n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, 
      n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, 
      n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, 
      n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, 
      n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, 
      n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, 
      n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, 
      n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, 
      n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, 
      n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, 
      n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, 
      n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, 
      n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, 
      n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, 
      n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, 
      n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, 
      n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, 
      n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, 
      n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, 
      n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, 
      n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, 
      n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, 
      n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, 
      n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, 
      n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, 
      n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, 
      n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, 
      n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, 
      n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, 
      n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, 
      n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, 
      n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, 
      n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, 
      n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, 
      n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, 
      n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, 
      n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, 
      n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, 
      n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, 
      n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, 
      n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, 
      n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, 
      n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, 
      n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, 
      n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, 
      n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, 
      n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, 
      n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, 
      n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, 
      n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, 
      n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, 
      n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, 
      n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, 
      n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, 
      n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, 
      n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, 
      n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, 
      n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, 
      n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, 
      n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, 
      n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, 
      n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, 
      n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, 
      n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, 
      n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, 
      n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, 
      n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, 
      n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, 
      n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, 
      n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, 
      n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, 
      n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, 
      n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, 
      n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, 
      n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, 
      n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, 
      n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, 
      n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, 
      n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, 
      n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, 
      n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, 
      n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, 
      n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, 
      n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, 
      n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, 
      n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, 
      n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, 
      n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, 
      n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, 
      n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, 
      n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, 
      n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, 
      n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, 
      n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, 
      n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, 
      n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, 
      n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, 
      n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, 
      n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, 
      n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, 
      n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, 
      n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, 
      n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, 
      n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, 
      n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, 
      n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, 
      n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, 
      n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, 
      n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, 
      n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, 
      n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, 
      n8442, n8443, n8444, n8445, n8446, n8447, n_1349, n_1350, n_1351, n_1352,
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412 : std_logic;

begin
   
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n7429);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n7430);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n8192);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n7692);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n7944);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n7431);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n7432);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n8193);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n7945);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n8194);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n7433);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n8195);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n7693);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n7946);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n7434);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n7694);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n8196);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n8197);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n7695);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n8198);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n8199);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n7435);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n8200);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n7947);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n7436);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n7948);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n7949);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n7437);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n7950);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n7951);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n8201);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n7696);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n7697);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n7438);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n7439);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n7698);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n7699);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n7440);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n7700);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n7441);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n7701);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n7702);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n7442);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n7443);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n7444);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n7445);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n7703);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n7446);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n7704);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n7447);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n7448);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n7449);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n7450);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n7705);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n7451);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n7706);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n7707);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n7708);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n7709);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n7710);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n7452);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n7711);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n7712);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n7713);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n7714);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n8202);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n7715);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n7952);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n7453);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n7716);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n7717);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n7454);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n7718);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n7455);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n8203);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n7719);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n7953);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n7456);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n7457);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n7458);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n7720);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n7721);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n7954);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n7722);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n7723);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n7459);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n7460);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n7461);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n7724);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n7462);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n7725);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n7726);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n7727);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n7463);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n7728);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n7729);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n7955);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n7730);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n7464);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n7465);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n7466);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n8204);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n7467);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n7468);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n8205);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n7469);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n7731);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n7956);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n7732);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n7957);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n7733);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n7734);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n7470);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n7958);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n7735);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n7736);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n7471);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n7737);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n7738);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n8206);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n7472);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n7473);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n7474);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n7475);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n7959);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n7476);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n7477);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n7960);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n7961);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n8207);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n7962);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n8208);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n8209);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n7963);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n7964);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n7965);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n7966);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n7967);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n7478);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n7479);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n7968);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n8210);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n7969);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n8211);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n7970);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n8212);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n7971);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n7972);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n8213);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n7973);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n8214);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n7974);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n8215);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n8216);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n7975);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n7976);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n8217);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n7739);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n7977);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n7978);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n8218);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n8219);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n7740);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n7979);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n7741);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n7742);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n7980);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n8220);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n7743);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n8221);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n7981);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n8222);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n8223);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n7744);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n7982);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n7983);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n8224);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n7745);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n8225);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n7480);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n7481);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n8226);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n7482);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n7746);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n7984);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n7985);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n8227);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n8228);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n7747);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n7986);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n7987);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n7988);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n7989);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n7990);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n8229);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n7991);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n8230);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n7992);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n8231);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n8232);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n7993);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n7994);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n8233);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n8234);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n7995);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n8235);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n8236);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n8237);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n7996);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n7997);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n7998);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n7999);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n8000);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n8001);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n8002);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n8238);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n8003);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n8239);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n8240);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n8241);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n8004);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n8242);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n8005);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n8243);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n7748);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n7483);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n8006);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n7749);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n8007);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n8244);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n8245);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n7750);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n7484);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n7751);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n8246);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n7485);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n7752);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n7753);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n8247);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n8008);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n7486);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n7487);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n7754);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n8248);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n8249);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n8250);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n8251);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n7488);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n8252);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n7755);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n7489);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n8009);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n7756);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n8253);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n7757);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n7490);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n8254);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n7758);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n8010);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n7759);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n7760);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n7761);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n8255);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n7762);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n8256);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n8257);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n8258);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n8011);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n7491);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n7763);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n8259);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n7492);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n7764);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n7765);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n7766);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n7493);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n8012);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n8260);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n8261);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n8013);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n7494);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n7767);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n7495);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n8262);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n8014);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n7768);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n7769);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n7770);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n7496);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n7497);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n7771);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n7772);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n7498);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n7773);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n7774);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n7499);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n7500);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n7775);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n7501);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n7776);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n7777);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n7502);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n7503);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n7778);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n7504);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n7779);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n7505);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n7780);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n7506);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n7507);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n7508);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n7509);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n7781);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n7510);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n7511);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n7782);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n7512);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n7513);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n7514);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n8263);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n7783);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n7515);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n7784);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n7516);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n7785);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n7517);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n8015);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n8016);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n7518);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n7519);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n7520);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n7786);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n8264);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n7787);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n7788);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n7521);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n7522);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n7789);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n8017);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n7790);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n7523);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n7791);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n7792);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n7793);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n8265);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n7524);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n7794);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n7795);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n8018);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n8019);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n8020);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n7796);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n7525);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n8021);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n7526);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n8266);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n7797);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n8267);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n7798);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n7527);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n8022);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n7528);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n7799);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n7800);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n7529);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n7530);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n7531);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n7801);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n7802);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n8268);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n7803);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n8269);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n7804);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n7532);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n7533);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n7805);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n7534);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n7806);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n7535);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n7536);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n7537);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n7807);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n7808);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n8023);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n8024);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n8270);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n8271);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n8025);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n8026);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n8272);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n8027);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n8273);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n8274);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n7538);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n8275);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n8276);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n8028);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n8277);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n8029);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n8030);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n8278);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n8031);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n8032);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n8033);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n8279);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n8034);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n8035);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n7539);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n8280);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n8036);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n8281);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n7540);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n8282);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n8283);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n8284);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n7541);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n8037);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n8285);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n8038);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n8039);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n8040);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n7542);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n7809);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n8041);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n7810);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n8286);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n7543);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n8042);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n8287);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n8043);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n8044);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n8045);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n8288);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n7544);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n8046);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n8289);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n7811);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n7812);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n8290);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n8291);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n8047);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n8048);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n8292);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n8293);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n7813);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n7545);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n8294);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n8049);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n8295);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n8050);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n8296);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n8051);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n8052);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n8053);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n8054);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n8297);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n8298);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n8055);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n8299);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n8056);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n8300);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n8301);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n8302);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n8303);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n8057);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n8058);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n8304);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n8059);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n8060);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n8305);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n8306);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n8061);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n8307);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n8308);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n8062);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n8063);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n8309);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n8310);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n8064);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n8311);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n7814);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n7815);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n7546);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n7816);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n8312);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n8065);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n7547);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n7817);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n7548);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n8313);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n8066);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n7549);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n7550);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n8067);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n7818);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n8314);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n8068);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n8069);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n7819);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n7551);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n8315);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n8070);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n7552);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n8316);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n7553);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n8317);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n8318);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n8071);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n7820);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n8072);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n7554);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n7940);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n8073);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n8319);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n8320);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n7555);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n7821);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n8074);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n7556);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n8321);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n8075);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n8322);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n7822);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n8323);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n8324);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n7557);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n7823);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n7824);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n7825);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n8325);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n8326);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n7826);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n7827);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n7558);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n8076);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n7828);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n7829);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n7559);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n7830);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n7831);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n7560);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n8077);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n7561);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n7684);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n7832);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n7833);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n7562);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n8078);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n8079);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n7563);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n8327);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n7564);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n7565);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n7566);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n7567);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n7568);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n7569);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n7570);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n7834);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n7835);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n8328);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n7571);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n7836);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n7572);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n7573);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n8329);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n7574);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n8080);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n7837);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n7575);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n8081);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n7576);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n7577);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n7578);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n7838);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n7685);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n8330);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n8331);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n7839);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n8082);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n7579);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n7840);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n8332);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n7580);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n7581);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n8083);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n7582);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n7841);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n7583);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n8084);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n8085);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n8086);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n8333);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n8087);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n8334);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n8335);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n8336);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n8337);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n8088);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n7842);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n8089);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n8090);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n7584);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n8091);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n7843);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n8338);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n7844);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n7424);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n7585);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n7845);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n7846);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n8339);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n7847);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n8340);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n8341);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n8342);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n7848);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n8092);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n8093);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n7586);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n8343);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n8094);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n8095);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n7587);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n8096);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n8344);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n7588);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n7589);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n7590);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n7849);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n8345);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n7591);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n7592);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n7593);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n8346);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n8347);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n8348);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n8097);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n8349);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n7686);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n8098);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n8099);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n7594);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n7850);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n8350);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n8351);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n8100);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n8101);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n8102);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n8103);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n8104);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n8352);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n8105);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n8353);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n8354);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n8106);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n8355);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n8356);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n8107);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n8108);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n8357);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n8109);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n8358);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n8110);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n8359);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n8360);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n8361);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n8362);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n8111);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n8363);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n8364);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n7941);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n8112);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n8113);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n8365);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n8114);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n8115);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n8366);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n8116);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n8117);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n8118);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n7851);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n8367);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n8119);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n8368);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n8369);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n8370);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n8120);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n8371);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n8372);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n8121);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n8373);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n8122);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n8374);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n8375);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n8376);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n8377);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n8378);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n8123);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n8379);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n8124);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n8380);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n8125);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n7942);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n8381);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n8382);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n8126);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n8383);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n8127);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n8384);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n8128);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n8129);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n8385);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n8386);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n8387);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n8388);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n8130);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n8389);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n8131);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n8132);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n8390);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n8133);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n8134);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n8135);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n8136);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n8137);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n8138);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n8391);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n8392);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n8393);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n8394);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n8139);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n8395);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n8140);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n8141);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n7687);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n7852);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n7853);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n8142);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n7595);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n7596);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n7597);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n7854);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n7855);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n8396);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n7856);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n7598);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n7599);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n7600);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n7857);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n7858);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n7859);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n7860);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n7861);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n7601);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n7862);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n8143);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n8144);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n7602);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n7603);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n7863);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n7864);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n7604);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n7605);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n7606);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n7865);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n7607);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n7425);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n8397);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n8145);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n8398);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n8399);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n8146);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n8400);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n7608);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n8147);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n8401);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n8402);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n8403);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n8404);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n8405);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n7866);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n7867);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n8406);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n8407);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n8148);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n8408);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n8149);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n8409);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n7609);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n8410);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n8411);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n8150);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n8151);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n7868);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n7610);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n8412);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n7869);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n7870);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n7688);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n7611);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n8152);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n7871);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n7612);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n7872);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n7873);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n7613);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n7874);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n7875);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n7876);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n7877);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n7614);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n7878);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n8413);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n7615);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n7616);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n7617);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n7879);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n7880);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n7618);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n7881);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n7882);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n7619);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n7620);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n8414);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n8415);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n7621);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n7622);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n7623);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n7624);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n7625);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n7689);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n8416);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n8153);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n8154);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n8417);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n8418);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n8155);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n7883);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n7884);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n8419);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n7885);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n7886);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n8156);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n8157);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n7626);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n7887);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n8420);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n7627);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n8421);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n8422);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n7628);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n8423);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n7888);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n7629);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n8158);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n8159);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n8424);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n8160);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n7889);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n8425);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n8426);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n8161);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n7426);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n7630);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n7631);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n7890);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n8162);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n7632);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n8163);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n7891);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n8164);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n7633);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n8165);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n7634);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n7892);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n7635);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n7636);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n7637);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n7893);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n7638);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n7639);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n7640);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n8427);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n7641);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n7894);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n7895);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n7642);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n7643);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n7896);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n7897);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n8428);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n7898);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n7644);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n8429);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n7690);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n7645);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n7899);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n8166);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n7646);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n8430);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n7647);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n8167);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n7900);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n7901);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n7902);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n8431);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n8432);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n8433);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n8168);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n8169);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n7648);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n7649);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n7650);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n7651);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n7652);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n7903);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n8170);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n8434);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n8171);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n7904);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n7905);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n8435);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n8436);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n8172);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n7906);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n8173);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n7691);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n7907);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n7653);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n7654);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n7908);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n7909);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n7655);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n7910);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n7656);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n7657);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n7658);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n8174);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n7911);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n7912);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n7913);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n8437);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n8438);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n7659);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n7914);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n7915);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n8439);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n7660);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n7661);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n7916);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n7917);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n7662);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n8175);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n7663);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n7918);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n7919);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n7664);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n7665);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n7427);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n7666);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n7667);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n7920);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n7921);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n7668);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n7669);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n7922);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n7923);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n7924);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n7670);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n7925);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n7671);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n7672);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n7673);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n7674);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n7926);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n7675);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n7676);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n7927);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n7928);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n7929);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n7930);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n7677);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n7931);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n7678);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n7679);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n7932);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n7680);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n7681);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n7933);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n7934);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n7943);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n8440);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n7935);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n8176);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n7936);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n8441);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n7937);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n8177);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n8442);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n8178);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n8179);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n8180);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n8181);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n7938);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n8443);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n8182);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n8183);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n8184);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n7682);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n8185);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n8444);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n8186);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n8187);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n7939);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n8445);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n8188);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n7683);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n8189);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n8190);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n8446);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n8191);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n8447);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1349);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1350);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1351);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1352);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1353);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1354);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1355);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1356);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1357);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1358);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1359);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1360);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1361);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1362);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1363);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1364);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1365);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1366);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1367);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1368);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1369);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1370);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1371);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1372);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1373);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1374);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1375);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1376);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1377);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1378);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1379);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1380);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1381);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1382);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1383);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1384);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1385);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1386);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1387);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1388);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1389);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1390);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1391);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1392);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1393);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1394);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1395);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1396);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1397);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1398);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1399);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1400);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1401);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1402);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1403);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1404);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1405);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1406);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1407);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1408);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1409);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1410);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1411);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1412);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n7428);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n5672);
   U4 : CLKBUF_X1 port map( A => RESET_BAR, Z => n5673);
   U5 : CLKBUF_X1 port map( A => RESET_BAR, Z => n5674);
   U6 : CLKBUF_X1 port map( A => RESET_BAR, Z => n5675);
   U7 : NAND2_X2 port map( A1 => n5672, A2 => n5730, ZN => n5732);
   U8 : NAND2_X2 port map( A1 => n5675, A2 => n5726, ZN => n5728);
   U9 : NAND2_X2 port map( A1 => n5675, A2 => n5723, ZN => n5725);
   U10 : NAND2_X2 port map( A1 => n5672, A2 => n5720, ZN => n5722);
   U11 : NAND2_X2 port map( A1 => n5675, A2 => n5717, ZN => n5719);
   U12 : NAND2_X2 port map( A1 => n5672, A2 => n5714, ZN => n5716);
   U13 : NAND2_X2 port map( A1 => n5675, A2 => n5711, ZN => n5713);
   U14 : NAND2_X2 port map( A1 => n5675, A2 => n5708, ZN => n5710);
   U15 : NAND2_X2 port map( A1 => n5672, A2 => n5847, ZN => n5859);
   U16 : NAND2_X2 port map( A1 => n5675, A2 => n5820, ZN => n5822);
   U17 : NAND2_X2 port map( A1 => n5672, A2 => n5816, ZN => n5818);
   U18 : NAND2_X2 port map( A1 => n5675, A2 => n5812, ZN => n5814);
   U19 : NAND2_X2 port map( A1 => n5674, A2 => n5808, ZN => n5810);
   U20 : NAND2_X2 port map( A1 => n5672, A2 => n5799, ZN => n5801);
   U21 : NAND2_X2 port map( A1 => n5672, A2 => n5795, ZN => n5797);
   U22 : NAND2_X2 port map( A1 => n5673, A2 => n5789, ZN => n5791);
   U23 : NAND2_X2 port map( A1 => n5673, A2 => n5780, ZN => n5782);
   U24 : NAND2_X2 port map( A1 => n5673, A2 => n5777, ZN => n5779);
   U25 : NAND2_X2 port map( A1 => n5673, A2 => n5774, ZN => n5776);
   U26 : NAND2_X2 port map( A1 => n5672, A2 => n5761, ZN => n5773);
   U27 : NAND2_X2 port map( A1 => n5672, A2 => n5737, ZN => n5739);
   U28 : NAND2_X2 port map( A1 => n5672, A2 => n5734, ZN => n5736);
   U29 : NAND2_X2 port map( A1 => n5672, A2 => n5705, ZN => n5707);
   U30 : NAND2_X2 port map( A1 => n5672, A2 => n5699, ZN => n5701);
   U31 : NAND2_X2 port map( A1 => n5672, A2 => n5695, ZN => n5697);
   U32 : NAND2_X2 port map( A1 => n5673, A2 => n5691, ZN => n5693);
   U33 : INV_X1 port map( A => ADD_WR(4), ZN => n5793);
   U34 : INV_X1 port map( A => ADD_WR(2), ZN => n5703);
   U35 : NOR2_X1 port map( A1 => n5793, A2 => n5792, ZN => n5823);
   U36 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n5694, ZN =>
                           n5798);
   U37 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n5733, ZN => n5704);
   U38 : CLKBUF_X1 port map( A => n6641, Z => n6586);
   U39 : CLKBUF_X1 port map( A => n7423, Z => n7367);
   U40 : CLKBUF_X1 port map( A => n5820, Z => n5821);
   U41 : NAND2_X1 port map( A1 => n5673, A2 => n5803, ZN => n5806);
   U42 : NAND2_X1 port map( A1 => n5673, A2 => n5783, ZN => n5786);
   U43 : CLKBUF_X1 port map( A => n5730, Z => n5731);
   U44 : CLKBUF_X1 port map( A => n5770, Z => n5856);
   U45 : CLKBUF_X1 port map( A => n5754, Z => n5840);
   U46 : CLKBUF_X1 port map( A => n5740, Z => n5826);
   U47 : CLKBUF_X1 port map( A => n5691, Z => n5692);
   U48 : NAND2_X1 port map( A1 => n5675, A2 => n5681, ZN => n5684);
   U49 : CLKBUF_X1 port map( A => n5680, Z => n5677);
   U50 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n5794);
   U51 : INV_X1 port map( A => ADD_WR(3), ZN => n5676);
   U52 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n5676, ZN => n5733);
   U53 : NAND2_X1 port map( A1 => n5794, A2 => n5704, ZN => n5678);
   U54 : CLKBUF_X1 port map( A => n5678, Z => n5679);
   U55 : NAND2_X1 port map( A1 => n5675, A2 => n5679, ZN => n5680);
   U56 : NAND2_X1 port map( A1 => n5675, A2 => DATAIN(31), ZN => n5825);
   U57 : CLKBUF_X1 port map( A => n5825, Z => n5788);
   U58 : OAI22_X1 port map( A1 => n7428, A2 => n5677, B1 => n5788, B2 => n5679,
                           ZN => n2166);
   U59 : NAND2_X1 port map( A1 => n5675, A2 => DATAIN(30), ZN => n5740);
   U60 : OAI22_X1 port map( A1 => n7429, A2 => n5680, B1 => n5679, B2 => n5740,
                           ZN => n2165);
   U61 : NAND2_X1 port map( A1 => n5675, A2 => DATAIN(29), ZN => n5741);
   U62 : OAI22_X1 port map( A1 => n7430, A2 => n5677, B1 => n5679, B2 => n5741,
                           ZN => n2164);
   U63 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(28), ZN => n5742);
   U64 : OAI22_X1 port map( A1 => n8192, A2 => n5680, B1 => n5679, B2 => n5742,
                           ZN => n2163);
   U65 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(27), ZN => n5743);
   U66 : OAI22_X1 port map( A1 => n7692, A2 => n5677, B1 => n5679, B2 => n5743,
                           ZN => n2162);
   U67 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(26), ZN => n5744);
   U68 : OAI22_X1 port map( A1 => n7944, A2 => n5680, B1 => n5679, B2 => n5744,
                           ZN => n2161);
   U69 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(25), ZN => n5745);
   U70 : OAI22_X1 port map( A1 => n7431, A2 => n5677, B1 => n5679, B2 => n5745,
                           ZN => n2160);
   U71 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(24), ZN => n5746);
   U72 : OAI22_X1 port map( A1 => n7432, A2 => n5680, B1 => n5679, B2 => n5746,
                           ZN => n2159);
   U73 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(23), ZN => n5747);
   U74 : OAI22_X1 port map( A1 => n8193, A2 => n5677, B1 => n5678, B2 => n5747,
                           ZN => n2158);
   U75 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(22), ZN => n5748);
   U76 : OAI22_X1 port map( A1 => n7945, A2 => n5680, B1 => n5678, B2 => n5748,
                           ZN => n2157);
   U77 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(21), ZN => n5749);
   U78 : OAI22_X1 port map( A1 => n8194, A2 => n5680, B1 => n5678, B2 => n5749,
                           ZN => n2156);
   U79 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(20), ZN => n5750);
   U80 : OAI22_X1 port map( A1 => n7433, A2 => n5680, B1 => n5678, B2 => n5750,
                           ZN => n2155);
   U81 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(19), ZN => n5751);
   U82 : OAI22_X1 port map( A1 => n8195, A2 => n5677, B1 => n5678, B2 => n5751,
                           ZN => n2154);
   U83 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(18), ZN => n5752);
   U84 : OAI22_X1 port map( A1 => n7693, A2 => n5677, B1 => n5678, B2 => n5752,
                           ZN => n2153);
   U85 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(17), ZN => n5753);
   U86 : OAI22_X1 port map( A1 => n7946, A2 => n5677, B1 => n5678, B2 => n5753,
                           ZN => n2152);
   U87 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(16), ZN => n5754);
   U88 : OAI22_X1 port map( A1 => n7434, A2 => n5677, B1 => n5678, B2 => n5754,
                           ZN => n2151);
   U89 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(15), ZN => n5755);
   U90 : OAI22_X1 port map( A1 => n7694, A2 => n5677, B1 => n5679, B2 => n5755,
                           ZN => n2150);
   U91 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(14), ZN => n5756);
   U92 : OAI22_X1 port map( A1 => n8196, A2 => n5677, B1 => n5678, B2 => n5756,
                           ZN => n2149);
   U93 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(13), ZN => n5757);
   U94 : OAI22_X1 port map( A1 => n8197, A2 => n5677, B1 => n5679, B2 => n5757,
                           ZN => n2148);
   U95 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(12), ZN => n5758);
   U96 : OAI22_X1 port map( A1 => n7695, A2 => n5677, B1 => n5678, B2 => n5758,
                           ZN => n2147);
   U97 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(11), ZN => n5759);
   U98 : OAI22_X1 port map( A1 => n8198, A2 => n5677, B1 => n5678, B2 => n5759,
                           ZN => n2146);
   U99 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(10), ZN => n5760);
   U100 : OAI22_X1 port map( A1 => n8199, A2 => n5677, B1 => n5678, B2 => n5760
                           , ZN => n2145);
   U101 : NAND2_X1 port map( A1 => n5674, A2 => DATAIN(9), ZN => n5762);
   U102 : OAI22_X1 port map( A1 => n7435, A2 => n5677, B1 => n5679, B2 => n5762
                           , ZN => n2144);
   U103 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(8), ZN => n5763);
   U104 : OAI22_X1 port map( A1 => n8200, A2 => n5677, B1 => n5678, B2 => n5763
                           , ZN => n2143);
   U105 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(7), ZN => n5764);
   U106 : OAI22_X1 port map( A1 => n7947, A2 => n5680, B1 => n5679, B2 => n5764
                           , ZN => n2142);
   U107 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(6), ZN => n5765);
   U108 : OAI22_X1 port map( A1 => n7436, A2 => n5680, B1 => n5678, B2 => n5765
                           , ZN => n2141);
   U109 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(5), ZN => n5766);
   U110 : OAI22_X1 port map( A1 => n7948, A2 => n5680, B1 => n5679, B2 => n5766
                           , ZN => n2140);
   U111 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(4), ZN => n5767);
   U112 : OAI22_X1 port map( A1 => n7949, A2 => n5680, B1 => n5678, B2 => n5767
                           , ZN => n2139);
   U113 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(3), ZN => n5768);
   U114 : OAI22_X1 port map( A1 => n7437, A2 => n5680, B1 => n5679, B2 => n5768
                           , ZN => n2138);
   U115 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(2), ZN => n5769);
   U116 : OAI22_X1 port map( A1 => n7950, A2 => n5680, B1 => n5678, B2 => n5769
                           , ZN => n2137);
   U117 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(1), ZN => n5770);
   U118 : OAI22_X1 port map( A1 => n7951, A2 => n5680, B1 => n5679, B2 => n5770
                           , ZN => n2136);
   U119 : NAND2_X1 port map( A1 => n5673, A2 => DATAIN(0), ZN => n5772);
   U120 : OAI22_X1 port map( A1 => n8201, A2 => n5680, B1 => n5679, B2 => n5772
                           , ZN => n2135);
   U121 : INV_X1 port map( A => ADD_WR(0), ZN => n5694);
   U122 : NAND2_X1 port map( A1 => n5704, A2 => n5798, ZN => n5681);
   U123 : CLKBUF_X1 port map( A => n5684, Z => n5682);
   U124 : CLKBUF_X1 port map( A => n5681, Z => n5683);
   U125 : OAI22_X1 port map( A1 => n7696, A2 => n5682, B1 => n5825, B2 => n5683
                           , ZN => n2134);
   U126 : OAI22_X1 port map( A1 => n7697, A2 => n5684, B1 => n5740, B2 => n5681
                           , ZN => n2133);
   U127 : OAI22_X1 port map( A1 => n7438, A2 => n5682, B1 => n5741, B2 => n5683
                           , ZN => n2132);
   U128 : OAI22_X1 port map( A1 => n7439, A2 => n5684, B1 => n5742, B2 => n5681
                           , ZN => n2131);
   U129 : OAI22_X1 port map( A1 => n7698, A2 => n5682, B1 => n5743, B2 => n5683
                           , ZN => n2130);
   U130 : OAI22_X1 port map( A1 => n7699, A2 => n5684, B1 => n5744, B2 => n5681
                           , ZN => n2129);
   U131 : OAI22_X1 port map( A1 => n7440, A2 => n5682, B1 => n5745, B2 => n5683
                           , ZN => n2128);
   U132 : OAI22_X1 port map( A1 => n7700, A2 => n5684, B1 => n5746, B2 => n5681
                           , ZN => n2127);
   U133 : OAI22_X1 port map( A1 => n7441, A2 => n5682, B1 => n5747, B2 => n5683
                           , ZN => n2126);
   U134 : OAI22_X1 port map( A1 => n7701, A2 => n5684, B1 => n5748, B2 => n5681
                           , ZN => n2125);
   U135 : OAI22_X1 port map( A1 => n7702, A2 => n5684, B1 => n5749, B2 => n5681
                           , ZN => n2124);
   U136 : OAI22_X1 port map( A1 => n7442, A2 => n5684, B1 => n5750, B2 => n5683
                           , ZN => n2123);
   U137 : OAI22_X1 port map( A1 => n7443, A2 => n5682, B1 => n5751, B2 => n5681
                           , ZN => n2122);
   U138 : OAI22_X1 port map( A1 => n7444, A2 => n5682, B1 => n5752, B2 => n5683
                           , ZN => n2121);
   U139 : OAI22_X1 port map( A1 => n7445, A2 => n5682, B1 => n5753, B2 => n5681
                           , ZN => n2120);
   U140 : OAI22_X1 port map( A1 => n7703, A2 => n5682, B1 => n5754, B2 => n5683
                           , ZN => n2119);
   U141 : OAI22_X1 port map( A1 => n7446, A2 => n5682, B1 => n5755, B2 => n5681
                           , ZN => n2118);
   U142 : OAI22_X1 port map( A1 => n7704, A2 => n5682, B1 => n5756, B2 => n5681
                           , ZN => n2117);
   U143 : OAI22_X1 port map( A1 => n7447, A2 => n5682, B1 => n5757, B2 => n5681
                           , ZN => n2116);
   U144 : OAI22_X1 port map( A1 => n7448, A2 => n5682, B1 => n5758, B2 => n5681
                           , ZN => n2115);
   U145 : OAI22_X1 port map( A1 => n7449, A2 => n5682, B1 => n5759, B2 => n5681
                           , ZN => n2114);
   U146 : OAI22_X1 port map( A1 => n7450, A2 => n5682, B1 => n5760, B2 => n5681
                           , ZN => n2113);
   U147 : OAI22_X1 port map( A1 => n7705, A2 => n5682, B1 => n5762, B2 => n5681
                           , ZN => n2112);
   U148 : OAI22_X1 port map( A1 => n7451, A2 => n5682, B1 => n5763, B2 => n5683
                           , ZN => n2111);
   U149 : OAI22_X1 port map( A1 => n7706, A2 => n5684, B1 => n5764, B2 => n5683
                           , ZN => n2110);
   U150 : OAI22_X1 port map( A1 => n7707, A2 => n5684, B1 => n5765, B2 => n5683
                           , ZN => n2109);
   U151 : OAI22_X1 port map( A1 => n7708, A2 => n5684, B1 => n5766, B2 => n5683
                           , ZN => n2108);
   U152 : OAI22_X1 port map( A1 => n7709, A2 => n5684, B1 => n5767, B2 => n5683
                           , ZN => n2107);
   U153 : OAI22_X1 port map( A1 => n7710, A2 => n5684, B1 => n5768, B2 => n5683
                           , ZN => n2106);
   U154 : OAI22_X1 port map( A1 => n7452, A2 => n5684, B1 => n5769, B2 => n5683
                           , ZN => n2105);
   U155 : OAI22_X1 port map( A1 => n7711, A2 => n5684, B1 => n5770, B2 => n5683
                           , ZN => n2104);
   U156 : OAI22_X1 port map( A1 => n7712, A2 => n5684, B1 => n5772, B2 => n5683
                           , ZN => n2103);
   U157 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n5694, ZN => n5698);
   U158 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n5698, ZN => n5802);
   U159 : NAND2_X1 port map( A1 => n5704, A2 => n5802, ZN => n5685);
   U160 : NAND2_X2 port map( A1 => n5675, A2 => n5685, ZN => n5687);
   U161 : CLKBUF_X1 port map( A => n5685, Z => n5686);
   U162 : OAI22_X1 port map( A1 => n7713, A2 => n5687, B1 => n5788, B2 => n5686
                           , ZN => n2102);
   U163 : OAI22_X1 port map( A1 => n7714, A2 => n5687, B1 => n5740, B2 => n5685
                           , ZN => n2101);
   U164 : OAI22_X1 port map( A1 => n8202, A2 => n5687, B1 => n5741, B2 => n5686
                           , ZN => n2100);
   U165 : OAI22_X1 port map( A1 => n7715, A2 => n5687, B1 => n5742, B2 => n5685
                           , ZN => n2099);
   U166 : OAI22_X1 port map( A1 => n7952, A2 => n5687, B1 => n5743, B2 => n5686
                           , ZN => n2098);
   U167 : OAI22_X1 port map( A1 => n7453, A2 => n5687, B1 => n5744, B2 => n5685
                           , ZN => n2097);
   U168 : OAI22_X1 port map( A1 => n7716, A2 => n5687, B1 => n5745, B2 => n5686
                           , ZN => n2096);
   U169 : OAI22_X1 port map( A1 => n7717, A2 => n5687, B1 => n5746, B2 => n5685
                           , ZN => n2095);
   U170 : OAI22_X1 port map( A1 => n7454, A2 => n5687, B1 => n5747, B2 => n5686
                           , ZN => n2094);
   U171 : OAI22_X1 port map( A1 => n7718, A2 => n5687, B1 => n5748, B2 => n5685
                           , ZN => n2093);
   U172 : OAI22_X1 port map( A1 => n7455, A2 => n5687, B1 => n5749, B2 => n5685
                           , ZN => n2092);
   U173 : OAI22_X1 port map( A1 => n8203, A2 => n5687, B1 => n5750, B2 => n5686
                           , ZN => n2091);
   U174 : OAI22_X1 port map( A1 => n7719, A2 => n5687, B1 => n5751, B2 => n5685
                           , ZN => n2090);
   U175 : OAI22_X1 port map( A1 => n7953, A2 => n5687, B1 => n5752, B2 => n5686
                           , ZN => n2089);
   U176 : OAI22_X1 port map( A1 => n7456, A2 => n5687, B1 => n5753, B2 => n5685
                           , ZN => n2088);
   U177 : OAI22_X1 port map( A1 => n7457, A2 => n5687, B1 => n5754, B2 => n5686
                           , ZN => n2087);
   U178 : OAI22_X1 port map( A1 => n7458, A2 => n5687, B1 => n5755, B2 => n5685
                           , ZN => n2086);
   U179 : OAI22_X1 port map( A1 => n7720, A2 => n5687, B1 => n5756, B2 => n5685
                           , ZN => n2085);
   U180 : OAI22_X1 port map( A1 => n7721, A2 => n5687, B1 => n5757, B2 => n5685
                           , ZN => n2084);
   U181 : OAI22_X1 port map( A1 => n7954, A2 => n5687, B1 => n5758, B2 => n5685
                           , ZN => n2083);
   U182 : OAI22_X1 port map( A1 => n7722, A2 => n5687, B1 => n5759, B2 => n5685
                           , ZN => n2082);
   U183 : OAI22_X1 port map( A1 => n7723, A2 => n5687, B1 => n5760, B2 => n5685
                           , ZN => n2081);
   U184 : OAI22_X1 port map( A1 => n7459, A2 => n5687, B1 => n5762, B2 => n5685
                           , ZN => n2080);
   U185 : OAI22_X1 port map( A1 => n7460, A2 => n5687, B1 => n5763, B2 => n5686
                           , ZN => n2079);
   U186 : OAI22_X1 port map( A1 => n7461, A2 => n5687, B1 => n5764, B2 => n5686
                           , ZN => n2078);
   U187 : OAI22_X1 port map( A1 => n7724, A2 => n5687, B1 => n5765, B2 => n5686
                           , ZN => n2077);
   U188 : OAI22_X1 port map( A1 => n7462, A2 => n5687, B1 => n5766, B2 => n5686
                           , ZN => n2076);
   U189 : OAI22_X1 port map( A1 => n7725, A2 => n5687, B1 => n5767, B2 => n5686
                           , ZN => n2075);
   U190 : OAI22_X1 port map( A1 => n7726, A2 => n5687, B1 => n5768, B2 => n5686
                           , ZN => n2074);
   U191 : OAI22_X1 port map( A1 => n7727, A2 => n5687, B1 => n5769, B2 => n5686
                           , ZN => n2073);
   U192 : OAI22_X1 port map( A1 => n7463, A2 => n5687, B1 => n5770, B2 => n5686
                           , ZN => n2072);
   U193 : OAI22_X1 port map( A1 => n7728, A2 => n5687, B1 => n5772, B2 => n5686
                           , ZN => n2071);
   U194 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n5702);
   U195 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n5702, ZN => n5807);
   U196 : NAND2_X1 port map( A1 => n5704, A2 => n5807, ZN => n5688);
   U197 : NAND2_X2 port map( A1 => n5675, A2 => n5688, ZN => n5690);
   U198 : CLKBUF_X1 port map( A => n5688, Z => n5689);
   U199 : OAI22_X1 port map( A1 => n7729, A2 => n5690, B1 => n5825, B2 => n5689
                           , ZN => n2070);
   U200 : OAI22_X1 port map( A1 => n7955, A2 => n5690, B1 => n5740, B2 => n5688
                           , ZN => n2069);
   U201 : OAI22_X1 port map( A1 => n7730, A2 => n5690, B1 => n5741, B2 => n5689
                           , ZN => n2068);
   U202 : OAI22_X1 port map( A1 => n7464, A2 => n5690, B1 => n5742, B2 => n5688
                           , ZN => n2067);
   U203 : OAI22_X1 port map( A1 => n7465, A2 => n5690, B1 => n5743, B2 => n5689
                           , ZN => n2066);
   U204 : OAI22_X1 port map( A1 => n7466, A2 => n5690, B1 => n5744, B2 => n5688
                           , ZN => n2065);
   U205 : OAI22_X1 port map( A1 => n8204, A2 => n5690, B1 => n5745, B2 => n5689
                           , ZN => n2064);
   U206 : OAI22_X1 port map( A1 => n7467, A2 => n5690, B1 => n5746, B2 => n5688
                           , ZN => n2063);
   U207 : OAI22_X1 port map( A1 => n7468, A2 => n5690, B1 => n5747, B2 => n5689
                           , ZN => n2062);
   U208 : OAI22_X1 port map( A1 => n8205, A2 => n5690, B1 => n5748, B2 => n5688
                           , ZN => n2061);
   U209 : OAI22_X1 port map( A1 => n7469, A2 => n5690, B1 => n5749, B2 => n5688
                           , ZN => n2060);
   U210 : OAI22_X1 port map( A1 => n7731, A2 => n5690, B1 => n5750, B2 => n5689
                           , ZN => n2059);
   U211 : OAI22_X1 port map( A1 => n7956, A2 => n5690, B1 => n5751, B2 => n5688
                           , ZN => n2058);
   U212 : OAI22_X1 port map( A1 => n7732, A2 => n5690, B1 => n5752, B2 => n5689
                           , ZN => n2057);
   U213 : OAI22_X1 port map( A1 => n7957, A2 => n5690, B1 => n5753, B2 => n5688
                           , ZN => n2056);
   U214 : OAI22_X1 port map( A1 => n7733, A2 => n5690, B1 => n5754, B2 => n5689
                           , ZN => n2055);
   U215 : OAI22_X1 port map( A1 => n7734, A2 => n5690, B1 => n5755, B2 => n5688
                           , ZN => n2054);
   U216 : OAI22_X1 port map( A1 => n7470, A2 => n5690, B1 => n5756, B2 => n5688
                           , ZN => n2053);
   U217 : OAI22_X1 port map( A1 => n7958, A2 => n5690, B1 => n5757, B2 => n5688
                           , ZN => n2052);
   U218 : OAI22_X1 port map( A1 => n7735, A2 => n5690, B1 => n5758, B2 => n5688
                           , ZN => n2051);
   U219 : OAI22_X1 port map( A1 => n7736, A2 => n5690, B1 => n5759, B2 => n5688
                           , ZN => n2050);
   U220 : OAI22_X1 port map( A1 => n7471, A2 => n5690, B1 => n5760, B2 => n5688
                           , ZN => n2049);
   U221 : OAI22_X1 port map( A1 => n7737, A2 => n5690, B1 => n5762, B2 => n5688
                           , ZN => n2048);
   U222 : OAI22_X1 port map( A1 => n7738, A2 => n5690, B1 => n5763, B2 => n5689
                           , ZN => n2047);
   U223 : OAI22_X1 port map( A1 => n8206, A2 => n5690, B1 => n5764, B2 => n5689
                           , ZN => n2046);
   U224 : OAI22_X1 port map( A1 => n7472, A2 => n5690, B1 => n5765, B2 => n5689
                           , ZN => n2045);
   U225 : OAI22_X1 port map( A1 => n7473, A2 => n5690, B1 => n5766, B2 => n5689
                           , ZN => n2044);
   U226 : OAI22_X1 port map( A1 => n7474, A2 => n5690, B1 => n5767, B2 => n5689
                           , ZN => n2043);
   U227 : OAI22_X1 port map( A1 => n7475, A2 => n5690, B1 => n5768, B2 => n5689
                           , ZN => n2042);
   U228 : OAI22_X1 port map( A1 => n7959, A2 => n5690, B1 => n5769, B2 => n5689
                           , ZN => n2041);
   U229 : OAI22_X1 port map( A1 => n7476, A2 => n5690, B1 => n5770, B2 => n5689
                           , ZN => n2040);
   U230 : OAI22_X1 port map( A1 => n7477, A2 => n5690, B1 => n5772, B2 => n5689
                           , ZN => n2039);
   U231 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n5703, ZN 
                           => n5811);
   U232 : NAND2_X1 port map( A1 => n5704, A2 => n5811, ZN => n5691);
   U233 : OAI22_X1 port map( A1 => n7960, A2 => n5693, B1 => n5788, B2 => n5692
                           , ZN => n2038);
   U234 : OAI22_X1 port map( A1 => n7961, A2 => n5693, B1 => n5740, B2 => n5691
                           , ZN => n2037);
   U235 : OAI22_X1 port map( A1 => n8207, A2 => n5693, B1 => n5741, B2 => n5692
                           , ZN => n2036);
   U236 : OAI22_X1 port map( A1 => n7962, A2 => n5693, B1 => n5742, B2 => n5691
                           , ZN => n2035);
   U237 : OAI22_X1 port map( A1 => n8208, A2 => n5693, B1 => n5743, B2 => n5692
                           , ZN => n2034);
   U238 : OAI22_X1 port map( A1 => n8209, A2 => n5693, B1 => n5744, B2 => n5691
                           , ZN => n2033);
   U239 : OAI22_X1 port map( A1 => n7963, A2 => n5693, B1 => n5745, B2 => n5692
                           , ZN => n2032);
   U240 : OAI22_X1 port map( A1 => n7964, A2 => n5693, B1 => n5746, B2 => n5691
                           , ZN => n2031);
   U241 : OAI22_X1 port map( A1 => n7965, A2 => n5693, B1 => n5747, B2 => n5692
                           , ZN => n2030);
   U242 : OAI22_X1 port map( A1 => n7966, A2 => n5693, B1 => n5748, B2 => n5691
                           , ZN => n2029);
   U243 : OAI22_X1 port map( A1 => n7967, A2 => n5693, B1 => n5749, B2 => n5691
                           , ZN => n2028);
   U244 : OAI22_X1 port map( A1 => n7478, A2 => n5693, B1 => n5750, B2 => n5692
                           , ZN => n2027);
   U245 : OAI22_X1 port map( A1 => n7479, A2 => n5693, B1 => n5751, B2 => n5691
                           , ZN => n2026);
   U246 : OAI22_X1 port map( A1 => n7968, A2 => n5693, B1 => n5752, B2 => n5692
                           , ZN => n2025);
   U247 : OAI22_X1 port map( A1 => n8210, A2 => n5693, B1 => n5753, B2 => n5691
                           , ZN => n2024);
   U248 : OAI22_X1 port map( A1 => n7969, A2 => n5693, B1 => n5754, B2 => n5692
                           , ZN => n2023);
   U249 : OAI22_X1 port map( A1 => n8211, A2 => n5693, B1 => n5755, B2 => n5691
                           , ZN => n2022);
   U250 : OAI22_X1 port map( A1 => n7970, A2 => n5693, B1 => n5756, B2 => n5691
                           , ZN => n2021);
   U251 : OAI22_X1 port map( A1 => n8212, A2 => n5693, B1 => n5757, B2 => n5691
                           , ZN => n2020);
   U252 : OAI22_X1 port map( A1 => n7971, A2 => n5693, B1 => n5758, B2 => n5691
                           , ZN => n2019);
   U253 : OAI22_X1 port map( A1 => n7972, A2 => n5693, B1 => n5759, B2 => n5691
                           , ZN => n2018);
   U254 : OAI22_X1 port map( A1 => n8213, A2 => n5693, B1 => n5760, B2 => n5691
                           , ZN => n2017);
   U255 : OAI22_X1 port map( A1 => n7973, A2 => n5693, B1 => n5762, B2 => n5691
                           , ZN => n2016);
   U256 : OAI22_X1 port map( A1 => n8214, A2 => n5693, B1 => n5763, B2 => n5692
                           , ZN => n2015);
   U257 : OAI22_X1 port map( A1 => n7974, A2 => n5693, B1 => n5764, B2 => n5692
                           , ZN => n2014);
   U258 : OAI22_X1 port map( A1 => n8215, A2 => n5693, B1 => n5765, B2 => n5692
                           , ZN => n2013);
   U259 : OAI22_X1 port map( A1 => n8216, A2 => n5693, B1 => n5766, B2 => n5692
                           , ZN => n2012);
   U260 : OAI22_X1 port map( A1 => n7975, A2 => n5693, B1 => n5767, B2 => n5692
                           , ZN => n2011);
   U261 : OAI22_X1 port map( A1 => n7976, A2 => n5693, B1 => n5768, B2 => n5692
                           , ZN => n2010);
   U262 : OAI22_X1 port map( A1 => n8217, A2 => n5693, B1 => n5769, B2 => n5692
                           , ZN => n2009);
   U263 : OAI22_X1 port map( A1 => n7739, A2 => n5693, B1 => n5770, B2 => n5692
                           , ZN => n2008);
   U264 : OAI22_X1 port map( A1 => n7977, A2 => n5693, B1 => n5772, B2 => n5692
                           , ZN => n2007);
   U265 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n5694, A3 => n5703, ZN => 
                           n5815);
   U266 : NAND2_X1 port map( A1 => n5704, A2 => n5815, ZN => n5695);
   U267 : CLKBUF_X1 port map( A => n5695, Z => n5696);
   U268 : OAI22_X1 port map( A1 => n7978, A2 => n5697, B1 => n5825, B2 => n5696
                           , ZN => n2006);
   U269 : OAI22_X1 port map( A1 => n8218, A2 => n5697, B1 => n5740, B2 => n5695
                           , ZN => n2005);
   U270 : OAI22_X1 port map( A1 => n8219, A2 => n5697, B1 => n5741, B2 => n5696
                           , ZN => n2004);
   U271 : OAI22_X1 port map( A1 => n7740, A2 => n5697, B1 => n5742, B2 => n5695
                           , ZN => n2003);
   U272 : OAI22_X1 port map( A1 => n7979, A2 => n5697, B1 => n5743, B2 => n5696
                           , ZN => n2002);
   U273 : OAI22_X1 port map( A1 => n7741, A2 => n5697, B1 => n5744, B2 => n5695
                           , ZN => n2001);
   U274 : OAI22_X1 port map( A1 => n7742, A2 => n5697, B1 => n5745, B2 => n5696
                           , ZN => n2000);
   U275 : OAI22_X1 port map( A1 => n7980, A2 => n5697, B1 => n5746, B2 => n5695
                           , ZN => n1999);
   U276 : OAI22_X1 port map( A1 => n8220, A2 => n5697, B1 => n5747, B2 => n5696
                           , ZN => n1998);
   U277 : OAI22_X1 port map( A1 => n7743, A2 => n5697, B1 => n5748, B2 => n5695
                           , ZN => n1997);
   U278 : OAI22_X1 port map( A1 => n8221, A2 => n5697, B1 => n5749, B2 => n5695
                           , ZN => n1996);
   U279 : OAI22_X1 port map( A1 => n7981, A2 => n5697, B1 => n5750, B2 => n5696
                           , ZN => n1995);
   U280 : OAI22_X1 port map( A1 => n8222, A2 => n5697, B1 => n5751, B2 => n5695
                           , ZN => n1994);
   U281 : OAI22_X1 port map( A1 => n8223, A2 => n5697, B1 => n5752, B2 => n5696
                           , ZN => n1993);
   U282 : OAI22_X1 port map( A1 => n7744, A2 => n5697, B1 => n5753, B2 => n5695
                           , ZN => n1992);
   U283 : OAI22_X1 port map( A1 => n7982, A2 => n5697, B1 => n5754, B2 => n5696
                           , ZN => n1991);
   U284 : OAI22_X1 port map( A1 => n7983, A2 => n5697, B1 => n5755, B2 => n5695
                           , ZN => n1990);
   U285 : OAI22_X1 port map( A1 => n8224, A2 => n5697, B1 => n5756, B2 => n5695
                           , ZN => n1989);
   U286 : OAI22_X1 port map( A1 => n7745, A2 => n5697, B1 => n5757, B2 => n5695
                           , ZN => n1988);
   U287 : OAI22_X1 port map( A1 => n8225, A2 => n5697, B1 => n5758, B2 => n5695
                           , ZN => n1987);
   U288 : OAI22_X1 port map( A1 => n7480, A2 => n5697, B1 => n5759, B2 => n5695
                           , ZN => n1986);
   U289 : OAI22_X1 port map( A1 => n7481, A2 => n5697, B1 => n5760, B2 => n5695
                           , ZN => n1985);
   U290 : OAI22_X1 port map( A1 => n8226, A2 => n5697, B1 => n5762, B2 => n5695
                           , ZN => n1984);
   U291 : OAI22_X1 port map( A1 => n7482, A2 => n5697, B1 => n5763, B2 => n5696
                           , ZN => n1983);
   U292 : OAI22_X1 port map( A1 => n7746, A2 => n5697, B1 => n5764, B2 => n5696
                           , ZN => n1982);
   U293 : OAI22_X1 port map( A1 => n7984, A2 => n5697, B1 => n5765, B2 => n5696
                           , ZN => n1981);
   U294 : OAI22_X1 port map( A1 => n7985, A2 => n5697, B1 => n5766, B2 => n5696
                           , ZN => n1980);
   U295 : OAI22_X1 port map( A1 => n8227, A2 => n5697, B1 => n5767, B2 => n5696
                           , ZN => n1979);
   U296 : OAI22_X1 port map( A1 => n8228, A2 => n5697, B1 => n5768, B2 => n5696
                           , ZN => n1978);
   U297 : OAI22_X1 port map( A1 => n7747, A2 => n5697, B1 => n5769, B2 => n5696
                           , ZN => n1977);
   U298 : OAI22_X1 port map( A1 => n7986, A2 => n5697, B1 => n5770, B2 => n5696
                           , ZN => n1976);
   U299 : OAI22_X1 port map( A1 => n7987, A2 => n5697, B1 => n5772, B2 => n5696
                           , ZN => n1975);
   U300 : NOR2_X1 port map( A1 => n5703, A2 => n5698, ZN => n5819);
   U301 : NAND2_X1 port map( A1 => n5704, A2 => n5819, ZN => n5699);
   U302 : CLKBUF_X1 port map( A => n5699, Z => n5700);
   U303 : OAI22_X1 port map( A1 => n7988, A2 => n5701, B1 => n5788, B2 => n5700
                           , ZN => n1974);
   U304 : OAI22_X1 port map( A1 => n7989, A2 => n5701, B1 => n5740, B2 => n5699
                           , ZN => n1973);
   U305 : OAI22_X1 port map( A1 => n7990, A2 => n5701, B1 => n5741, B2 => n5700
                           , ZN => n1972);
   U306 : OAI22_X1 port map( A1 => n8229, A2 => n5701, B1 => n5742, B2 => n5699
                           , ZN => n1971);
   U307 : OAI22_X1 port map( A1 => n7991, A2 => n5701, B1 => n5743, B2 => n5700
                           , ZN => n1970);
   U308 : OAI22_X1 port map( A1 => n8230, A2 => n5701, B1 => n5744, B2 => n5699
                           , ZN => n1969);
   U309 : OAI22_X1 port map( A1 => n7992, A2 => n5701, B1 => n5745, B2 => n5700
                           , ZN => n1968);
   U310 : OAI22_X1 port map( A1 => n8231, A2 => n5701, B1 => n5746, B2 => n5699
                           , ZN => n1967);
   U311 : OAI22_X1 port map( A1 => n8232, A2 => n5701, B1 => n5747, B2 => n5700
                           , ZN => n1966);
   U312 : OAI22_X1 port map( A1 => n7993, A2 => n5701, B1 => n5748, B2 => n5699
                           , ZN => n1965);
   U313 : OAI22_X1 port map( A1 => n7994, A2 => n5701, B1 => n5749, B2 => n5699
                           , ZN => n1964);
   U314 : OAI22_X1 port map( A1 => n8233, A2 => n5701, B1 => n5750, B2 => n5700
                           , ZN => n1963);
   U315 : OAI22_X1 port map( A1 => n8234, A2 => n5701, B1 => n5751, B2 => n5699
                           , ZN => n1962);
   U316 : OAI22_X1 port map( A1 => n7995, A2 => n5701, B1 => n5752, B2 => n5700
                           , ZN => n1961);
   U317 : OAI22_X1 port map( A1 => n8235, A2 => n5701, B1 => n5753, B2 => n5699
                           , ZN => n1960);
   U318 : OAI22_X1 port map( A1 => n8236, A2 => n5701, B1 => n5754, B2 => n5700
                           , ZN => n1959);
   U319 : OAI22_X1 port map( A1 => n8237, A2 => n5701, B1 => n5755, B2 => n5699
                           , ZN => n1958);
   U320 : OAI22_X1 port map( A1 => n7996, A2 => n5701, B1 => n5756, B2 => n5699
                           , ZN => n1957);
   U321 : OAI22_X1 port map( A1 => n7997, A2 => n5701, B1 => n5757, B2 => n5699
                           , ZN => n1956);
   U322 : OAI22_X1 port map( A1 => n7998, A2 => n5701, B1 => n5758, B2 => n5699
                           , ZN => n1955);
   U323 : OAI22_X1 port map( A1 => n7999, A2 => n5701, B1 => n5759, B2 => n5699
                           , ZN => n1954);
   U324 : OAI22_X1 port map( A1 => n8000, A2 => n5701, B1 => n5760, B2 => n5699
                           , ZN => n1953);
   U325 : OAI22_X1 port map( A1 => n8001, A2 => n5701, B1 => n5762, B2 => n5699
                           , ZN => n1952);
   U326 : OAI22_X1 port map( A1 => n8002, A2 => n5701, B1 => n5763, B2 => n5700
                           , ZN => n1951);
   U327 : OAI22_X1 port map( A1 => n8238, A2 => n5701, B1 => n5764, B2 => n5700
                           , ZN => n1950);
   U328 : OAI22_X1 port map( A1 => n8003, A2 => n5701, B1 => n5765, B2 => n5700
                           , ZN => n1949);
   U329 : OAI22_X1 port map( A1 => n8239, A2 => n5701, B1 => n5766, B2 => n5700
                           , ZN => n1948);
   U330 : OAI22_X1 port map( A1 => n8240, A2 => n5701, B1 => n5767, B2 => n5700
                           , ZN => n1947);
   U331 : OAI22_X1 port map( A1 => n8241, A2 => n5701, B1 => n5768, B2 => n5700
                           , ZN => n1946);
   U332 : OAI22_X1 port map( A1 => n8004, A2 => n5701, B1 => n5769, B2 => n5700
                           , ZN => n1945);
   U333 : OAI22_X1 port map( A1 => n8242, A2 => n5701, B1 => n5770, B2 => n5700
                           , ZN => n1944);
   U334 : OAI22_X1 port map( A1 => n8005, A2 => n5701, B1 => n5772, B2 => n5700
                           , ZN => n1943);
   U335 : NOR2_X1 port map( A1 => n5703, A2 => n5702, ZN => n5824);
   U336 : NAND2_X1 port map( A1 => n5704, A2 => n5824, ZN => n5705);
   U337 : CLKBUF_X1 port map( A => n5705, Z => n5706);
   U338 : OAI22_X1 port map( A1 => n8243, A2 => n5707, B1 => n5825, B2 => n5706
                           , ZN => n1942);
   U339 : OAI22_X1 port map( A1 => n7748, A2 => n5707, B1 => n5740, B2 => n5705
                           , ZN => n1941);
   U340 : OAI22_X1 port map( A1 => n7483, A2 => n5707, B1 => n5741, B2 => n5706
                           , ZN => n1940);
   U341 : OAI22_X1 port map( A1 => n8006, A2 => n5707, B1 => n5742, B2 => n5705
                           , ZN => n1939);
   U342 : OAI22_X1 port map( A1 => n7749, A2 => n5707, B1 => n5743, B2 => n5706
                           , ZN => n1938);
   U343 : OAI22_X1 port map( A1 => n8007, A2 => n5707, B1 => n5744, B2 => n5705
                           , ZN => n1937);
   U344 : OAI22_X1 port map( A1 => n8244, A2 => n5707, B1 => n5745, B2 => n5706
                           , ZN => n1936);
   U345 : OAI22_X1 port map( A1 => n8245, A2 => n5707, B1 => n5746, B2 => n5705
                           , ZN => n1935);
   U346 : OAI22_X1 port map( A1 => n7750, A2 => n5707, B1 => n5747, B2 => n5706
                           , ZN => n1934);
   U347 : OAI22_X1 port map( A1 => n7484, A2 => n5707, B1 => n5748, B2 => n5705
                           , ZN => n1933);
   U348 : OAI22_X1 port map( A1 => n7751, A2 => n5707, B1 => n5749, B2 => n5705
                           , ZN => n1932);
   U349 : OAI22_X1 port map( A1 => n8246, A2 => n5707, B1 => n5750, B2 => n5706
                           , ZN => n1931);
   U350 : OAI22_X1 port map( A1 => n7485, A2 => n5707, B1 => n5751, B2 => n5705
                           , ZN => n1930);
   U351 : OAI22_X1 port map( A1 => n7752, A2 => n5707, B1 => n5752, B2 => n5706
                           , ZN => n1929);
   U352 : OAI22_X1 port map( A1 => n7753, A2 => n5707, B1 => n5753, B2 => n5705
                           , ZN => n1928);
   U353 : OAI22_X1 port map( A1 => n8247, A2 => n5707, B1 => n5754, B2 => n5706
                           , ZN => n1927);
   U354 : OAI22_X1 port map( A1 => n8008, A2 => n5707, B1 => n5755, B2 => n5705
                           , ZN => n1926);
   U355 : OAI22_X1 port map( A1 => n7486, A2 => n5707, B1 => n5756, B2 => n5705
                           , ZN => n1925);
   U356 : OAI22_X1 port map( A1 => n7487, A2 => n5707, B1 => n5757, B2 => n5705
                           , ZN => n1924);
   U357 : OAI22_X1 port map( A1 => n7754, A2 => n5707, B1 => n5758, B2 => n5705
                           , ZN => n1923);
   U358 : OAI22_X1 port map( A1 => n8248, A2 => n5707, B1 => n5759, B2 => n5705
                           , ZN => n1922);
   U359 : OAI22_X1 port map( A1 => n8249, A2 => n5707, B1 => n5760, B2 => n5705
                           , ZN => n1921);
   U360 : OAI22_X1 port map( A1 => n8250, A2 => n5707, B1 => n5762, B2 => n5705
                           , ZN => n1920);
   U361 : OAI22_X1 port map( A1 => n8251, A2 => n5707, B1 => n5763, B2 => n5706
                           , ZN => n1919);
   U362 : OAI22_X1 port map( A1 => n7488, A2 => n5707, B1 => n5764, B2 => n5706
                           , ZN => n1918);
   U363 : OAI22_X1 port map( A1 => n8252, A2 => n5707, B1 => n5765, B2 => n5706
                           , ZN => n1917);
   U364 : OAI22_X1 port map( A1 => n7755, A2 => n5707, B1 => n5766, B2 => n5706
                           , ZN => n1916);
   U365 : OAI22_X1 port map( A1 => n7489, A2 => n5707, B1 => n5767, B2 => n5706
                           , ZN => n1915);
   U366 : OAI22_X1 port map( A1 => n8009, A2 => n5707, B1 => n5768, B2 => n5706
                           , ZN => n1914);
   U367 : OAI22_X1 port map( A1 => n7756, A2 => n5707, B1 => n5769, B2 => n5706
                           , ZN => n1913);
   U368 : OAI22_X1 port map( A1 => n8253, A2 => n5707, B1 => n5770, B2 => n5706
                           , ZN => n1912);
   U369 : OAI22_X1 port map( A1 => n7757, A2 => n5707, B1 => n5772, B2 => n5706
                           , ZN => n1911);
   U370 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(3), ZN => 
                           n5792);
   U371 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n5792, ZN => n5729);
   U372 : NAND2_X1 port map( A1 => n5794, A2 => n5729, ZN => n5708);
   U373 : CLKBUF_X1 port map( A => n5708, Z => n5709);
   U374 : OAI22_X1 port map( A1 => n7490, A2 => n5710, B1 => n5788, B2 => n5709
                           , ZN => n1910);
   U375 : OAI22_X1 port map( A1 => n8254, A2 => n5710, B1 => n5740, B2 => n5708
                           , ZN => n1909);
   U376 : OAI22_X1 port map( A1 => n7758, A2 => n5710, B1 => n5741, B2 => n5709
                           , ZN => n1908);
   U377 : OAI22_X1 port map( A1 => n8010, A2 => n5710, B1 => n5742, B2 => n5708
                           , ZN => n1907);
   U378 : OAI22_X1 port map( A1 => n7759, A2 => n5710, B1 => n5743, B2 => n5709
                           , ZN => n1906);
   U379 : OAI22_X1 port map( A1 => n7760, A2 => n5710, B1 => n5744, B2 => n5708
                           , ZN => n1905);
   U380 : OAI22_X1 port map( A1 => n7761, A2 => n5710, B1 => n5745, B2 => n5709
                           , ZN => n1904);
   U381 : OAI22_X1 port map( A1 => n8255, A2 => n5710, B1 => n5746, B2 => n5708
                           , ZN => n1903);
   U382 : OAI22_X1 port map( A1 => n7762, A2 => n5710, B1 => n5747, B2 => n5709
                           , ZN => n1902);
   U383 : OAI22_X1 port map( A1 => n8256, A2 => n5710, B1 => n5748, B2 => n5708
                           , ZN => n1901);
   U384 : OAI22_X1 port map( A1 => n8257, A2 => n5710, B1 => n5749, B2 => n5708
                           , ZN => n1900);
   U385 : OAI22_X1 port map( A1 => n8258, A2 => n5710, B1 => n5750, B2 => n5709
                           , ZN => n1899);
   U386 : OAI22_X1 port map( A1 => n8011, A2 => n5710, B1 => n5751, B2 => n5708
                           , ZN => n1898);
   U387 : OAI22_X1 port map( A1 => n7491, A2 => n5710, B1 => n5752, B2 => n5709
                           , ZN => n1897);
   U388 : OAI22_X1 port map( A1 => n7763, A2 => n5710, B1 => n5753, B2 => n5708
                           , ZN => n1896);
   U389 : OAI22_X1 port map( A1 => n8259, A2 => n5710, B1 => n5754, B2 => n5709
                           , ZN => n1895);
   U390 : OAI22_X1 port map( A1 => n7492, A2 => n5710, B1 => n5755, B2 => n5708
                           , ZN => n1894);
   U391 : OAI22_X1 port map( A1 => n7764, A2 => n5710, B1 => n5756, B2 => n5708
                           , ZN => n1893);
   U392 : OAI22_X1 port map( A1 => n7765, A2 => n5710, B1 => n5757, B2 => n5708
                           , ZN => n1892);
   U393 : OAI22_X1 port map( A1 => n7766, A2 => n5710, B1 => n5758, B2 => n5708
                           , ZN => n1891);
   U394 : OAI22_X1 port map( A1 => n7493, A2 => n5710, B1 => n5759, B2 => n5708
                           , ZN => n1890);
   U395 : OAI22_X1 port map( A1 => n8012, A2 => n5710, B1 => n5760, B2 => n5708
                           , ZN => n1889);
   U396 : OAI22_X1 port map( A1 => n8260, A2 => n5710, B1 => n5762, B2 => n5708
                           , ZN => n1888);
   U397 : OAI22_X1 port map( A1 => n8261, A2 => n5710, B1 => n5763, B2 => n5709
                           , ZN => n1887);
   U398 : OAI22_X1 port map( A1 => n8013, A2 => n5710, B1 => n5764, B2 => n5709
                           , ZN => n1886);
   U399 : OAI22_X1 port map( A1 => n7494, A2 => n5710, B1 => n5765, B2 => n5709
                           , ZN => n1885);
   U400 : OAI22_X1 port map( A1 => n7767, A2 => n5710, B1 => n5766, B2 => n5709
                           , ZN => n1884);
   U401 : OAI22_X1 port map( A1 => n7495, A2 => n5710, B1 => n5767, B2 => n5709
                           , ZN => n1883);
   U402 : OAI22_X1 port map( A1 => n8262, A2 => n5710, B1 => n5768, B2 => n5709
                           , ZN => n1882);
   U403 : OAI22_X1 port map( A1 => n8014, A2 => n5710, B1 => n5769, B2 => n5709
                           , ZN => n1881);
   U404 : OAI22_X1 port map( A1 => n7768, A2 => n5710, B1 => n5770, B2 => n5709
                           , ZN => n1880);
   U405 : OAI22_X1 port map( A1 => n7769, A2 => n5710, B1 => n5772, B2 => n5709
                           , ZN => n1879);
   U406 : NAND2_X1 port map( A1 => n5798, A2 => n5729, ZN => n5711);
   U407 : CLKBUF_X1 port map( A => n5711, Z => n5712);
   U408 : OAI22_X1 port map( A1 => n7770, A2 => n5713, B1 => n5825, B2 => n5712
                           , ZN => n1878);
   U409 : OAI22_X1 port map( A1 => n7496, A2 => n5713, B1 => n5740, B2 => n5711
                           , ZN => n1877);
   U410 : OAI22_X1 port map( A1 => n7497, A2 => n5713, B1 => n5741, B2 => n5712
                           , ZN => n1876);
   U411 : OAI22_X1 port map( A1 => n7771, A2 => n5713, B1 => n5742, B2 => n5711
                           , ZN => n1875);
   U412 : OAI22_X1 port map( A1 => n7772, A2 => n5713, B1 => n5743, B2 => n5712
                           , ZN => n1874);
   U413 : OAI22_X1 port map( A1 => n7498, A2 => n5713, B1 => n5744, B2 => n5711
                           , ZN => n1873);
   U414 : OAI22_X1 port map( A1 => n7773, A2 => n5713, B1 => n5745, B2 => n5712
                           , ZN => n1872);
   U415 : OAI22_X1 port map( A1 => n7774, A2 => n5713, B1 => n5746, B2 => n5711
                           , ZN => n1871);
   U416 : OAI22_X1 port map( A1 => n7499, A2 => n5713, B1 => n5747, B2 => n5712
                           , ZN => n1870);
   U417 : OAI22_X1 port map( A1 => n7500, A2 => n5713, B1 => n5748, B2 => n5711
                           , ZN => n1869);
   U418 : OAI22_X1 port map( A1 => n7775, A2 => n5713, B1 => n5749, B2 => n5711
                           , ZN => n1868);
   U419 : OAI22_X1 port map( A1 => n7501, A2 => n5713, B1 => n5750, B2 => n5712
                           , ZN => n1867);
   U420 : OAI22_X1 port map( A1 => n7776, A2 => n5713, B1 => n5751, B2 => n5711
                           , ZN => n1866);
   U421 : OAI22_X1 port map( A1 => n7777, A2 => n5713, B1 => n5752, B2 => n5712
                           , ZN => n1865);
   U422 : OAI22_X1 port map( A1 => n7502, A2 => n5713, B1 => n5753, B2 => n5711
                           , ZN => n1864);
   U423 : OAI22_X1 port map( A1 => n7503, A2 => n5713, B1 => n5754, B2 => n5712
                           , ZN => n1863);
   U424 : OAI22_X1 port map( A1 => n7778, A2 => n5713, B1 => n5755, B2 => n5711
                           , ZN => n1862);
   U425 : OAI22_X1 port map( A1 => n7504, A2 => n5713, B1 => n5756, B2 => n5711
                           , ZN => n1861);
   U426 : OAI22_X1 port map( A1 => n7779, A2 => n5713, B1 => n5757, B2 => n5711
                           , ZN => n1860);
   U427 : OAI22_X1 port map( A1 => n7505, A2 => n5713, B1 => n5758, B2 => n5711
                           , ZN => n1859);
   U428 : OAI22_X1 port map( A1 => n7780, A2 => n5713, B1 => n5759, B2 => n5711
                           , ZN => n1858);
   U429 : OAI22_X1 port map( A1 => n7506, A2 => n5713, B1 => n5760, B2 => n5711
                           , ZN => n1857);
   U430 : OAI22_X1 port map( A1 => n7507, A2 => n5713, B1 => n5762, B2 => n5711
                           , ZN => n1856);
   U431 : OAI22_X1 port map( A1 => n7508, A2 => n5713, B1 => n5763, B2 => n5712
                           , ZN => n1855);
   U432 : OAI22_X1 port map( A1 => n7509, A2 => n5713, B1 => n5764, B2 => n5712
                           , ZN => n1854);
   U433 : OAI22_X1 port map( A1 => n7781, A2 => n5713, B1 => n5765, B2 => n5712
                           , ZN => n1853);
   U434 : OAI22_X1 port map( A1 => n7510, A2 => n5713, B1 => n5766, B2 => n5712
                           , ZN => n1852);
   U435 : OAI22_X1 port map( A1 => n7511, A2 => n5713, B1 => n5767, B2 => n5712
                           , ZN => n1851);
   U436 : OAI22_X1 port map( A1 => n7782, A2 => n5713, B1 => n5768, B2 => n5712
                           , ZN => n1850);
   U437 : OAI22_X1 port map( A1 => n7512, A2 => n5713, B1 => n5769, B2 => n5712
                           , ZN => n1849);
   U438 : OAI22_X1 port map( A1 => n7513, A2 => n5713, B1 => n5770, B2 => n5712
                           , ZN => n1848);
   U439 : OAI22_X1 port map( A1 => n7514, A2 => n5713, B1 => n5772, B2 => n5712
                           , ZN => n1847);
   U440 : NAND2_X1 port map( A1 => n5802, A2 => n5729, ZN => n5714);
   U441 : CLKBUF_X1 port map( A => n5714, Z => n5715);
   U442 : OAI22_X1 port map( A1 => n8263, A2 => n5716, B1 => n5825, B2 => n5715
                           , ZN => n1846);
   U443 : OAI22_X1 port map( A1 => n7783, A2 => n5716, B1 => n5740, B2 => n5714
                           , ZN => n1845);
   U444 : OAI22_X1 port map( A1 => n7515, A2 => n5716, B1 => n5741, B2 => n5715
                           , ZN => n1844);
   U445 : OAI22_X1 port map( A1 => n7784, A2 => n5716, B1 => n5742, B2 => n5714
                           , ZN => n1843);
   U446 : OAI22_X1 port map( A1 => n7516, A2 => n5716, B1 => n5743, B2 => n5715
                           , ZN => n1842);
   U447 : OAI22_X1 port map( A1 => n7785, A2 => n5716, B1 => n5744, B2 => n5714
                           , ZN => n1841);
   U448 : OAI22_X1 port map( A1 => n7517, A2 => n5716, B1 => n5745, B2 => n5715
                           , ZN => n1840);
   U449 : OAI22_X1 port map( A1 => n8015, A2 => n5716, B1 => n5746, B2 => n5714
                           , ZN => n1839);
   U450 : OAI22_X1 port map( A1 => n8016, A2 => n5716, B1 => n5747, B2 => n5715
                           , ZN => n1838);
   U451 : OAI22_X1 port map( A1 => n7518, A2 => n5716, B1 => n5748, B2 => n5714
                           , ZN => n1837);
   U452 : OAI22_X1 port map( A1 => n7519, A2 => n5716, B1 => n5749, B2 => n5714
                           , ZN => n1836);
   U453 : OAI22_X1 port map( A1 => n7520, A2 => n5716, B1 => n5750, B2 => n5715
                           , ZN => n1835);
   U454 : OAI22_X1 port map( A1 => n7786, A2 => n5716, B1 => n5751, B2 => n5714
                           , ZN => n1834);
   U455 : OAI22_X1 port map( A1 => n8264, A2 => n5716, B1 => n5752, B2 => n5715
                           , ZN => n1833);
   U456 : OAI22_X1 port map( A1 => n7787, A2 => n5716, B1 => n5753, B2 => n5714
                           , ZN => n1832);
   U457 : OAI22_X1 port map( A1 => n7788, A2 => n5716, B1 => n5754, B2 => n5715
                           , ZN => n1831);
   U458 : OAI22_X1 port map( A1 => n7521, A2 => n5716, B1 => n5755, B2 => n5714
                           , ZN => n1830);
   U459 : OAI22_X1 port map( A1 => n7522, A2 => n5716, B1 => n5756, B2 => n5714
                           , ZN => n1829);
   U460 : OAI22_X1 port map( A1 => n7789, A2 => n5716, B1 => n5757, B2 => n5714
                           , ZN => n1828);
   U461 : OAI22_X1 port map( A1 => n8017, A2 => n5716, B1 => n5758, B2 => n5714
                           , ZN => n1827);
   U462 : OAI22_X1 port map( A1 => n7790, A2 => n5716, B1 => n5759, B2 => n5714
                           , ZN => n1826);
   U463 : OAI22_X1 port map( A1 => n7523, A2 => n5716, B1 => n5760, B2 => n5714
                           , ZN => n1825);
   U464 : OAI22_X1 port map( A1 => n7791, A2 => n5716, B1 => n5762, B2 => n5714
                           , ZN => n1824);
   U465 : OAI22_X1 port map( A1 => n7792, A2 => n5716, B1 => n5763, B2 => n5715
                           , ZN => n1823);
   U466 : OAI22_X1 port map( A1 => n7793, A2 => n5716, B1 => n5764, B2 => n5715
                           , ZN => n1822);
   U467 : OAI22_X1 port map( A1 => n8265, A2 => n5716, B1 => n5765, B2 => n5715
                           , ZN => n1821);
   U468 : OAI22_X1 port map( A1 => n7524, A2 => n5716, B1 => n5766, B2 => n5715
                           , ZN => n1820);
   U469 : OAI22_X1 port map( A1 => n7794, A2 => n5716, B1 => n5767, B2 => n5715
                           , ZN => n1819);
   U470 : OAI22_X1 port map( A1 => n7795, A2 => n5716, B1 => n5768, B2 => n5715
                           , ZN => n1818);
   U471 : OAI22_X1 port map( A1 => n8018, A2 => n5716, B1 => n5769, B2 => n5715
                           , ZN => n1817);
   U472 : OAI22_X1 port map( A1 => n8019, A2 => n5716, B1 => n5770, B2 => n5715
                           , ZN => n1816);
   U473 : OAI22_X1 port map( A1 => n8020, A2 => n5716, B1 => n5772, B2 => n5715
                           , ZN => n1815);
   U474 : NAND2_X1 port map( A1 => n5807, A2 => n5729, ZN => n5717);
   U475 : CLKBUF_X1 port map( A => n5717, Z => n5718);
   U476 : OAI22_X1 port map( A1 => n7796, A2 => n5719, B1 => n5825, B2 => n5718
                           , ZN => n1814);
   U477 : OAI22_X1 port map( A1 => n7525, A2 => n5719, B1 => n5826, B2 => n5717
                           , ZN => n1813);
   U478 : CLKBUF_X1 port map( A => n5741, Z => n5827);
   U479 : OAI22_X1 port map( A1 => n8021, A2 => n5719, B1 => n5827, B2 => n5718
                           , ZN => n1812);
   U480 : CLKBUF_X1 port map( A => n5742, Z => n5828);
   U481 : OAI22_X1 port map( A1 => n7526, A2 => n5719, B1 => n5828, B2 => n5717
                           , ZN => n1811);
   U482 : CLKBUF_X1 port map( A => n5743, Z => n5829);
   U483 : OAI22_X1 port map( A1 => n8266, A2 => n5719, B1 => n5829, B2 => n5718
                           , ZN => n1810);
   U484 : CLKBUF_X1 port map( A => n5744, Z => n5830);
   U485 : OAI22_X1 port map( A1 => n7797, A2 => n5719, B1 => n5830, B2 => n5717
                           , ZN => n1809);
   U486 : CLKBUF_X1 port map( A => n5745, Z => n5831);
   U487 : OAI22_X1 port map( A1 => n8267, A2 => n5719, B1 => n5831, B2 => n5718
                           , ZN => n1808);
   U488 : CLKBUF_X1 port map( A => n5746, Z => n5832);
   U489 : OAI22_X1 port map( A1 => n7798, A2 => n5719, B1 => n5832, B2 => n5717
                           , ZN => n1807);
   U490 : CLKBUF_X1 port map( A => n5747, Z => n5833);
   U491 : OAI22_X1 port map( A1 => n7527, A2 => n5719, B1 => n5833, B2 => n5718
                           , ZN => n1806);
   U492 : CLKBUF_X1 port map( A => n5748, Z => n5834);
   U493 : OAI22_X1 port map( A1 => n8022, A2 => n5719, B1 => n5834, B2 => n5717
                           , ZN => n1805);
   U494 : CLKBUF_X1 port map( A => n5749, Z => n5835);
   U495 : OAI22_X1 port map( A1 => n7528, A2 => n5719, B1 => n5835, B2 => n5717
                           , ZN => n1804);
   U496 : CLKBUF_X1 port map( A => n5750, Z => n5836);
   U497 : OAI22_X1 port map( A1 => n7799, A2 => n5719, B1 => n5836, B2 => n5718
                           , ZN => n1803);
   U498 : CLKBUF_X1 port map( A => n5751, Z => n5837);
   U499 : OAI22_X1 port map( A1 => n7800, A2 => n5719, B1 => n5837, B2 => n5717
                           , ZN => n1802);
   U500 : CLKBUF_X1 port map( A => n5752, Z => n5838);
   U501 : OAI22_X1 port map( A1 => n7529, A2 => n5719, B1 => n5838, B2 => n5718
                           , ZN => n1801);
   U502 : CLKBUF_X1 port map( A => n5753, Z => n5839);
   U503 : OAI22_X1 port map( A1 => n7530, A2 => n5719, B1 => n5839, B2 => n5717
                           , ZN => n1800);
   U504 : OAI22_X1 port map( A1 => n7531, A2 => n5719, B1 => n5840, B2 => n5718
                           , ZN => n1799);
   U505 : CLKBUF_X1 port map( A => n5755, Z => n5841);
   U506 : OAI22_X1 port map( A1 => n7801, A2 => n5719, B1 => n5841, B2 => n5717
                           , ZN => n1798);
   U507 : CLKBUF_X1 port map( A => n5756, Z => n5842);
   U508 : OAI22_X1 port map( A1 => n7802, A2 => n5719, B1 => n5842, B2 => n5717
                           , ZN => n1797);
   U509 : CLKBUF_X1 port map( A => n5757, Z => n5843);
   U510 : OAI22_X1 port map( A1 => n8268, A2 => n5719, B1 => n5843, B2 => n5717
                           , ZN => n1796);
   U511 : CLKBUF_X1 port map( A => n5758, Z => n5844);
   U512 : OAI22_X1 port map( A1 => n7803, A2 => n5719, B1 => n5844, B2 => n5717
                           , ZN => n1795);
   U513 : CLKBUF_X1 port map( A => n5759, Z => n5845);
   U514 : OAI22_X1 port map( A1 => n8269, A2 => n5719, B1 => n5845, B2 => n5717
                           , ZN => n1794);
   U515 : CLKBUF_X1 port map( A => n5760, Z => n5846);
   U516 : OAI22_X1 port map( A1 => n7804, A2 => n5719, B1 => n5846, B2 => n5717
                           , ZN => n1793);
   U517 : CLKBUF_X1 port map( A => n5762, Z => n5848);
   U518 : OAI22_X1 port map( A1 => n7532, A2 => n5719, B1 => n5848, B2 => n5717
                           , ZN => n1792);
   U519 : CLKBUF_X1 port map( A => n5763, Z => n5849);
   U520 : OAI22_X1 port map( A1 => n7533, A2 => n5719, B1 => n5849, B2 => n5718
                           , ZN => n1791);
   U521 : CLKBUF_X1 port map( A => n5764, Z => n5850);
   U522 : OAI22_X1 port map( A1 => n7805, A2 => n5719, B1 => n5850, B2 => n5718
                           , ZN => n1790);
   U523 : CLKBUF_X1 port map( A => n5765, Z => n5851);
   U524 : OAI22_X1 port map( A1 => n7534, A2 => n5719, B1 => n5851, B2 => n5718
                           , ZN => n1789);
   U525 : CLKBUF_X1 port map( A => n5766, Z => n5852);
   U526 : OAI22_X1 port map( A1 => n7806, A2 => n5719, B1 => n5852, B2 => n5718
                           , ZN => n1788);
   U527 : CLKBUF_X1 port map( A => n5767, Z => n5853);
   U528 : OAI22_X1 port map( A1 => n7535, A2 => n5719, B1 => n5853, B2 => n5718
                           , ZN => n1787);
   U529 : CLKBUF_X1 port map( A => n5768, Z => n5854);
   U530 : OAI22_X1 port map( A1 => n7536, A2 => n5719, B1 => n5854, B2 => n5718
                           , ZN => n1786);
   U531 : CLKBUF_X1 port map( A => n5769, Z => n5855);
   U532 : OAI22_X1 port map( A1 => n7537, A2 => n5719, B1 => n5855, B2 => n5718
                           , ZN => n1785);
   U533 : OAI22_X1 port map( A1 => n7807, A2 => n5719, B1 => n5856, B2 => n5718
                           , ZN => n1784);
   U534 : CLKBUF_X1 port map( A => n5772, Z => n5858);
   U535 : OAI22_X1 port map( A1 => n7808, A2 => n5719, B1 => n5858, B2 => n5718
                           , ZN => n1783);
   U536 : NAND2_X1 port map( A1 => n5811, A2 => n5729, ZN => n5720);
   U537 : CLKBUF_X1 port map( A => n5720, Z => n5721);
   U538 : OAI22_X1 port map( A1 => n8023, A2 => n5722, B1 => n5788, B2 => n5721
                           , ZN => n1782);
   U539 : OAI22_X1 port map( A1 => n8024, A2 => n5722, B1 => n5740, B2 => n5720
                           , ZN => n1781);
   U540 : OAI22_X1 port map( A1 => n8270, A2 => n5722, B1 => n5741, B2 => n5721
                           , ZN => n1780);
   U541 : OAI22_X1 port map( A1 => n8271, A2 => n5722, B1 => n5742, B2 => n5720
                           , ZN => n1779);
   U542 : OAI22_X1 port map( A1 => n8025, A2 => n5722, B1 => n5743, B2 => n5721
                           , ZN => n1778);
   U543 : OAI22_X1 port map( A1 => n8026, A2 => n5722, B1 => n5744, B2 => n5720
                           , ZN => n1777);
   U544 : OAI22_X1 port map( A1 => n8272, A2 => n5722, B1 => n5745, B2 => n5721
                           , ZN => n1776);
   U545 : OAI22_X1 port map( A1 => n8027, A2 => n5722, B1 => n5746, B2 => n5720
                           , ZN => n1775);
   U546 : OAI22_X1 port map( A1 => n8273, A2 => n5722, B1 => n5747, B2 => n5721
                           , ZN => n1774);
   U547 : OAI22_X1 port map( A1 => n8274, A2 => n5722, B1 => n5748, B2 => n5720
                           , ZN => n1773);
   U548 : OAI22_X1 port map( A1 => n7538, A2 => n5722, B1 => n5749, B2 => n5720
                           , ZN => n1772);
   U549 : OAI22_X1 port map( A1 => n8275, A2 => n5722, B1 => n5750, B2 => n5721
                           , ZN => n1771);
   U550 : OAI22_X1 port map( A1 => n8276, A2 => n5722, B1 => n5751, B2 => n5720
                           , ZN => n1770);
   U551 : OAI22_X1 port map( A1 => n8028, A2 => n5722, B1 => n5752, B2 => n5721
                           , ZN => n1769);
   U552 : OAI22_X1 port map( A1 => n8277, A2 => n5722, B1 => n5753, B2 => n5720
                           , ZN => n1768);
   U553 : OAI22_X1 port map( A1 => n8029, A2 => n5722, B1 => n5754, B2 => n5721
                           , ZN => n1767);
   U554 : OAI22_X1 port map( A1 => n8030, A2 => n5722, B1 => n5755, B2 => n5720
                           , ZN => n1766);
   U555 : OAI22_X1 port map( A1 => n8278, A2 => n5722, B1 => n5756, B2 => n5720
                           , ZN => n1765);
   U556 : OAI22_X1 port map( A1 => n8031, A2 => n5722, B1 => n5757, B2 => n5720
                           , ZN => n1764);
   U557 : OAI22_X1 port map( A1 => n8032, A2 => n5722, B1 => n5758, B2 => n5720
                           , ZN => n1763);
   U558 : OAI22_X1 port map( A1 => n8033, A2 => n5722, B1 => n5759, B2 => n5720
                           , ZN => n1762);
   U559 : OAI22_X1 port map( A1 => n8279, A2 => n5722, B1 => n5760, B2 => n5720
                           , ZN => n1761);
   U560 : OAI22_X1 port map( A1 => n8034, A2 => n5722, B1 => n5762, B2 => n5720
                           , ZN => n1760);
   U561 : OAI22_X1 port map( A1 => n8035, A2 => n5722, B1 => n5763, B2 => n5721
                           , ZN => n1759);
   U562 : OAI22_X1 port map( A1 => n7539, A2 => n5722, B1 => n5764, B2 => n5721
                           , ZN => n1758);
   U563 : OAI22_X1 port map( A1 => n8280, A2 => n5722, B1 => n5765, B2 => n5721
                           , ZN => n1757);
   U564 : OAI22_X1 port map( A1 => n8036, A2 => n5722, B1 => n5766, B2 => n5721
                           , ZN => n1756);
   U565 : OAI22_X1 port map( A1 => n8281, A2 => n5722, B1 => n5767, B2 => n5721
                           , ZN => n1755);
   U566 : OAI22_X1 port map( A1 => n7540, A2 => n5722, B1 => n5768, B2 => n5721
                           , ZN => n1754);
   U567 : OAI22_X1 port map( A1 => n8282, A2 => n5722, B1 => n5769, B2 => n5721
                           , ZN => n1753);
   U568 : OAI22_X1 port map( A1 => n8283, A2 => n5722, B1 => n5770, B2 => n5721
                           , ZN => n1752);
   U569 : OAI22_X1 port map( A1 => n8284, A2 => n5722, B1 => n5772, B2 => n5721
                           , ZN => n1751);
   U570 : NAND2_X1 port map( A1 => n5815, A2 => n5729, ZN => n5723);
   U571 : CLKBUF_X1 port map( A => n5723, Z => n5724);
   U572 : OAI22_X1 port map( A1 => n7541, A2 => n5725, B1 => n5788, B2 => n5724
                           , ZN => n1750);
   U573 : OAI22_X1 port map( A1 => n8037, A2 => n5725, B1 => n5826, B2 => n5723
                           , ZN => n1749);
   U574 : OAI22_X1 port map( A1 => n8285, A2 => n5725, B1 => n5827, B2 => n5724
                           , ZN => n1748);
   U575 : OAI22_X1 port map( A1 => n8038, A2 => n5725, B1 => n5828, B2 => n5723
                           , ZN => n1747);
   U576 : OAI22_X1 port map( A1 => n8039, A2 => n5725, B1 => n5829, B2 => n5724
                           , ZN => n1746);
   U577 : OAI22_X1 port map( A1 => n8040, A2 => n5725, B1 => n5830, B2 => n5723
                           , ZN => n1745);
   U578 : OAI22_X1 port map( A1 => n7542, A2 => n5725, B1 => n5831, B2 => n5724
                           , ZN => n1744);
   U579 : OAI22_X1 port map( A1 => n7809, A2 => n5725, B1 => n5832, B2 => n5723
                           , ZN => n1743);
   U580 : OAI22_X1 port map( A1 => n8041, A2 => n5725, B1 => n5833, B2 => n5724
                           , ZN => n1742);
   U581 : OAI22_X1 port map( A1 => n7810, A2 => n5725, B1 => n5834, B2 => n5723
                           , ZN => n1741);
   U582 : OAI22_X1 port map( A1 => n8286, A2 => n5725, B1 => n5835, B2 => n5723
                           , ZN => n1740);
   U583 : OAI22_X1 port map( A1 => n7543, A2 => n5725, B1 => n5836, B2 => n5724
                           , ZN => n1739);
   U584 : OAI22_X1 port map( A1 => n8042, A2 => n5725, B1 => n5837, B2 => n5723
                           , ZN => n1738);
   U585 : OAI22_X1 port map( A1 => n8287, A2 => n5725, B1 => n5838, B2 => n5724
                           , ZN => n1737);
   U586 : OAI22_X1 port map( A1 => n8043, A2 => n5725, B1 => n5839, B2 => n5723
                           , ZN => n1736);
   U587 : OAI22_X1 port map( A1 => n8044, A2 => n5725, B1 => n5840, B2 => n5724
                           , ZN => n1735);
   U588 : OAI22_X1 port map( A1 => n8045, A2 => n5725, B1 => n5841, B2 => n5723
                           , ZN => n1734);
   U589 : OAI22_X1 port map( A1 => n8288, A2 => n5725, B1 => n5842, B2 => n5723
                           , ZN => n1733);
   U590 : OAI22_X1 port map( A1 => n7544, A2 => n5725, B1 => n5843, B2 => n5723
                           , ZN => n1732);
   U591 : OAI22_X1 port map( A1 => n8046, A2 => n5725, B1 => n5844, B2 => n5723
                           , ZN => n1731);
   U592 : OAI22_X1 port map( A1 => n8289, A2 => n5725, B1 => n5845, B2 => n5723
                           , ZN => n1730);
   U593 : OAI22_X1 port map( A1 => n7811, A2 => n5725, B1 => n5846, B2 => n5723
                           , ZN => n1729);
   U594 : OAI22_X1 port map( A1 => n7812, A2 => n5725, B1 => n5848, B2 => n5723
                           , ZN => n1728);
   U595 : OAI22_X1 port map( A1 => n8290, A2 => n5725, B1 => n5849, B2 => n5724
                           , ZN => n1727);
   U596 : OAI22_X1 port map( A1 => n8291, A2 => n5725, B1 => n5850, B2 => n5724
                           , ZN => n1726);
   U597 : OAI22_X1 port map( A1 => n8047, A2 => n5725, B1 => n5851, B2 => n5724
                           , ZN => n1725);
   U598 : OAI22_X1 port map( A1 => n8048, A2 => n5725, B1 => n5852, B2 => n5724
                           , ZN => n1724);
   U599 : OAI22_X1 port map( A1 => n8292, A2 => n5725, B1 => n5853, B2 => n5724
                           , ZN => n1723);
   U600 : OAI22_X1 port map( A1 => n8293, A2 => n5725, B1 => n5854, B2 => n5724
                           , ZN => n1722);
   U601 : OAI22_X1 port map( A1 => n7813, A2 => n5725, B1 => n5855, B2 => n5724
                           , ZN => n1721);
   U602 : OAI22_X1 port map( A1 => n7545, A2 => n5725, B1 => n5856, B2 => n5724
                           , ZN => n1720);
   U603 : OAI22_X1 port map( A1 => n8294, A2 => n5725, B1 => n5858, B2 => n5724
                           , ZN => n1719);
   U604 : NAND2_X1 port map( A1 => n5819, A2 => n5729, ZN => n5726);
   U605 : CLKBUF_X1 port map( A => n5726, Z => n5727);
   U606 : OAI22_X1 port map( A1 => n8049, A2 => n5728, B1 => n5788, B2 => n5727
                           , ZN => n1718);
   U607 : OAI22_X1 port map( A1 => n8295, A2 => n5728, B1 => n5740, B2 => n5726
                           , ZN => n1717);
   U608 : OAI22_X1 port map( A1 => n8050, A2 => n5728, B1 => n5741, B2 => n5727
                           , ZN => n1716);
   U609 : OAI22_X1 port map( A1 => n8296, A2 => n5728, B1 => n5742, B2 => n5726
                           , ZN => n1715);
   U610 : OAI22_X1 port map( A1 => n8051, A2 => n5728, B1 => n5743, B2 => n5727
                           , ZN => n1714);
   U611 : OAI22_X1 port map( A1 => n8052, A2 => n5728, B1 => n5744, B2 => n5726
                           , ZN => n1713);
   U612 : OAI22_X1 port map( A1 => n8053, A2 => n5728, B1 => n5745, B2 => n5727
                           , ZN => n1712);
   U613 : OAI22_X1 port map( A1 => n8054, A2 => n5728, B1 => n5746, B2 => n5726
                           , ZN => n1711);
   U614 : OAI22_X1 port map( A1 => n8297, A2 => n5728, B1 => n5747, B2 => n5727
                           , ZN => n1710);
   U615 : OAI22_X1 port map( A1 => n8298, A2 => n5728, B1 => n5748, B2 => n5726
                           , ZN => n1709);
   U616 : OAI22_X1 port map( A1 => n8055, A2 => n5728, B1 => n5749, B2 => n5726
                           , ZN => n1708);
   U617 : OAI22_X1 port map( A1 => n8299, A2 => n5728, B1 => n5750, B2 => n5727
                           , ZN => n1707);
   U618 : OAI22_X1 port map( A1 => n8056, A2 => n5728, B1 => n5751, B2 => n5726
                           , ZN => n1706);
   U619 : OAI22_X1 port map( A1 => n8300, A2 => n5728, B1 => n5752, B2 => n5727
                           , ZN => n1705);
   U620 : OAI22_X1 port map( A1 => n8301, A2 => n5728, B1 => n5753, B2 => n5726
                           , ZN => n1704);
   U621 : OAI22_X1 port map( A1 => n8302, A2 => n5728, B1 => n5754, B2 => n5727
                           , ZN => n1703);
   U622 : OAI22_X1 port map( A1 => n8303, A2 => n5728, B1 => n5755, B2 => n5726
                           , ZN => n1702);
   U623 : OAI22_X1 port map( A1 => n8057, A2 => n5728, B1 => n5756, B2 => n5726
                           , ZN => n1701);
   U624 : OAI22_X1 port map( A1 => n8058, A2 => n5728, B1 => n5757, B2 => n5726
                           , ZN => n1700);
   U625 : OAI22_X1 port map( A1 => n8304, A2 => n5728, B1 => n5758, B2 => n5726
                           , ZN => n1699);
   U626 : OAI22_X1 port map( A1 => n8059, A2 => n5728, B1 => n5759, B2 => n5726
                           , ZN => n1698);
   U627 : OAI22_X1 port map( A1 => n8060, A2 => n5728, B1 => n5760, B2 => n5726
                           , ZN => n1697);
   U628 : OAI22_X1 port map( A1 => n8305, A2 => n5728, B1 => n5762, B2 => n5726
                           , ZN => n1696);
   U629 : OAI22_X1 port map( A1 => n8306, A2 => n5728, B1 => n5763, B2 => n5727
                           , ZN => n1695);
   U630 : OAI22_X1 port map( A1 => n8061, A2 => n5728, B1 => n5764, B2 => n5727
                           , ZN => n1694);
   U631 : OAI22_X1 port map( A1 => n8307, A2 => n5728, B1 => n5765, B2 => n5727
                           , ZN => n1693);
   U632 : OAI22_X1 port map( A1 => n8308, A2 => n5728, B1 => n5766, B2 => n5727
                           , ZN => n1692);
   U633 : OAI22_X1 port map( A1 => n8062, A2 => n5728, B1 => n5767, B2 => n5727
                           , ZN => n1691);
   U634 : OAI22_X1 port map( A1 => n8063, A2 => n5728, B1 => n5768, B2 => n5727
                           , ZN => n1690);
   U635 : OAI22_X1 port map( A1 => n8309, A2 => n5728, B1 => n5769, B2 => n5727
                           , ZN => n1689);
   U636 : OAI22_X1 port map( A1 => n8310, A2 => n5728, B1 => n5770, B2 => n5727
                           , ZN => n1688);
   U637 : OAI22_X1 port map( A1 => n8064, A2 => n5728, B1 => n5772, B2 => n5727
                           , ZN => n1687);
   U638 : NAND2_X1 port map( A1 => n5824, A2 => n5729, ZN => n5730);
   U639 : OAI22_X1 port map( A1 => n8311, A2 => n5732, B1 => n5788, B2 => n5731
                           , ZN => n1686);
   U640 : OAI22_X1 port map( A1 => n7814, A2 => n5732, B1 => n5826, B2 => n5730
                           , ZN => n1685);
   U641 : OAI22_X1 port map( A1 => n7815, A2 => n5732, B1 => n5827, B2 => n5731
                           , ZN => n1684);
   U642 : OAI22_X1 port map( A1 => n7546, A2 => n5732, B1 => n5828, B2 => n5730
                           , ZN => n1683);
   U643 : OAI22_X1 port map( A1 => n7816, A2 => n5732, B1 => n5829, B2 => n5731
                           , ZN => n1682);
   U644 : OAI22_X1 port map( A1 => n8312, A2 => n5732, B1 => n5830, B2 => n5730
                           , ZN => n1681);
   U645 : OAI22_X1 port map( A1 => n8065, A2 => n5732, B1 => n5831, B2 => n5731
                           , ZN => n1680);
   U646 : OAI22_X1 port map( A1 => n7547, A2 => n5732, B1 => n5832, B2 => n5730
                           , ZN => n1679);
   U647 : OAI22_X1 port map( A1 => n7817, A2 => n5732, B1 => n5833, B2 => n5731
                           , ZN => n1678);
   U648 : OAI22_X1 port map( A1 => n7548, A2 => n5732, B1 => n5834, B2 => n5730
                           , ZN => n1677);
   U649 : OAI22_X1 port map( A1 => n8313, A2 => n5732, B1 => n5835, B2 => n5730
                           , ZN => n1676);
   U650 : OAI22_X1 port map( A1 => n8066, A2 => n5732, B1 => n5836, B2 => n5731
                           , ZN => n1675);
   U651 : OAI22_X1 port map( A1 => n7549, A2 => n5732, B1 => n5837, B2 => n5730
                           , ZN => n1674);
   U652 : OAI22_X1 port map( A1 => n7550, A2 => n5732, B1 => n5838, B2 => n5731
                           , ZN => n1673);
   U653 : OAI22_X1 port map( A1 => n8067, A2 => n5732, B1 => n5839, B2 => n5730
                           , ZN => n1672);
   U654 : OAI22_X1 port map( A1 => n7818, A2 => n5732, B1 => n5840, B2 => n5731
                           , ZN => n1671);
   U655 : OAI22_X1 port map( A1 => n8314, A2 => n5732, B1 => n5841, B2 => n5730
                           , ZN => n1670);
   U656 : OAI22_X1 port map( A1 => n8068, A2 => n5732, B1 => n5842, B2 => n5730
                           , ZN => n1669);
   U657 : OAI22_X1 port map( A1 => n8069, A2 => n5732, B1 => n5843, B2 => n5730
                           , ZN => n1668);
   U658 : OAI22_X1 port map( A1 => n7819, A2 => n5732, B1 => n5844, B2 => n5730
                           , ZN => n1667);
   U659 : OAI22_X1 port map( A1 => n7551, A2 => n5732, B1 => n5845, B2 => n5730
                           , ZN => n1666);
   U660 : OAI22_X1 port map( A1 => n8315, A2 => n5732, B1 => n5846, B2 => n5730
                           , ZN => n1665);
   U661 : OAI22_X1 port map( A1 => n8070, A2 => n5732, B1 => n5848, B2 => n5730
                           , ZN => n1664);
   U662 : OAI22_X1 port map( A1 => n7552, A2 => n5732, B1 => n5849, B2 => n5731
                           , ZN => n1663);
   U663 : OAI22_X1 port map( A1 => n8316, A2 => n5732, B1 => n5850, B2 => n5731
                           , ZN => n1662);
   U664 : OAI22_X1 port map( A1 => n7553, A2 => n5732, B1 => n5851, B2 => n5731
                           , ZN => n1661);
   U665 : OAI22_X1 port map( A1 => n8317, A2 => n5732, B1 => n5852, B2 => n5731
                           , ZN => n1660);
   U666 : OAI22_X1 port map( A1 => n8318, A2 => n5732, B1 => n5853, B2 => n5731
                           , ZN => n1659);
   U667 : OAI22_X1 port map( A1 => n8071, A2 => n5732, B1 => n5854, B2 => n5731
                           , ZN => n1658);
   U668 : OAI22_X1 port map( A1 => n7820, A2 => n5732, B1 => n5855, B2 => n5731
                           , ZN => n1657);
   U669 : OAI22_X1 port map( A1 => n8072, A2 => n5732, B1 => n5856, B2 => n5731
                           , ZN => n1656);
   U670 : OAI22_X1 port map( A1 => n7554, A2 => n5732, B1 => n5858, B2 => n5731
                           , ZN => n1655);
   U671 : NOR2_X1 port map( A1 => n5793, A2 => n5733, ZN => n5787);
   U672 : NAND2_X1 port map( A1 => n5794, A2 => n5787, ZN => n5734);
   U673 : CLKBUF_X1 port map( A => n5734, Z => n5735);
   U674 : OAI22_X1 port map( A1 => n7940, A2 => n5736, B1 => n5788, B2 => n5735
                           , ZN => n1654);
   U675 : OAI22_X1 port map( A1 => n8073, A2 => n5736, B1 => n5740, B2 => n5734
                           , ZN => n1653);
   U676 : OAI22_X1 port map( A1 => n8319, A2 => n5736, B1 => n5741, B2 => n5735
                           , ZN => n1652);
   U677 : OAI22_X1 port map( A1 => n8320, A2 => n5736, B1 => n5742, B2 => n5734
                           , ZN => n1651);
   U678 : OAI22_X1 port map( A1 => n7555, A2 => n5736, B1 => n5743, B2 => n5735
                           , ZN => n1650);
   U679 : OAI22_X1 port map( A1 => n7821, A2 => n5736, B1 => n5744, B2 => n5734
                           , ZN => n1649);
   U680 : OAI22_X1 port map( A1 => n8074, A2 => n5736, B1 => n5745, B2 => n5735
                           , ZN => n1648);
   U681 : OAI22_X1 port map( A1 => n7556, A2 => n5736, B1 => n5746, B2 => n5734
                           , ZN => n1647);
   U682 : OAI22_X1 port map( A1 => n8321, A2 => n5736, B1 => n5747, B2 => n5735
                           , ZN => n1646);
   U683 : OAI22_X1 port map( A1 => n8075, A2 => n5736, B1 => n5748, B2 => n5734
                           , ZN => n1645);
   U684 : OAI22_X1 port map( A1 => n8322, A2 => n5736, B1 => n5749, B2 => n5734
                           , ZN => n1644);
   U685 : OAI22_X1 port map( A1 => n7822, A2 => n5736, B1 => n5750, B2 => n5735
                           , ZN => n1643);
   U686 : OAI22_X1 port map( A1 => n8323, A2 => n5736, B1 => n5751, B2 => n5734
                           , ZN => n1642);
   U687 : OAI22_X1 port map( A1 => n8324, A2 => n5736, B1 => n5752, B2 => n5735
                           , ZN => n1641);
   U688 : OAI22_X1 port map( A1 => n7557, A2 => n5736, B1 => n5753, B2 => n5734
                           , ZN => n1640);
   U689 : OAI22_X1 port map( A1 => n7823, A2 => n5736, B1 => n5754, B2 => n5735
                           , ZN => n1639);
   U690 : OAI22_X1 port map( A1 => n7824, A2 => n5736, B1 => n5755, B2 => n5734
                           , ZN => n1638);
   U691 : OAI22_X1 port map( A1 => n7825, A2 => n5736, B1 => n5756, B2 => n5734
                           , ZN => n1637);
   U692 : OAI22_X1 port map( A1 => n8325, A2 => n5736, B1 => n5757, B2 => n5734
                           , ZN => n1636);
   U693 : OAI22_X1 port map( A1 => n8326, A2 => n5736, B1 => n5758, B2 => n5734
                           , ZN => n1635);
   U694 : OAI22_X1 port map( A1 => n7826, A2 => n5736, B1 => n5759, B2 => n5734
                           , ZN => n1634);
   U695 : OAI22_X1 port map( A1 => n7827, A2 => n5736, B1 => n5760, B2 => n5734
                           , ZN => n1633);
   U696 : OAI22_X1 port map( A1 => n7558, A2 => n5736, B1 => n5762, B2 => n5734
                           , ZN => n1632);
   U697 : OAI22_X1 port map( A1 => n8076, A2 => n5736, B1 => n5763, B2 => n5735
                           , ZN => n1631);
   U698 : OAI22_X1 port map( A1 => n7828, A2 => n5736, B1 => n5764, B2 => n5735
                           , ZN => n1630);
   U699 : OAI22_X1 port map( A1 => n7829, A2 => n5736, B1 => n5765, B2 => n5735
                           , ZN => n1629);
   U700 : OAI22_X1 port map( A1 => n7559, A2 => n5736, B1 => n5766, B2 => n5735
                           , ZN => n1628);
   U701 : OAI22_X1 port map( A1 => n7830, A2 => n5736, B1 => n5767, B2 => n5735
                           , ZN => n1627);
   U702 : OAI22_X1 port map( A1 => n7831, A2 => n5736, B1 => n5768, B2 => n5735
                           , ZN => n1626);
   U703 : OAI22_X1 port map( A1 => n7560, A2 => n5736, B1 => n5769, B2 => n5735
                           , ZN => n1625);
   U704 : OAI22_X1 port map( A1 => n8077, A2 => n5736, B1 => n5770, B2 => n5735
                           , ZN => n1624);
   U705 : OAI22_X1 port map( A1 => n7561, A2 => n5736, B1 => n5772, B2 => n5735
                           , ZN => n1623);
   U706 : NAND2_X1 port map( A1 => n5798, A2 => n5787, ZN => n5737);
   U707 : CLKBUF_X1 port map( A => n5737, Z => n5738);
   U708 : OAI22_X1 port map( A1 => n7684, A2 => n5739, B1 => n5788, B2 => n5738
                           , ZN => n1622);
   U709 : OAI22_X1 port map( A1 => n7832, A2 => n5739, B1 => n5826, B2 => n5737
                           , ZN => n1621);
   U710 : OAI22_X1 port map( A1 => n7833, A2 => n5739, B1 => n5827, B2 => n5738
                           , ZN => n1620);
   U711 : OAI22_X1 port map( A1 => n7562, A2 => n5739, B1 => n5828, B2 => n5737
                           , ZN => n1619);
   U712 : OAI22_X1 port map( A1 => n8078, A2 => n5739, B1 => n5829, B2 => n5738
                           , ZN => n1618);
   U713 : OAI22_X1 port map( A1 => n8079, A2 => n5739, B1 => n5830, B2 => n5737
                           , ZN => n1617);
   U714 : OAI22_X1 port map( A1 => n7563, A2 => n5739, B1 => n5831, B2 => n5738
                           , ZN => n1616);
   U715 : OAI22_X1 port map( A1 => n8327, A2 => n5739, B1 => n5832, B2 => n5737
                           , ZN => n1615);
   U716 : OAI22_X1 port map( A1 => n7564, A2 => n5739, B1 => n5833, B2 => n5738
                           , ZN => n1614);
   U717 : OAI22_X1 port map( A1 => n7565, A2 => n5739, B1 => n5834, B2 => n5737
                           , ZN => n1613);
   U718 : OAI22_X1 port map( A1 => n7566, A2 => n5739, B1 => n5835, B2 => n5737
                           , ZN => n1612);
   U719 : OAI22_X1 port map( A1 => n7567, A2 => n5739, B1 => n5836, B2 => n5738
                           , ZN => n1611);
   U720 : OAI22_X1 port map( A1 => n7568, A2 => n5739, B1 => n5837, B2 => n5737
                           , ZN => n1610);
   U721 : OAI22_X1 port map( A1 => n7569, A2 => n5739, B1 => n5838, B2 => n5738
                           , ZN => n1609);
   U722 : OAI22_X1 port map( A1 => n7570, A2 => n5739, B1 => n5839, B2 => n5737
                           , ZN => n1608);
   U723 : OAI22_X1 port map( A1 => n7834, A2 => n5739, B1 => n5840, B2 => n5738
                           , ZN => n1607);
   U724 : OAI22_X1 port map( A1 => n7835, A2 => n5739, B1 => n5841, B2 => n5737
                           , ZN => n1606);
   U725 : OAI22_X1 port map( A1 => n8328, A2 => n5739, B1 => n5842, B2 => n5737
                           , ZN => n1605);
   U726 : OAI22_X1 port map( A1 => n7571, A2 => n5739, B1 => n5843, B2 => n5737
                           , ZN => n1604);
   U727 : OAI22_X1 port map( A1 => n7836, A2 => n5739, B1 => n5844, B2 => n5737
                           , ZN => n1603);
   U728 : OAI22_X1 port map( A1 => n7572, A2 => n5739, B1 => n5845, B2 => n5737
                           , ZN => n1602);
   U729 : OAI22_X1 port map( A1 => n7573, A2 => n5739, B1 => n5846, B2 => n5737
                           , ZN => n1601);
   U730 : OAI22_X1 port map( A1 => n8329, A2 => n5739, B1 => n5848, B2 => n5737
                           , ZN => n1600);
   U731 : OAI22_X1 port map( A1 => n7574, A2 => n5739, B1 => n5849, B2 => n5738
                           , ZN => n1599);
   U732 : OAI22_X1 port map( A1 => n8080, A2 => n5739, B1 => n5850, B2 => n5738
                           , ZN => n1598);
   U733 : OAI22_X1 port map( A1 => n7837, A2 => n5739, B1 => n5851, B2 => n5738
                           , ZN => n1597);
   U734 : OAI22_X1 port map( A1 => n7575, A2 => n5739, B1 => n5852, B2 => n5738
                           , ZN => n1596);
   U735 : OAI22_X1 port map( A1 => n8081, A2 => n5739, B1 => n5853, B2 => n5738
                           , ZN => n1595);
   U736 : OAI22_X1 port map( A1 => n7576, A2 => n5739, B1 => n5854, B2 => n5738
                           , ZN => n1594);
   U737 : OAI22_X1 port map( A1 => n7577, A2 => n5739, B1 => n5855, B2 => n5738
                           , ZN => n1593);
   U738 : OAI22_X1 port map( A1 => n7578, A2 => n5739, B1 => n5856, B2 => n5738
                           , ZN => n1592);
   U739 : OAI22_X1 port map( A1 => n7838, A2 => n5739, B1 => n5858, B2 => n5738
                           , ZN => n1591);
   U740 : NAND2_X1 port map( A1 => n5802, A2 => n5787, ZN => n5761);
   U741 : CLKBUF_X1 port map( A => n5761, Z => n5771);
   U742 : OAI22_X1 port map( A1 => n7685, A2 => n5773, B1 => n5788, B2 => n5771
                           , ZN => n1590);
   U743 : OAI22_X1 port map( A1 => n8330, A2 => n5773, B1 => n5740, B2 => n5761
                           , ZN => n1589);
   U744 : OAI22_X1 port map( A1 => n8331, A2 => n5773, B1 => n5741, B2 => n5771
                           , ZN => n1588);
   U745 : OAI22_X1 port map( A1 => n7839, A2 => n5773, B1 => n5742, B2 => n5761
                           , ZN => n1587);
   U746 : OAI22_X1 port map( A1 => n8082, A2 => n5773, B1 => n5743, B2 => n5771
                           , ZN => n1586);
   U747 : OAI22_X1 port map( A1 => n7579, A2 => n5773, B1 => n5744, B2 => n5761
                           , ZN => n1585);
   U748 : OAI22_X1 port map( A1 => n7840, A2 => n5773, B1 => n5745, B2 => n5771
                           , ZN => n1584);
   U749 : OAI22_X1 port map( A1 => n8332, A2 => n5773, B1 => n5746, B2 => n5761
                           , ZN => n1583);
   U750 : OAI22_X1 port map( A1 => n7580, A2 => n5773, B1 => n5747, B2 => n5771
                           , ZN => n1582);
   U751 : OAI22_X1 port map( A1 => n7581, A2 => n5773, B1 => n5748, B2 => n5761
                           , ZN => n1581);
   U752 : OAI22_X1 port map( A1 => n8083, A2 => n5773, B1 => n5749, B2 => n5761
                           , ZN => n1580);
   U753 : OAI22_X1 port map( A1 => n7582, A2 => n5773, B1 => n5750, B2 => n5771
                           , ZN => n1579);
   U754 : OAI22_X1 port map( A1 => n7841, A2 => n5773, B1 => n5751, B2 => n5761
                           , ZN => n1578);
   U755 : OAI22_X1 port map( A1 => n7583, A2 => n5773, B1 => n5752, B2 => n5771
                           , ZN => n1577);
   U756 : OAI22_X1 port map( A1 => n8084, A2 => n5773, B1 => n5753, B2 => n5761
                           , ZN => n1576);
   U757 : OAI22_X1 port map( A1 => n8085, A2 => n5773, B1 => n5754, B2 => n5771
                           , ZN => n1575);
   U758 : OAI22_X1 port map( A1 => n8086, A2 => n5773, B1 => n5755, B2 => n5761
                           , ZN => n1574);
   U759 : OAI22_X1 port map( A1 => n8333, A2 => n5773, B1 => n5756, B2 => n5761
                           , ZN => n1573);
   U760 : OAI22_X1 port map( A1 => n8087, A2 => n5773, B1 => n5757, B2 => n5761
                           , ZN => n1572);
   U761 : OAI22_X1 port map( A1 => n8334, A2 => n5773, B1 => n5758, B2 => n5761
                           , ZN => n1571);
   U762 : OAI22_X1 port map( A1 => n8335, A2 => n5773, B1 => n5759, B2 => n5761
                           , ZN => n1570);
   U763 : OAI22_X1 port map( A1 => n8336, A2 => n5773, B1 => n5760, B2 => n5761
                           , ZN => n1569);
   U764 : OAI22_X1 port map( A1 => n8337, A2 => n5773, B1 => n5762, B2 => n5761
                           , ZN => n1568);
   U765 : OAI22_X1 port map( A1 => n8088, A2 => n5773, B1 => n5763, B2 => n5771
                           , ZN => n1567);
   U766 : OAI22_X1 port map( A1 => n7842, A2 => n5773, B1 => n5764, B2 => n5771
                           , ZN => n1566);
   U767 : OAI22_X1 port map( A1 => n8089, A2 => n5773, B1 => n5765, B2 => n5771
                           , ZN => n1565);
   U768 : OAI22_X1 port map( A1 => n8090, A2 => n5773, B1 => n5766, B2 => n5771
                           , ZN => n1564);
   U769 : OAI22_X1 port map( A1 => n7584, A2 => n5773, B1 => n5767, B2 => n5771
                           , ZN => n1563);
   U770 : OAI22_X1 port map( A1 => n8091, A2 => n5773, B1 => n5768, B2 => n5771
                           , ZN => n1562);
   U771 : OAI22_X1 port map( A1 => n7843, A2 => n5773, B1 => n5769, B2 => n5771
                           , ZN => n1561);
   U772 : OAI22_X1 port map( A1 => n8338, A2 => n5773, B1 => n5770, B2 => n5771
                           , ZN => n1560);
   U773 : OAI22_X1 port map( A1 => n7844, A2 => n5773, B1 => n5772, B2 => n5771
                           , ZN => n1559);
   U774 : NAND2_X1 port map( A1 => n5807, A2 => n5787, ZN => n5774);
   U775 : CLKBUF_X1 port map( A => n5774, Z => n5775);
   U776 : OAI22_X1 port map( A1 => n7424, A2 => n5776, B1 => n5788, B2 => n5775
                           , ZN => n1558);
   U777 : OAI22_X1 port map( A1 => n7585, A2 => n5776, B1 => n5826, B2 => n5774
                           , ZN => n1557);
   U778 : OAI22_X1 port map( A1 => n7845, A2 => n5776, B1 => n5827, B2 => n5775
                           , ZN => n1556);
   U779 : OAI22_X1 port map( A1 => n7846, A2 => n5776, B1 => n5828, B2 => n5774
                           , ZN => n1555);
   U780 : OAI22_X1 port map( A1 => n8339, A2 => n5776, B1 => n5829, B2 => n5775
                           , ZN => n1554);
   U781 : OAI22_X1 port map( A1 => n7847, A2 => n5776, B1 => n5830, B2 => n5774
                           , ZN => n1553);
   U782 : OAI22_X1 port map( A1 => n8340, A2 => n5776, B1 => n5831, B2 => n5775
                           , ZN => n1552);
   U783 : OAI22_X1 port map( A1 => n8341, A2 => n5776, B1 => n5832, B2 => n5774
                           , ZN => n1551);
   U784 : OAI22_X1 port map( A1 => n8342, A2 => n5776, B1 => n5833, B2 => n5775
                           , ZN => n1550);
   U785 : OAI22_X1 port map( A1 => n7848, A2 => n5776, B1 => n5834, B2 => n5774
                           , ZN => n1549);
   U786 : OAI22_X1 port map( A1 => n8092, A2 => n5776, B1 => n5835, B2 => n5774
                           , ZN => n1548);
   U787 : OAI22_X1 port map( A1 => n8093, A2 => n5776, B1 => n5836, B2 => n5775
                           , ZN => n1547);
   U788 : OAI22_X1 port map( A1 => n7586, A2 => n5776, B1 => n5837, B2 => n5774
                           , ZN => n1546);
   U789 : OAI22_X1 port map( A1 => n8343, A2 => n5776, B1 => n5838, B2 => n5775
                           , ZN => n1545);
   U790 : OAI22_X1 port map( A1 => n8094, A2 => n5776, B1 => n5839, B2 => n5774
                           , ZN => n1544);
   U791 : OAI22_X1 port map( A1 => n8095, A2 => n5776, B1 => n5840, B2 => n5775
                           , ZN => n1543);
   U792 : OAI22_X1 port map( A1 => n7587, A2 => n5776, B1 => n5841, B2 => n5774
                           , ZN => n1542);
   U793 : OAI22_X1 port map( A1 => n8096, A2 => n5776, B1 => n5842, B2 => n5774
                           , ZN => n1541);
   U794 : OAI22_X1 port map( A1 => n8344, A2 => n5776, B1 => n5843, B2 => n5774
                           , ZN => n1540);
   U795 : OAI22_X1 port map( A1 => n7588, A2 => n5776, B1 => n5844, B2 => n5774
                           , ZN => n1539);
   U796 : OAI22_X1 port map( A1 => n7589, A2 => n5776, B1 => n5845, B2 => n5774
                           , ZN => n1538);
   U797 : OAI22_X1 port map( A1 => n7590, A2 => n5776, B1 => n5846, B2 => n5774
                           , ZN => n1537);
   U798 : OAI22_X1 port map( A1 => n7849, A2 => n5776, B1 => n5848, B2 => n5774
                           , ZN => n1536);
   U799 : OAI22_X1 port map( A1 => n8345, A2 => n5776, B1 => n5849, B2 => n5775
                           , ZN => n1535);
   U800 : OAI22_X1 port map( A1 => n7591, A2 => n5776, B1 => n5850, B2 => n5775
                           , ZN => n1534);
   U801 : OAI22_X1 port map( A1 => n7592, A2 => n5776, B1 => n5851, B2 => n5775
                           , ZN => n1533);
   U802 : OAI22_X1 port map( A1 => n7593, A2 => n5776, B1 => n5852, B2 => n5775
                           , ZN => n1532);
   U803 : OAI22_X1 port map( A1 => n8346, A2 => n5776, B1 => n5853, B2 => n5775
                           , ZN => n1531);
   U804 : OAI22_X1 port map( A1 => n8347, A2 => n5776, B1 => n5854, B2 => n5775
                           , ZN => n1530);
   U805 : OAI22_X1 port map( A1 => n8348, A2 => n5776, B1 => n5855, B2 => n5775
                           , ZN => n1529);
   U806 : OAI22_X1 port map( A1 => n8097, A2 => n5776, B1 => n5856, B2 => n5775
                           , ZN => n1528);
   U807 : OAI22_X1 port map( A1 => n8349, A2 => n5776, B1 => n5858, B2 => n5775
                           , ZN => n1527);
   U808 : NAND2_X1 port map( A1 => n5811, A2 => n5787, ZN => n5777);
   U809 : CLKBUF_X1 port map( A => n5777, Z => n5778);
   U810 : OAI22_X1 port map( A1 => n7686, A2 => n5779, B1 => n5788, B2 => n5778
                           , ZN => n1526);
   U811 : OAI22_X1 port map( A1 => n8098, A2 => n5779, B1 => n5826, B2 => n5777
                           , ZN => n1525);
   U812 : OAI22_X1 port map( A1 => n8099, A2 => n5779, B1 => n5827, B2 => n5778
                           , ZN => n1524);
   U813 : OAI22_X1 port map( A1 => n7594, A2 => n5779, B1 => n5828, B2 => n5777
                           , ZN => n1523);
   U814 : OAI22_X1 port map( A1 => n7850, A2 => n5779, B1 => n5829, B2 => n5778
                           , ZN => n1522);
   U815 : OAI22_X1 port map( A1 => n8350, A2 => n5779, B1 => n5830, B2 => n5777
                           , ZN => n1521);
   U816 : OAI22_X1 port map( A1 => n8351, A2 => n5779, B1 => n5831, B2 => n5778
                           , ZN => n1520);
   U817 : OAI22_X1 port map( A1 => n8100, A2 => n5779, B1 => n5832, B2 => n5777
                           , ZN => n1519);
   U818 : OAI22_X1 port map( A1 => n8101, A2 => n5779, B1 => n5833, B2 => n5778
                           , ZN => n1518);
   U819 : OAI22_X1 port map( A1 => n8102, A2 => n5779, B1 => n5834, B2 => n5777
                           , ZN => n1517);
   U820 : OAI22_X1 port map( A1 => n8103, A2 => n5779, B1 => n5835, B2 => n5777
                           , ZN => n1516);
   U821 : OAI22_X1 port map( A1 => n8104, A2 => n5779, B1 => n5836, B2 => n5778
                           , ZN => n1515);
   U822 : OAI22_X1 port map( A1 => n8352, A2 => n5779, B1 => n5837, B2 => n5777
                           , ZN => n1514);
   U823 : OAI22_X1 port map( A1 => n8105, A2 => n5779, B1 => n5838, B2 => n5778
                           , ZN => n1513);
   U824 : OAI22_X1 port map( A1 => n8353, A2 => n5779, B1 => n5839, B2 => n5777
                           , ZN => n1512);
   U825 : OAI22_X1 port map( A1 => n8354, A2 => n5779, B1 => n5840, B2 => n5778
                           , ZN => n1511);
   U826 : OAI22_X1 port map( A1 => n8106, A2 => n5779, B1 => n5841, B2 => n5777
                           , ZN => n1510);
   U827 : OAI22_X1 port map( A1 => n8355, A2 => n5779, B1 => n5842, B2 => n5777
                           , ZN => n1509);
   U828 : OAI22_X1 port map( A1 => n8356, A2 => n5779, B1 => n5843, B2 => n5777
                           , ZN => n1508);
   U829 : OAI22_X1 port map( A1 => n8107, A2 => n5779, B1 => n5844, B2 => n5777
                           , ZN => n1507);
   U830 : OAI22_X1 port map( A1 => n8108, A2 => n5779, B1 => n5845, B2 => n5777
                           , ZN => n1506);
   U831 : OAI22_X1 port map( A1 => n8357, A2 => n5779, B1 => n5846, B2 => n5777
                           , ZN => n1505);
   U832 : OAI22_X1 port map( A1 => n8109, A2 => n5779, B1 => n5848, B2 => n5777
                           , ZN => n1504);
   U833 : OAI22_X1 port map( A1 => n8358, A2 => n5779, B1 => n5849, B2 => n5778
                           , ZN => n1503);
   U834 : OAI22_X1 port map( A1 => n8110, A2 => n5779, B1 => n5850, B2 => n5778
                           , ZN => n1502);
   U835 : OAI22_X1 port map( A1 => n8359, A2 => n5779, B1 => n5851, B2 => n5778
                           , ZN => n1501);
   U836 : OAI22_X1 port map( A1 => n8360, A2 => n5779, B1 => n5852, B2 => n5778
                           , ZN => n1500);
   U837 : OAI22_X1 port map( A1 => n8361, A2 => n5779, B1 => n5853, B2 => n5778
                           , ZN => n1499);
   U838 : OAI22_X1 port map( A1 => n8362, A2 => n5779, B1 => n5854, B2 => n5778
                           , ZN => n1498);
   U839 : OAI22_X1 port map( A1 => n8111, A2 => n5779, B1 => n5855, B2 => n5778
                           , ZN => n1497);
   U840 : OAI22_X1 port map( A1 => n8363, A2 => n5779, B1 => n5856, B2 => n5778
                           , ZN => n1496);
   U841 : OAI22_X1 port map( A1 => n8364, A2 => n5779, B1 => n5858, B2 => n5778
                           , ZN => n1495);
   U842 : NAND2_X1 port map( A1 => n5815, A2 => n5787, ZN => n5780);
   U843 : CLKBUF_X1 port map( A => n5780, Z => n5781);
   U844 : OAI22_X1 port map( A1 => n7941, A2 => n5782, B1 => n5788, B2 => n5781
                           , ZN => n1494);
   U845 : OAI22_X1 port map( A1 => n8112, A2 => n5782, B1 => n5826, B2 => n5780
                           , ZN => n1493);
   U846 : OAI22_X1 port map( A1 => n8113, A2 => n5782, B1 => n5827, B2 => n5781
                           , ZN => n1492);
   U847 : OAI22_X1 port map( A1 => n8365, A2 => n5782, B1 => n5828, B2 => n5780
                           , ZN => n1491);
   U848 : OAI22_X1 port map( A1 => n8114, A2 => n5782, B1 => n5829, B2 => n5781
                           , ZN => n1490);
   U849 : OAI22_X1 port map( A1 => n8115, A2 => n5782, B1 => n5830, B2 => n5780
                           , ZN => n1489);
   U850 : OAI22_X1 port map( A1 => n8366, A2 => n5782, B1 => n5831, B2 => n5781
                           , ZN => n1488);
   U851 : OAI22_X1 port map( A1 => n8116, A2 => n5782, B1 => n5832, B2 => n5780
                           , ZN => n1487);
   U852 : OAI22_X1 port map( A1 => n8117, A2 => n5782, B1 => n5833, B2 => n5781
                           , ZN => n1486);
   U853 : OAI22_X1 port map( A1 => n8118, A2 => n5782, B1 => n5834, B2 => n5780
                           , ZN => n1485);
   U854 : OAI22_X1 port map( A1 => n7851, A2 => n5782, B1 => n5835, B2 => n5780
                           , ZN => n1484);
   U855 : OAI22_X1 port map( A1 => n8367, A2 => n5782, B1 => n5836, B2 => n5781
                           , ZN => n1483);
   U856 : OAI22_X1 port map( A1 => n8119, A2 => n5782, B1 => n5837, B2 => n5780
                           , ZN => n1482);
   U857 : OAI22_X1 port map( A1 => n8368, A2 => n5782, B1 => n5838, B2 => n5781
                           , ZN => n1481);
   U858 : OAI22_X1 port map( A1 => n8369, A2 => n5782, B1 => n5839, B2 => n5780
                           , ZN => n1480);
   U859 : OAI22_X1 port map( A1 => n8370, A2 => n5782, B1 => n5840, B2 => n5781
                           , ZN => n1479);
   U860 : OAI22_X1 port map( A1 => n8120, A2 => n5782, B1 => n5841, B2 => n5780
                           , ZN => n1478);
   U861 : OAI22_X1 port map( A1 => n8371, A2 => n5782, B1 => n5842, B2 => n5780
                           , ZN => n1477);
   U862 : OAI22_X1 port map( A1 => n8372, A2 => n5782, B1 => n5843, B2 => n5780
                           , ZN => n1476);
   U863 : OAI22_X1 port map( A1 => n8121, A2 => n5782, B1 => n5844, B2 => n5780
                           , ZN => n1475);
   U864 : OAI22_X1 port map( A1 => n8373, A2 => n5782, B1 => n5845, B2 => n5780
                           , ZN => n1474);
   U865 : OAI22_X1 port map( A1 => n8122, A2 => n5782, B1 => n5846, B2 => n5780
                           , ZN => n1473);
   U866 : OAI22_X1 port map( A1 => n8374, A2 => n5782, B1 => n5848, B2 => n5780
                           , ZN => n1472);
   U867 : OAI22_X1 port map( A1 => n8375, A2 => n5782, B1 => n5849, B2 => n5781
                           , ZN => n1471);
   U868 : OAI22_X1 port map( A1 => n8376, A2 => n5782, B1 => n5850, B2 => n5781
                           , ZN => n1470);
   U869 : OAI22_X1 port map( A1 => n8377, A2 => n5782, B1 => n5851, B2 => n5781
                           , ZN => n1469);
   U870 : OAI22_X1 port map( A1 => n8378, A2 => n5782, B1 => n5852, B2 => n5781
                           , ZN => n1468);
   U871 : OAI22_X1 port map( A1 => n8123, A2 => n5782, B1 => n5853, B2 => n5781
                           , ZN => n1467);
   U872 : OAI22_X1 port map( A1 => n8379, A2 => n5782, B1 => n5854, B2 => n5781
                           , ZN => n1466);
   U873 : OAI22_X1 port map( A1 => n8124, A2 => n5782, B1 => n5855, B2 => n5781
                           , ZN => n1465);
   U874 : OAI22_X1 port map( A1 => n8380, A2 => n5782, B1 => n5856, B2 => n5781
                           , ZN => n1464);
   U875 : OAI22_X1 port map( A1 => n8125, A2 => n5782, B1 => n5858, B2 => n5781
                           , ZN => n1463);
   U876 : NAND2_X1 port map( A1 => n5819, A2 => n5787, ZN => n5783);
   U877 : CLKBUF_X1 port map( A => n5786, Z => n5784);
   U878 : CLKBUF_X1 port map( A => n5783, Z => n5785);
   U879 : OAI22_X1 port map( A1 => n7942, A2 => n5784, B1 => n5788, B2 => n5785
                           , ZN => n1462);
   U880 : OAI22_X1 port map( A1 => n8381, A2 => n5786, B1 => n5826, B2 => n5783
                           , ZN => n1461);
   U881 : OAI22_X1 port map( A1 => n8382, A2 => n5784, B1 => n5827, B2 => n5785
                           , ZN => n1460);
   U882 : OAI22_X1 port map( A1 => n8126, A2 => n5786, B1 => n5828, B2 => n5783
                           , ZN => n1459);
   U883 : OAI22_X1 port map( A1 => n8383, A2 => n5784, B1 => n5829, B2 => n5785
                           , ZN => n1458);
   U884 : OAI22_X1 port map( A1 => n8127, A2 => n5786, B1 => n5830, B2 => n5783
                           , ZN => n1457);
   U885 : OAI22_X1 port map( A1 => n8384, A2 => n5784, B1 => n5831, B2 => n5785
                           , ZN => n1456);
   U886 : OAI22_X1 port map( A1 => n8128, A2 => n5786, B1 => n5832, B2 => n5783
                           , ZN => n1455);
   U887 : OAI22_X1 port map( A1 => n8129, A2 => n5784, B1 => n5833, B2 => n5785
                           , ZN => n1454);
   U888 : OAI22_X1 port map( A1 => n8385, A2 => n5786, B1 => n5834, B2 => n5783
                           , ZN => n1453);
   U889 : OAI22_X1 port map( A1 => n8386, A2 => n5786, B1 => n5835, B2 => n5783
                           , ZN => n1452);
   U890 : OAI22_X1 port map( A1 => n8387, A2 => n5786, B1 => n5836, B2 => n5785
                           , ZN => n1451);
   U891 : OAI22_X1 port map( A1 => n8388, A2 => n5784, B1 => n5837, B2 => n5783
                           , ZN => n1450);
   U892 : OAI22_X1 port map( A1 => n8130, A2 => n5784, B1 => n5838, B2 => n5785
                           , ZN => n1449);
   U893 : OAI22_X1 port map( A1 => n8389, A2 => n5784, B1 => n5839, B2 => n5783
                           , ZN => n1448);
   U894 : OAI22_X1 port map( A1 => n8131, A2 => n5784, B1 => n5840, B2 => n5785
                           , ZN => n1447);
   U895 : OAI22_X1 port map( A1 => n8132, A2 => n5784, B1 => n5841, B2 => n5783
                           , ZN => n1446);
   U896 : OAI22_X1 port map( A1 => n8390, A2 => n5784, B1 => n5842, B2 => n5783
                           , ZN => n1445);
   U897 : OAI22_X1 port map( A1 => n8133, A2 => n5784, B1 => n5843, B2 => n5783
                           , ZN => n1444);
   U898 : OAI22_X1 port map( A1 => n8134, A2 => n5784, B1 => n5844, B2 => n5783
                           , ZN => n1443);
   U899 : OAI22_X1 port map( A1 => n8135, A2 => n5784, B1 => n5845, B2 => n5783
                           , ZN => n1442);
   U900 : OAI22_X1 port map( A1 => n8136, A2 => n5784, B1 => n5846, B2 => n5783
                           , ZN => n1441);
   U901 : OAI22_X1 port map( A1 => n8137, A2 => n5784, B1 => n5848, B2 => n5783
                           , ZN => n1440);
   U902 : OAI22_X1 port map( A1 => n8138, A2 => n5784, B1 => n5849, B2 => n5785
                           , ZN => n1439);
   U903 : OAI22_X1 port map( A1 => n8391, A2 => n5786, B1 => n5850, B2 => n5785
                           , ZN => n1438);
   U904 : OAI22_X1 port map( A1 => n8392, A2 => n5786, B1 => n5851, B2 => n5785
                           , ZN => n1437);
   U905 : OAI22_X1 port map( A1 => n8393, A2 => n5786, B1 => n5852, B2 => n5785
                           , ZN => n1436);
   U906 : OAI22_X1 port map( A1 => n8394, A2 => n5786, B1 => n5853, B2 => n5785
                           , ZN => n1435);
   U907 : OAI22_X1 port map( A1 => n8139, A2 => n5786, B1 => n5854, B2 => n5785
                           , ZN => n1434);
   U908 : OAI22_X1 port map( A1 => n8395, A2 => n5786, B1 => n5855, B2 => n5785
                           , ZN => n1433);
   U909 : OAI22_X1 port map( A1 => n8140, A2 => n5786, B1 => n5856, B2 => n5785
                           , ZN => n1432);
   U910 : OAI22_X1 port map( A1 => n8141, A2 => n5786, B1 => n5858, B2 => n5785
                           , ZN => n1431);
   U911 : NAND2_X1 port map( A1 => n5824, A2 => n5787, ZN => n5789);
   U912 : CLKBUF_X1 port map( A => n5789, Z => n5790);
   U913 : OAI22_X1 port map( A1 => n7687, A2 => n5791, B1 => n5788, B2 => n5790
                           , ZN => n1430);
   U914 : OAI22_X1 port map( A1 => n7852, A2 => n5791, B1 => n5826, B2 => n5789
                           , ZN => n1429);
   U915 : OAI22_X1 port map( A1 => n7853, A2 => n5791, B1 => n5827, B2 => n5790
                           , ZN => n1428);
   U916 : OAI22_X1 port map( A1 => n8142, A2 => n5791, B1 => n5828, B2 => n5789
                           , ZN => n1427);
   U917 : OAI22_X1 port map( A1 => n7595, A2 => n5791, B1 => n5829, B2 => n5790
                           , ZN => n1426);
   U918 : OAI22_X1 port map( A1 => n7596, A2 => n5791, B1 => n5830, B2 => n5789
                           , ZN => n1425);
   U919 : OAI22_X1 port map( A1 => n7597, A2 => n5791, B1 => n5831, B2 => n5790
                           , ZN => n1424);
   U920 : OAI22_X1 port map( A1 => n7854, A2 => n5791, B1 => n5832, B2 => n5789
                           , ZN => n1423);
   U921 : OAI22_X1 port map( A1 => n7855, A2 => n5791, B1 => n5833, B2 => n5790
                           , ZN => n1422);
   U922 : OAI22_X1 port map( A1 => n8396, A2 => n5791, B1 => n5834, B2 => n5789
                           , ZN => n1421);
   U923 : OAI22_X1 port map( A1 => n7856, A2 => n5791, B1 => n5835, B2 => n5789
                           , ZN => n1420);
   U924 : OAI22_X1 port map( A1 => n7598, A2 => n5791, B1 => n5836, B2 => n5790
                           , ZN => n1419);
   U925 : OAI22_X1 port map( A1 => n7599, A2 => n5791, B1 => n5837, B2 => n5789
                           , ZN => n1418);
   U926 : OAI22_X1 port map( A1 => n7600, A2 => n5791, B1 => n5838, B2 => n5790
                           , ZN => n1417);
   U927 : OAI22_X1 port map( A1 => n7857, A2 => n5791, B1 => n5839, B2 => n5789
                           , ZN => n1416);
   U928 : OAI22_X1 port map( A1 => n7858, A2 => n5791, B1 => n5840, B2 => n5790
                           , ZN => n1415);
   U929 : OAI22_X1 port map( A1 => n7859, A2 => n5791, B1 => n5841, B2 => n5789
                           , ZN => n1414);
   U930 : OAI22_X1 port map( A1 => n7860, A2 => n5791, B1 => n5842, B2 => n5789
                           , ZN => n1413);
   U931 : OAI22_X1 port map( A1 => n7861, A2 => n5791, B1 => n5843, B2 => n5789
                           , ZN => n1412);
   U932 : OAI22_X1 port map( A1 => n7601, A2 => n5791, B1 => n5844, B2 => n5789
                           , ZN => n1411);
   U933 : OAI22_X1 port map( A1 => n7862, A2 => n5791, B1 => n5845, B2 => n5789
                           , ZN => n1410);
   U934 : OAI22_X1 port map( A1 => n8143, A2 => n5791, B1 => n5846, B2 => n5789
                           , ZN => n1409);
   U935 : OAI22_X1 port map( A1 => n8144, A2 => n5791, B1 => n5848, B2 => n5789
                           , ZN => n1408);
   U936 : OAI22_X1 port map( A1 => n7602, A2 => n5791, B1 => n5849, B2 => n5790
                           , ZN => n1407);
   U937 : OAI22_X1 port map( A1 => n7603, A2 => n5791, B1 => n5850, B2 => n5790
                           , ZN => n1406);
   U938 : OAI22_X1 port map( A1 => n7863, A2 => n5791, B1 => n5851, B2 => n5790
                           , ZN => n1405);
   U939 : OAI22_X1 port map( A1 => n7864, A2 => n5791, B1 => n5852, B2 => n5790
                           , ZN => n1404);
   U940 : OAI22_X1 port map( A1 => n7604, A2 => n5791, B1 => n5853, B2 => n5790
                           , ZN => n1403);
   U941 : OAI22_X1 port map( A1 => n7605, A2 => n5791, B1 => n5854, B2 => n5790
                           , ZN => n1402);
   U942 : OAI22_X1 port map( A1 => n7606, A2 => n5791, B1 => n5855, B2 => n5790
                           , ZN => n1401);
   U943 : OAI22_X1 port map( A1 => n7865, A2 => n5791, B1 => n5856, B2 => n5790
                           , ZN => n1400);
   U944 : OAI22_X1 port map( A1 => n7607, A2 => n5791, B1 => n5858, B2 => n5790
                           , ZN => n1399);
   U945 : NAND2_X1 port map( A1 => n5794, A2 => n5823, ZN => n5795);
   U946 : CLKBUF_X1 port map( A => n5795, Z => n5796);
   U947 : OAI22_X1 port map( A1 => n7425, A2 => n5797, B1 => n5825, B2 => n5796
                           , ZN => n1398);
   U948 : OAI22_X1 port map( A1 => n8397, A2 => n5797, B1 => n5826, B2 => n5795
                           , ZN => n1397);
   U949 : OAI22_X1 port map( A1 => n8145, A2 => n5797, B1 => n5827, B2 => n5796
                           , ZN => n1396);
   U950 : OAI22_X1 port map( A1 => n8398, A2 => n5797, B1 => n5828, B2 => n5795
                           , ZN => n1395);
   U951 : OAI22_X1 port map( A1 => n8399, A2 => n5797, B1 => n5829, B2 => n5796
                           , ZN => n1394);
   U952 : OAI22_X1 port map( A1 => n8146, A2 => n5797, B1 => n5830, B2 => n5795
                           , ZN => n1393);
   U953 : OAI22_X1 port map( A1 => n8400, A2 => n5797, B1 => n5831, B2 => n5796
                           , ZN => n1392);
   U954 : OAI22_X1 port map( A1 => n7608, A2 => n5797, B1 => n5832, B2 => n5795
                           , ZN => n1391);
   U955 : OAI22_X1 port map( A1 => n8147, A2 => n5797, B1 => n5833, B2 => n5796
                           , ZN => n1390);
   U956 : OAI22_X1 port map( A1 => n8401, A2 => n5797, B1 => n5834, B2 => n5795
                           , ZN => n1389);
   U957 : OAI22_X1 port map( A1 => n8402, A2 => n5797, B1 => n5835, B2 => n5795
                           , ZN => n1388);
   U958 : OAI22_X1 port map( A1 => n8403, A2 => n5797, B1 => n5836, B2 => n5796
                           , ZN => n1387);
   U959 : OAI22_X1 port map( A1 => n8404, A2 => n5797, B1 => n5837, B2 => n5795
                           , ZN => n1386);
   U960 : OAI22_X1 port map( A1 => n8405, A2 => n5797, B1 => n5838, B2 => n5796
                           , ZN => n1385);
   U961 : OAI22_X1 port map( A1 => n7866, A2 => n5797, B1 => n5839, B2 => n5795
                           , ZN => n1384);
   U962 : OAI22_X1 port map( A1 => n7867, A2 => n5797, B1 => n5840, B2 => n5796
                           , ZN => n1383);
   U963 : OAI22_X1 port map( A1 => n8406, A2 => n5797, B1 => n5841, B2 => n5795
                           , ZN => n1382);
   U964 : OAI22_X1 port map( A1 => n8407, A2 => n5797, B1 => n5842, B2 => n5795
                           , ZN => n1381);
   U965 : OAI22_X1 port map( A1 => n8148, A2 => n5797, B1 => n5843, B2 => n5795
                           , ZN => n1380);
   U966 : OAI22_X1 port map( A1 => n8408, A2 => n5797, B1 => n5844, B2 => n5795
                           , ZN => n1379);
   U967 : OAI22_X1 port map( A1 => n8149, A2 => n5797, B1 => n5845, B2 => n5795
                           , ZN => n1378);
   U968 : OAI22_X1 port map( A1 => n8409, A2 => n5797, B1 => n5846, B2 => n5795
                           , ZN => n1377);
   U969 : OAI22_X1 port map( A1 => n7609, A2 => n5797, B1 => n5848, B2 => n5795
                           , ZN => n1376);
   U970 : OAI22_X1 port map( A1 => n8410, A2 => n5797, B1 => n5849, B2 => n5796
                           , ZN => n1375);
   U971 : OAI22_X1 port map( A1 => n8411, A2 => n5797, B1 => n5850, B2 => n5796
                           , ZN => n1374);
   U972 : OAI22_X1 port map( A1 => n8150, A2 => n5797, B1 => n5851, B2 => n5796
                           , ZN => n1373);
   U973 : OAI22_X1 port map( A1 => n8151, A2 => n5797, B1 => n5852, B2 => n5796
                           , ZN => n1372);
   U974 : OAI22_X1 port map( A1 => n7868, A2 => n5797, B1 => n5853, B2 => n5796
                           , ZN => n1371);
   U975 : OAI22_X1 port map( A1 => n7610, A2 => n5797, B1 => n5854, B2 => n5796
                           , ZN => n1370);
   U976 : OAI22_X1 port map( A1 => n8412, A2 => n5797, B1 => n5855, B2 => n5796
                           , ZN => n1369);
   U977 : OAI22_X1 port map( A1 => n7869, A2 => n5797, B1 => n5856, B2 => n5796
                           , ZN => n1368);
   U978 : OAI22_X1 port map( A1 => n7870, A2 => n5797, B1 => n5858, B2 => n5796
                           , ZN => n1367);
   U979 : NAND2_X1 port map( A1 => n5798, A2 => n5823, ZN => n5799);
   U980 : CLKBUF_X1 port map( A => n5799, Z => n5800);
   U981 : OAI22_X1 port map( A1 => n7688, A2 => n5801, B1 => n5825, B2 => n5800
                           , ZN => n1366);
   U982 : OAI22_X1 port map( A1 => n7611, A2 => n5801, B1 => n5826, B2 => n5799
                           , ZN => n1365);
   U983 : OAI22_X1 port map( A1 => n8152, A2 => n5801, B1 => n5827, B2 => n5800
                           , ZN => n1364);
   U984 : OAI22_X1 port map( A1 => n7871, A2 => n5801, B1 => n5828, B2 => n5799
                           , ZN => n1363);
   U985 : OAI22_X1 port map( A1 => n7612, A2 => n5801, B1 => n5829, B2 => n5800
                           , ZN => n1362);
   U986 : OAI22_X1 port map( A1 => n7872, A2 => n5801, B1 => n5830, B2 => n5799
                           , ZN => n1361);
   U987 : OAI22_X1 port map( A1 => n7873, A2 => n5801, B1 => n5831, B2 => n5800
                           , ZN => n1360);
   U988 : OAI22_X1 port map( A1 => n7613, A2 => n5801, B1 => n5832, B2 => n5799
                           , ZN => n1359);
   U989 : OAI22_X1 port map( A1 => n7874, A2 => n5801, B1 => n5833, B2 => n5800
                           , ZN => n1358);
   U990 : OAI22_X1 port map( A1 => n7875, A2 => n5801, B1 => n5834, B2 => n5799
                           , ZN => n1357);
   U991 : OAI22_X1 port map( A1 => n7876, A2 => n5801, B1 => n5835, B2 => n5799
                           , ZN => n1356);
   U992 : OAI22_X1 port map( A1 => n7877, A2 => n5801, B1 => n5836, B2 => n5800
                           , ZN => n1355);
   U993 : OAI22_X1 port map( A1 => n7614, A2 => n5801, B1 => n5837, B2 => n5799
                           , ZN => n1354);
   U994 : OAI22_X1 port map( A1 => n7878, A2 => n5801, B1 => n5838, B2 => n5800
                           , ZN => n1353);
   U995 : OAI22_X1 port map( A1 => n8413, A2 => n5801, B1 => n5839, B2 => n5799
                           , ZN => n1352);
   U996 : OAI22_X1 port map( A1 => n7615, A2 => n5801, B1 => n5840, B2 => n5800
                           , ZN => n1351);
   U997 : OAI22_X1 port map( A1 => n7616, A2 => n5801, B1 => n5841, B2 => n5799
                           , ZN => n1350);
   U998 : OAI22_X1 port map( A1 => n7617, A2 => n5801, B1 => n5842, B2 => n5799
                           , ZN => n1349);
   U999 : OAI22_X1 port map( A1 => n7879, A2 => n5801, B1 => n5843, B2 => n5799
                           , ZN => n1348);
   U1000 : OAI22_X1 port map( A1 => n7880, A2 => n5801, B1 => n5844, B2 => 
                           n5799, ZN => n1347);
   U1001 : OAI22_X1 port map( A1 => n7618, A2 => n5801, B1 => n5845, B2 => 
                           n5799, ZN => n1346);
   U1002 : OAI22_X1 port map( A1 => n7881, A2 => n5801, B1 => n5846, B2 => 
                           n5799, ZN => n1345);
   U1003 : OAI22_X1 port map( A1 => n7882, A2 => n5801, B1 => n5848, B2 => 
                           n5799, ZN => n1344);
   U1004 : OAI22_X1 port map( A1 => n7619, A2 => n5801, B1 => n5849, B2 => 
                           n5800, ZN => n1343);
   U1005 : OAI22_X1 port map( A1 => n7620, A2 => n5801, B1 => n5850, B2 => 
                           n5800, ZN => n1342);
   U1006 : OAI22_X1 port map( A1 => n8414, A2 => n5801, B1 => n5851, B2 => 
                           n5800, ZN => n1341);
   U1007 : OAI22_X1 port map( A1 => n8415, A2 => n5801, B1 => n5852, B2 => 
                           n5800, ZN => n1340);
   U1008 : OAI22_X1 port map( A1 => n7621, A2 => n5801, B1 => n5853, B2 => 
                           n5800, ZN => n1339);
   U1009 : OAI22_X1 port map( A1 => n7622, A2 => n5801, B1 => n5854, B2 => 
                           n5800, ZN => n1338);
   U1010 : OAI22_X1 port map( A1 => n7623, A2 => n5801, B1 => n5855, B2 => 
                           n5800, ZN => n1337);
   U1011 : OAI22_X1 port map( A1 => n7624, A2 => n5801, B1 => n5856, B2 => 
                           n5800, ZN => n1336);
   U1012 : OAI22_X1 port map( A1 => n7625, A2 => n5801, B1 => n5858, B2 => 
                           n5800, ZN => n1335);
   U1013 : NAND2_X1 port map( A1 => n5802, A2 => n5823, ZN => n5803);
   U1014 : CLKBUF_X1 port map( A => n5806, Z => n5804);
   U1015 : CLKBUF_X1 port map( A => n5803, Z => n5805);
   U1016 : OAI22_X1 port map( A1 => n7689, A2 => n5804, B1 => n5825, B2 => 
                           n5805, ZN => n1334);
   U1017 : OAI22_X1 port map( A1 => n8416, A2 => n5806, B1 => n5826, B2 => 
                           n5803, ZN => n1333);
   U1018 : OAI22_X1 port map( A1 => n8153, A2 => n5804, B1 => n5827, B2 => 
                           n5805, ZN => n1332);
   U1019 : OAI22_X1 port map( A1 => n8154, A2 => n5806, B1 => n5828, B2 => 
                           n5803, ZN => n1331);
   U1020 : OAI22_X1 port map( A1 => n8417, A2 => n5804, B1 => n5829, B2 => 
                           n5805, ZN => n1330);
   U1021 : OAI22_X1 port map( A1 => n8418, A2 => n5806, B1 => n5830, B2 => 
                           n5803, ZN => n1329);
   U1022 : OAI22_X1 port map( A1 => n8155, A2 => n5804, B1 => n5831, B2 => 
                           n5805, ZN => n1328);
   U1023 : OAI22_X1 port map( A1 => n7883, A2 => n5806, B1 => n5832, B2 => 
                           n5803, ZN => n1327);
   U1024 : OAI22_X1 port map( A1 => n7884, A2 => n5804, B1 => n5833, B2 => 
                           n5805, ZN => n1326);
   U1025 : OAI22_X1 port map( A1 => n8419, A2 => n5806, B1 => n5834, B2 => 
                           n5803, ZN => n1325);
   U1026 : OAI22_X1 port map( A1 => n7885, A2 => n5806, B1 => n5835, B2 => 
                           n5803, ZN => n1324);
   U1027 : OAI22_X1 port map( A1 => n7886, A2 => n5806, B1 => n5836, B2 => 
                           n5805, ZN => n1323);
   U1028 : OAI22_X1 port map( A1 => n8156, A2 => n5804, B1 => n5837, B2 => 
                           n5803, ZN => n1322);
   U1029 : OAI22_X1 port map( A1 => n8157, A2 => n5804, B1 => n5838, B2 => 
                           n5805, ZN => n1321);
   U1030 : OAI22_X1 port map( A1 => n7626, A2 => n5804, B1 => n5839, B2 => 
                           n5803, ZN => n1320);
   U1031 : OAI22_X1 port map( A1 => n7887, A2 => n5804, B1 => n5840, B2 => 
                           n5805, ZN => n1319);
   U1032 : OAI22_X1 port map( A1 => n8420, A2 => n5804, B1 => n5841, B2 => 
                           n5803, ZN => n1318);
   U1033 : OAI22_X1 port map( A1 => n7627, A2 => n5804, B1 => n5842, B2 => 
                           n5803, ZN => n1317);
   U1034 : OAI22_X1 port map( A1 => n8421, A2 => n5804, B1 => n5843, B2 => 
                           n5803, ZN => n1316);
   U1035 : OAI22_X1 port map( A1 => n8422, A2 => n5804, B1 => n5844, B2 => 
                           n5803, ZN => n1315);
   U1036 : OAI22_X1 port map( A1 => n7628, A2 => n5804, B1 => n5845, B2 => 
                           n5803, ZN => n1314);
   U1037 : OAI22_X1 port map( A1 => n8423, A2 => n5804, B1 => n5846, B2 => 
                           n5803, ZN => n1313);
   U1038 : OAI22_X1 port map( A1 => n7888, A2 => n5804, B1 => n5848, B2 => 
                           n5803, ZN => n1312);
   U1039 : OAI22_X1 port map( A1 => n7629, A2 => n5804, B1 => n5849, B2 => 
                           n5805, ZN => n1311);
   U1040 : OAI22_X1 port map( A1 => n8158, A2 => n5806, B1 => n5850, B2 => 
                           n5805, ZN => n1310);
   U1041 : OAI22_X1 port map( A1 => n8159, A2 => n5806, B1 => n5851, B2 => 
                           n5805, ZN => n1309);
   U1042 : OAI22_X1 port map( A1 => n8424, A2 => n5806, B1 => n5852, B2 => 
                           n5805, ZN => n1308);
   U1043 : OAI22_X1 port map( A1 => n8160, A2 => n5806, B1 => n5853, B2 => 
                           n5805, ZN => n1307);
   U1044 : OAI22_X1 port map( A1 => n7889, A2 => n5806, B1 => n5854, B2 => 
                           n5805, ZN => n1306);
   U1045 : OAI22_X1 port map( A1 => n8425, A2 => n5806, B1 => n5855, B2 => 
                           n5805, ZN => n1305);
   U1046 : OAI22_X1 port map( A1 => n8426, A2 => n5806, B1 => n5856, B2 => 
                           n5805, ZN => n1304);
   U1047 : OAI22_X1 port map( A1 => n8161, A2 => n5806, B1 => n5858, B2 => 
                           n5805, ZN => n1303);
   U1048 : NAND2_X1 port map( A1 => n5807, A2 => n5823, ZN => n5808);
   U1049 : CLKBUF_X1 port map( A => n5808, Z => n5809);
   U1050 : OAI22_X1 port map( A1 => n7426, A2 => n5810, B1 => n5825, B2 => 
                           n5809, ZN => n1302);
   U1051 : OAI22_X1 port map( A1 => n7630, A2 => n5810, B1 => n5826, B2 => 
                           n5808, ZN => n1301);
   U1052 : OAI22_X1 port map( A1 => n7631, A2 => n5810, B1 => n5827, B2 => 
                           n5809, ZN => n1300);
   U1053 : OAI22_X1 port map( A1 => n7890, A2 => n5810, B1 => n5828, B2 => 
                           n5808, ZN => n1299);
   U1054 : OAI22_X1 port map( A1 => n8162, A2 => n5810, B1 => n5829, B2 => 
                           n5809, ZN => n1298);
   U1055 : OAI22_X1 port map( A1 => n7632, A2 => n5810, B1 => n5830, B2 => 
                           n5808, ZN => n1297);
   U1056 : OAI22_X1 port map( A1 => n8163, A2 => n5810, B1 => n5831, B2 => 
                           n5809, ZN => n1296);
   U1057 : OAI22_X1 port map( A1 => n7891, A2 => n5810, B1 => n5832, B2 => 
                           n5808, ZN => n1295);
   U1058 : OAI22_X1 port map( A1 => n8164, A2 => n5810, B1 => n5833, B2 => 
                           n5809, ZN => n1294);
   U1059 : OAI22_X1 port map( A1 => n7633, A2 => n5810, B1 => n5834, B2 => 
                           n5808, ZN => n1293);
   U1060 : OAI22_X1 port map( A1 => n8165, A2 => n5810, B1 => n5835, B2 => 
                           n5808, ZN => n1292);
   U1061 : OAI22_X1 port map( A1 => n7634, A2 => n5810, B1 => n5836, B2 => 
                           n5809, ZN => n1291);
   U1062 : OAI22_X1 port map( A1 => n7892, A2 => n5810, B1 => n5837, B2 => 
                           n5808, ZN => n1290);
   U1063 : OAI22_X1 port map( A1 => n7635, A2 => n5810, B1 => n5838, B2 => 
                           n5809, ZN => n1289);
   U1064 : OAI22_X1 port map( A1 => n7636, A2 => n5810, B1 => n5839, B2 => 
                           n5808, ZN => n1288);
   U1065 : OAI22_X1 port map( A1 => n7637, A2 => n5810, B1 => n5840, B2 => 
                           n5809, ZN => n1287);
   U1066 : OAI22_X1 port map( A1 => n7893, A2 => n5810, B1 => n5841, B2 => 
                           n5808, ZN => n1286);
   U1067 : OAI22_X1 port map( A1 => n7638, A2 => n5810, B1 => n5842, B2 => 
                           n5808, ZN => n1285);
   U1068 : OAI22_X1 port map( A1 => n7639, A2 => n5810, B1 => n5843, B2 => 
                           n5808, ZN => n1284);
   U1069 : OAI22_X1 port map( A1 => n7640, A2 => n5810, B1 => n5844, B2 => 
                           n5808, ZN => n1283);
   U1070 : OAI22_X1 port map( A1 => n8427, A2 => n5810, B1 => n5845, B2 => 
                           n5808, ZN => n1282);
   U1071 : OAI22_X1 port map( A1 => n7641, A2 => n5810, B1 => n5846, B2 => 
                           n5808, ZN => n1281);
   U1072 : OAI22_X1 port map( A1 => n7894, A2 => n5810, B1 => n5848, B2 => 
                           n5808, ZN => n1280);
   U1073 : OAI22_X1 port map( A1 => n7895, A2 => n5810, B1 => n5849, B2 => 
                           n5809, ZN => n1279);
   U1074 : OAI22_X1 port map( A1 => n7642, A2 => n5810, B1 => n5850, B2 => 
                           n5809, ZN => n1278);
   U1075 : OAI22_X1 port map( A1 => n7643, A2 => n5810, B1 => n5851, B2 => 
                           n5809, ZN => n1277);
   U1076 : OAI22_X1 port map( A1 => n7896, A2 => n5810, B1 => n5852, B2 => 
                           n5809, ZN => n1276);
   U1077 : OAI22_X1 port map( A1 => n7897, A2 => n5810, B1 => n5853, B2 => 
                           n5809, ZN => n1275);
   U1078 : OAI22_X1 port map( A1 => n8428, A2 => n5810, B1 => n5854, B2 => 
                           n5809, ZN => n1274);
   U1079 : OAI22_X1 port map( A1 => n7898, A2 => n5810, B1 => n5855, B2 => 
                           n5809, ZN => n1273);
   U1080 : OAI22_X1 port map( A1 => n7644, A2 => n5810, B1 => n5856, B2 => 
                           n5809, ZN => n1272);
   U1081 : OAI22_X1 port map( A1 => n8429, A2 => n5810, B1 => n5858, B2 => 
                           n5809, ZN => n1271);
   U1082 : NAND2_X1 port map( A1 => n5811, A2 => n5823, ZN => n5812);
   U1083 : CLKBUF_X1 port map( A => n5812, Z => n5813);
   U1084 : OAI22_X1 port map( A1 => n7690, A2 => n5814, B1 => n5825, B2 => 
                           n5813, ZN => n1270);
   U1085 : OAI22_X1 port map( A1 => n7645, A2 => n5814, B1 => n5826, B2 => 
                           n5812, ZN => n1269);
   U1086 : OAI22_X1 port map( A1 => n7899, A2 => n5814, B1 => n5827, B2 => 
                           n5813, ZN => n1268);
   U1087 : OAI22_X1 port map( A1 => n8166, A2 => n5814, B1 => n5828, B2 => 
                           n5812, ZN => n1267);
   U1088 : OAI22_X1 port map( A1 => n7646, A2 => n5814, B1 => n5829, B2 => 
                           n5813, ZN => n1266);
   U1089 : OAI22_X1 port map( A1 => n8430, A2 => n5814, B1 => n5830, B2 => 
                           n5812, ZN => n1265);
   U1090 : OAI22_X1 port map( A1 => n7647, A2 => n5814, B1 => n5831, B2 => 
                           n5813, ZN => n1264);
   U1091 : OAI22_X1 port map( A1 => n8167, A2 => n5814, B1 => n5832, B2 => 
                           n5812, ZN => n1263);
   U1092 : OAI22_X1 port map( A1 => n7900, A2 => n5814, B1 => n5833, B2 => 
                           n5813, ZN => n1262);
   U1093 : OAI22_X1 port map( A1 => n7901, A2 => n5814, B1 => n5834, B2 => 
                           n5812, ZN => n1261);
   U1094 : OAI22_X1 port map( A1 => n7902, A2 => n5814, B1 => n5835, B2 => 
                           n5812, ZN => n1260);
   U1095 : OAI22_X1 port map( A1 => n8431, A2 => n5814, B1 => n5836, B2 => 
                           n5813, ZN => n1259);
   U1096 : OAI22_X1 port map( A1 => n8432, A2 => n5814, B1 => n5837, B2 => 
                           n5812, ZN => n1258);
   U1097 : OAI22_X1 port map( A1 => n8433, A2 => n5814, B1 => n5838, B2 => 
                           n5813, ZN => n1257);
   U1098 : OAI22_X1 port map( A1 => n8168, A2 => n5814, B1 => n5839, B2 => 
                           n5812, ZN => n1256);
   U1099 : OAI22_X1 port map( A1 => n8169, A2 => n5814, B1 => n5840, B2 => 
                           n5813, ZN => n1255);
   U1100 : OAI22_X1 port map( A1 => n7648, A2 => n5814, B1 => n5841, B2 => 
                           n5812, ZN => n1254);
   U1101 : OAI22_X1 port map( A1 => n7649, A2 => n5814, B1 => n5842, B2 => 
                           n5812, ZN => n1253);
   U1102 : OAI22_X1 port map( A1 => n7650, A2 => n5814, B1 => n5843, B2 => 
                           n5812, ZN => n1252);
   U1103 : OAI22_X1 port map( A1 => n7651, A2 => n5814, B1 => n5844, B2 => 
                           n5812, ZN => n1251);
   U1104 : OAI22_X1 port map( A1 => n7652, A2 => n5814, B1 => n5845, B2 => 
                           n5812, ZN => n1250);
   U1105 : OAI22_X1 port map( A1 => n7903, A2 => n5814, B1 => n5846, B2 => 
                           n5812, ZN => n1249);
   U1106 : OAI22_X1 port map( A1 => n8170, A2 => n5814, B1 => n5848, B2 => 
                           n5812, ZN => n1248);
   U1107 : OAI22_X1 port map( A1 => n8434, A2 => n5814, B1 => n5849, B2 => 
                           n5813, ZN => n1247);
   U1108 : OAI22_X1 port map( A1 => n8171, A2 => n5814, B1 => n5850, B2 => 
                           n5813, ZN => n1246);
   U1109 : OAI22_X1 port map( A1 => n7904, A2 => n5814, B1 => n5851, B2 => 
                           n5813, ZN => n1245);
   U1110 : OAI22_X1 port map( A1 => n7905, A2 => n5814, B1 => n5852, B2 => 
                           n5813, ZN => n1244);
   U1111 : OAI22_X1 port map( A1 => n8435, A2 => n5814, B1 => n5853, B2 => 
                           n5813, ZN => n1243);
   U1112 : OAI22_X1 port map( A1 => n8436, A2 => n5814, B1 => n5854, B2 => 
                           n5813, ZN => n1242);
   U1113 : OAI22_X1 port map( A1 => n8172, A2 => n5814, B1 => n5855, B2 => 
                           n5813, ZN => n1241);
   U1114 : OAI22_X1 port map( A1 => n7906, A2 => n5814, B1 => n5856, B2 => 
                           n5813, ZN => n1240);
   U1115 : OAI22_X1 port map( A1 => n8173, A2 => n5814, B1 => n5858, B2 => 
                           n5813, ZN => n1239);
   U1116 : NAND2_X1 port map( A1 => n5815, A2 => n5823, ZN => n5816);
   U1117 : CLKBUF_X1 port map( A => n5816, Z => n5817);
   U1118 : OAI22_X1 port map( A1 => n7691, A2 => n5818, B1 => n5825, B2 => 
                           n5817, ZN => n1238);
   U1119 : OAI22_X1 port map( A1 => n7907, A2 => n5818, B1 => n5826, B2 => 
                           n5816, ZN => n1237);
   U1120 : OAI22_X1 port map( A1 => n7653, A2 => n5818, B1 => n5827, B2 => 
                           n5817, ZN => n1236);
   U1121 : OAI22_X1 port map( A1 => n7654, A2 => n5818, B1 => n5828, B2 => 
                           n5816, ZN => n1235);
   U1122 : OAI22_X1 port map( A1 => n7908, A2 => n5818, B1 => n5829, B2 => 
                           n5817, ZN => n1234);
   U1123 : OAI22_X1 port map( A1 => n7909, A2 => n5818, B1 => n5830, B2 => 
                           n5816, ZN => n1233);
   U1124 : OAI22_X1 port map( A1 => n7655, A2 => n5818, B1 => n5831, B2 => 
                           n5817, ZN => n1232);
   U1125 : OAI22_X1 port map( A1 => n7910, A2 => n5818, B1 => n5832, B2 => 
                           n5816, ZN => n1231);
   U1126 : OAI22_X1 port map( A1 => n7656, A2 => n5818, B1 => n5833, B2 => 
                           n5817, ZN => n1230);
   U1127 : OAI22_X1 port map( A1 => n7657, A2 => n5818, B1 => n5834, B2 => 
                           n5816, ZN => n1229);
   U1128 : OAI22_X1 port map( A1 => n7658, A2 => n5818, B1 => n5835, B2 => 
                           n5816, ZN => n1228);
   U1129 : OAI22_X1 port map( A1 => n8174, A2 => n5818, B1 => n5836, B2 => 
                           n5817, ZN => n1227);
   U1130 : OAI22_X1 port map( A1 => n7911, A2 => n5818, B1 => n5837, B2 => 
                           n5816, ZN => n1226);
   U1131 : OAI22_X1 port map( A1 => n7912, A2 => n5818, B1 => n5838, B2 => 
                           n5817, ZN => n1225);
   U1132 : OAI22_X1 port map( A1 => n7913, A2 => n5818, B1 => n5839, B2 => 
                           n5816, ZN => n1224);
   U1133 : OAI22_X1 port map( A1 => n8437, A2 => n5818, B1 => n5840, B2 => 
                           n5817, ZN => n1223);
   U1134 : OAI22_X1 port map( A1 => n8438, A2 => n5818, B1 => n5841, B2 => 
                           n5816, ZN => n1222);
   U1135 : OAI22_X1 port map( A1 => n7659, A2 => n5818, B1 => n5842, B2 => 
                           n5816, ZN => n1221);
   U1136 : OAI22_X1 port map( A1 => n7914, A2 => n5818, B1 => n5843, B2 => 
                           n5816, ZN => n1220);
   U1137 : OAI22_X1 port map( A1 => n7915, A2 => n5818, B1 => n5844, B2 => 
                           n5816, ZN => n1219);
   U1138 : OAI22_X1 port map( A1 => n8439, A2 => n5818, B1 => n5845, B2 => 
                           n5816, ZN => n1218);
   U1139 : OAI22_X1 port map( A1 => n7660, A2 => n5818, B1 => n5846, B2 => 
                           n5816, ZN => n1217);
   U1140 : OAI22_X1 port map( A1 => n7661, A2 => n5818, B1 => n5848, B2 => 
                           n5816, ZN => n1216);
   U1141 : OAI22_X1 port map( A1 => n7916, A2 => n5818, B1 => n5849, B2 => 
                           n5817, ZN => n1215);
   U1142 : OAI22_X1 port map( A1 => n7917, A2 => n5818, B1 => n5850, B2 => 
                           n5817, ZN => n1214);
   U1143 : OAI22_X1 port map( A1 => n7662, A2 => n5818, B1 => n5851, B2 => 
                           n5817, ZN => n1213);
   U1144 : OAI22_X1 port map( A1 => n8175, A2 => n5818, B1 => n5852, B2 => 
                           n5817, ZN => n1212);
   U1145 : OAI22_X1 port map( A1 => n7663, A2 => n5818, B1 => n5853, B2 => 
                           n5817, ZN => n1211);
   U1146 : OAI22_X1 port map( A1 => n7918, A2 => n5818, B1 => n5854, B2 => 
                           n5817, ZN => n1210);
   U1147 : OAI22_X1 port map( A1 => n7919, A2 => n5818, B1 => n5855, B2 => 
                           n5817, ZN => n1209);
   U1148 : OAI22_X1 port map( A1 => n7664, A2 => n5818, B1 => n5856, B2 => 
                           n5817, ZN => n1208);
   U1149 : OAI22_X1 port map( A1 => n7665, A2 => n5818, B1 => n5858, B2 => 
                           n5817, ZN => n1207);
   U1150 : NAND2_X1 port map( A1 => n5819, A2 => n5823, ZN => n5820);
   U1151 : OAI22_X1 port map( A1 => n7427, A2 => n5822, B1 => n5825, B2 => 
                           n5821, ZN => n1206);
   U1152 : OAI22_X1 port map( A1 => n7666, A2 => n5822, B1 => n5826, B2 => 
                           n5820, ZN => n1205);
   U1153 : OAI22_X1 port map( A1 => n7667, A2 => n5822, B1 => n5827, B2 => 
                           n5821, ZN => n1204);
   U1154 : OAI22_X1 port map( A1 => n7920, A2 => n5822, B1 => n5828, B2 => 
                           n5820, ZN => n1203);
   U1155 : OAI22_X1 port map( A1 => n7921, A2 => n5822, B1 => n5829, B2 => 
                           n5821, ZN => n1202);
   U1156 : OAI22_X1 port map( A1 => n7668, A2 => n5822, B1 => n5830, B2 => 
                           n5820, ZN => n1201);
   U1157 : OAI22_X1 port map( A1 => n7669, A2 => n5822, B1 => n5831, B2 => 
                           n5821, ZN => n1200);
   U1158 : OAI22_X1 port map( A1 => n7922, A2 => n5822, B1 => n5832, B2 => 
                           n5820, ZN => n1199);
   U1159 : OAI22_X1 port map( A1 => n7923, A2 => n5822, B1 => n5833, B2 => 
                           n5821, ZN => n1198);
   U1160 : OAI22_X1 port map( A1 => n7924, A2 => n5822, B1 => n5834, B2 => 
                           n5820, ZN => n1197);
   U1161 : OAI22_X1 port map( A1 => n7670, A2 => n5822, B1 => n5835, B2 => 
                           n5820, ZN => n1196);
   U1162 : OAI22_X1 port map( A1 => n7925, A2 => n5822, B1 => n5836, B2 => 
                           n5821, ZN => n1195);
   U1163 : OAI22_X1 port map( A1 => n7671, A2 => n5822, B1 => n5837, B2 => 
                           n5820, ZN => n1194);
   U1164 : OAI22_X1 port map( A1 => n7672, A2 => n5822, B1 => n5838, B2 => 
                           n5821, ZN => n1193);
   U1165 : OAI22_X1 port map( A1 => n7673, A2 => n5822, B1 => n5839, B2 => 
                           n5820, ZN => n1192);
   U1166 : OAI22_X1 port map( A1 => n7674, A2 => n5822, B1 => n5840, B2 => 
                           n5821, ZN => n1191);
   U1167 : OAI22_X1 port map( A1 => n7926, A2 => n5822, B1 => n5841, B2 => 
                           n5820, ZN => n1190);
   U1168 : OAI22_X1 port map( A1 => n7675, A2 => n5822, B1 => n5842, B2 => 
                           n5820, ZN => n1189);
   U1169 : OAI22_X1 port map( A1 => n7676, A2 => n5822, B1 => n5843, B2 => 
                           n5820, ZN => n1188);
   U1170 : OAI22_X1 port map( A1 => n7927, A2 => n5822, B1 => n5844, B2 => 
                           n5820, ZN => n1187);
   U1171 : OAI22_X1 port map( A1 => n7928, A2 => n5822, B1 => n5845, B2 => 
                           n5820, ZN => n1186);
   U1172 : OAI22_X1 port map( A1 => n7929, A2 => n5822, B1 => n5846, B2 => 
                           n5820, ZN => n1185);
   U1173 : OAI22_X1 port map( A1 => n7930, A2 => n5822, B1 => n5848, B2 => 
                           n5820, ZN => n1184);
   U1174 : OAI22_X1 port map( A1 => n7677, A2 => n5822, B1 => n5849, B2 => 
                           n5821, ZN => n1183);
   U1175 : OAI22_X1 port map( A1 => n7931, A2 => n5822, B1 => n5850, B2 => 
                           n5821, ZN => n1182);
   U1176 : OAI22_X1 port map( A1 => n7678, A2 => n5822, B1 => n5851, B2 => 
                           n5821, ZN => n1181);
   U1177 : OAI22_X1 port map( A1 => n7679, A2 => n5822, B1 => n5852, B2 => 
                           n5821, ZN => n1180);
   U1178 : OAI22_X1 port map( A1 => n7932, A2 => n5822, B1 => n5853, B2 => 
                           n5821, ZN => n1179);
   U1179 : OAI22_X1 port map( A1 => n7680, A2 => n5822, B1 => n5854, B2 => 
                           n5821, ZN => n1178);
   U1180 : OAI22_X1 port map( A1 => n7681, A2 => n5822, B1 => n5855, B2 => 
                           n5821, ZN => n1177);
   U1181 : OAI22_X1 port map( A1 => n7933, A2 => n5822, B1 => n5856, B2 => 
                           n5821, ZN => n1176);
   U1182 : OAI22_X1 port map( A1 => n7934, A2 => n5822, B1 => n5858, B2 => 
                           n5821, ZN => n1175);
   U1183 : NAND2_X1 port map( A1 => n5824, A2 => n5823, ZN => n5847);
   U1184 : CLKBUF_X1 port map( A => n5847, Z => n5857);
   U1185 : OAI22_X1 port map( A1 => n7943, A2 => n5859, B1 => n5825, B2 => 
                           n5857, ZN => n1174);
   U1186 : OAI22_X1 port map( A1 => n8440, A2 => n5859, B1 => n5826, B2 => 
                           n5847, ZN => n1173);
   U1187 : OAI22_X1 port map( A1 => n7935, A2 => n5859, B1 => n5827, B2 => 
                           n5857, ZN => n1172);
   U1188 : OAI22_X1 port map( A1 => n8176, A2 => n5859, B1 => n5828, B2 => 
                           n5847, ZN => n1171);
   U1189 : OAI22_X1 port map( A1 => n7936, A2 => n5859, B1 => n5829, B2 => 
                           n5857, ZN => n1170);
   U1190 : OAI22_X1 port map( A1 => n8441, A2 => n5859, B1 => n5830, B2 => 
                           n5847, ZN => n1169);
   U1191 : OAI22_X1 port map( A1 => n7937, A2 => n5859, B1 => n5831, B2 => 
                           n5857, ZN => n1168);
   U1192 : OAI22_X1 port map( A1 => n8177, A2 => n5859, B1 => n5832, B2 => 
                           n5847, ZN => n1167);
   U1193 : OAI22_X1 port map( A1 => n8442, A2 => n5859, B1 => n5833, B2 => 
                           n5857, ZN => n1166);
   U1194 : OAI22_X1 port map( A1 => n8178, A2 => n5859, B1 => n5834, B2 => 
                           n5847, ZN => n1165);
   U1195 : OAI22_X1 port map( A1 => n8179, A2 => n5859, B1 => n5835, B2 => 
                           n5847, ZN => n1164);
   U1196 : OAI22_X1 port map( A1 => n8180, A2 => n5859, B1 => n5836, B2 => 
                           n5857, ZN => n1163);
   U1197 : OAI22_X1 port map( A1 => n8181, A2 => n5859, B1 => n5837, B2 => 
                           n5847, ZN => n1162);
   U1198 : OAI22_X1 port map( A1 => n7938, A2 => n5859, B1 => n5838, B2 => 
                           n5857, ZN => n1161);
   U1199 : OAI22_X1 port map( A1 => n8443, A2 => n5859, B1 => n5839, B2 => 
                           n5847, ZN => n1160);
   U1200 : OAI22_X1 port map( A1 => n8182, A2 => n5859, B1 => n5840, B2 => 
                           n5857, ZN => n1159);
   U1201 : OAI22_X1 port map( A1 => n8183, A2 => n5859, B1 => n5841, B2 => 
                           n5847, ZN => n1158);
   U1202 : OAI22_X1 port map( A1 => n8184, A2 => n5859, B1 => n5842, B2 => 
                           n5847, ZN => n1157);
   U1203 : OAI22_X1 port map( A1 => n7682, A2 => n5859, B1 => n5843, B2 => 
                           n5847, ZN => n1156);
   U1204 : OAI22_X1 port map( A1 => n8185, A2 => n5859, B1 => n5844, B2 => 
                           n5847, ZN => n1155);
   U1205 : OAI22_X1 port map( A1 => n8444, A2 => n5859, B1 => n5845, B2 => 
                           n5847, ZN => n1154);
   U1206 : OAI22_X1 port map( A1 => n8186, A2 => n5859, B1 => n5846, B2 => 
                           n5847, ZN => n1153);
   U1207 : OAI22_X1 port map( A1 => n8187, A2 => n5859, B1 => n5848, B2 => 
                           n5847, ZN => n1152);
   U1208 : OAI22_X1 port map( A1 => n7939, A2 => n5859, B1 => n5849, B2 => 
                           n5857, ZN => n1151);
   U1209 : OAI22_X1 port map( A1 => n8445, A2 => n5859, B1 => n5850, B2 => 
                           n5857, ZN => n1150);
   U1210 : OAI22_X1 port map( A1 => n8188, A2 => n5859, B1 => n5851, B2 => 
                           n5857, ZN => n1149);
   U1211 : OAI22_X1 port map( A1 => n7683, A2 => n5859, B1 => n5852, B2 => 
                           n5857, ZN => n1148);
   U1212 : OAI22_X1 port map( A1 => n8189, A2 => n5859, B1 => n5853, B2 => 
                           n5857, ZN => n1147);
   U1213 : OAI22_X1 port map( A1 => n8190, A2 => n5859, B1 => n5854, B2 => 
                           n5857, ZN => n1146);
   U1214 : OAI22_X1 port map( A1 => n8446, A2 => n5859, B1 => n5855, B2 => 
                           n5857, ZN => n1145);
   U1215 : OAI22_X1 port map( A1 => n8191, A2 => n5859, B1 => n5856, B2 => 
                           n5857, ZN => n1144);
   U1216 : OAI22_X1 port map( A1 => n8447, A2 => n5859, B1 => n5858, B2 => 
                           n5857, ZN => n1143);
   U1217 : NAND3_X1 port map( A1 => n5675, A2 => ENABLE, A3 => RD2, ZN => n6641
                           );
   U1218 : INV_X1 port map( A => ADD_RD2(3), ZN => n5888);
   U1219 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n5888, ZN => n5869);
   U1220 : INV_X1 port map( A => ADD_RD2(1), ZN => n5866);
   U1221 : INV_X1 port map( A => ADD_RD2(2), ZN => n5860);
   U1222 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n5866, A3 => n5860, ZN =>
                           n5879);
   U1223 : NOR2_X1 port map( A1 => n5869, A2 => n5879, ZN => n6416);
   U1224 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => n5866, 
                           ZN => n5876);
   U1225 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n5868);
   U1226 : NOR2_X1 port map( A1 => n5876, A2 => n5868, ZN => n6315);
   U1227 : CLKBUF_X1 port map( A => n6315, Z => n6603);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n6416, B1 => 
                           REGISTERS_29_31_port, B2 => n6603, ZN => n5865);
   U1229 : INV_X1 port map( A => ADD_RD2(0), ZN => n5861);
   U1230 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => n5866, A3 => n5861, ZN =>
                           n5880);
   U1231 : NOR2_X1 port map( A1 => n5880, A2 => n5868, ZN => n6561);
   U1232 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => n5860, 
                           ZN => n5881);
   U1233 : NOR2_X1 port map( A1 => n5869, A2 => n5881, ZN => n6604);
   U1234 : CLKBUF_X1 port map( A => n6604, Z => n6562);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n6561, B1 => 
                           REGISTERS_19_31_port, B2 => n6562, ZN => n5864);
   U1236 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n5878);
   U1237 : NOR2_X1 port map( A1 => n5869, A2 => n5878, ZN => n6364);
   U1238 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => n5861, 
                           ZN => n5882);
   U1239 : NOR2_X1 port map( A1 => n5882, A2 => n5868, ZN => n6589);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n6364, B1 => 
                           REGISTERS_30_31_port, B2 => n6589, ZN => n5863);
   U1241 : NOR2_X1 port map( A1 => n5868, A2 => n5879, ZN => n6439);
   U1242 : NOR2_X1 port map( A1 => n5868, A2 => n5881, ZN => n6590);
   U1243 : CLKBUF_X1 port map( A => n6590, Z => n6555);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n6439, B1 => 
                           REGISTERS_27_31_port, B2 => n6555, ZN => n5862);
   U1245 : NAND4_X1 port map( A1 => n5865, A2 => n5864, A3 => n5863, A4 => 
                           n5862, ZN => n5875);
   U1246 : NOR2_X1 port map( A1 => n5869, A2 => n5876, ZN => n6369);
   U1247 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), ZN => n5867);
   U1248 : NAND2_X1 port map( A1 => n5867, A2 => n5866, ZN => n5883);
   U1249 : NOR2_X1 port map( A1 => n5868, A2 => n5883, ZN => n6605);
   U1250 : CLKBUF_X1 port map( A => n6605, Z => n6534);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n6369, B1 => 
                           REGISTERS_24_31_port, B2 => n6534, ZN => n5873);
   U1252 : NOR2_X1 port map( A1 => n5869, A2 => n5882, ZN => n6592);
   U1253 : NOR2_X1 port map( A1 => n5869, A2 => n5880, ZN => n6341);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n6592, B1 => 
                           REGISTERS_20_31_port, B2 => n6341, ZN => n5872);
   U1255 : NOR2_X1 port map( A1 => n5869, A2 => n5883, ZN => n6320);
   U1256 : NAND2_X1 port map( A1 => ADD_RD2(1), A2 => n5867, ZN => n5877);
   U1257 : NOR2_X1 port map( A1 => n5868, A2 => n5877, ZN => n6507);
   U1258 : CLKBUF_X1 port map( A => n6507, Z => n6594);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n6320, B1 => 
                           REGISTERS_26_31_port, B2 => n6594, ZN => n5871);
   U1260 : NOR2_X1 port map( A1 => n5868, A2 => n5878, ZN => n6459);
   U1261 : NOR2_X1 port map( A1 => n5869, A2 => n5877, ZN => n6601);
   U1262 : CLKBUF_X1 port map( A => n6601, Z => n6560);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_31_31_port, A2 => n6459, B1 => 
                           REGISTERS_18_31_port, B2 => n6560, ZN => n5870);
   U1264 : NAND4_X1 port map( A1 => n5873, A2 => n5872, A3 => n5871, A4 => 
                           n5870, ZN => n5874);
   U1265 : NOR2_X1 port map( A1 => n5875, A2 => n5874, ZN => n5896);
   U1266 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n6586, 
                           ZN => n6638);
   U1267 : CLKBUF_X1 port map( A => n6638, Z => n6456);
   U1268 : INV_X1 port map( A => n5876, ZN => n6624);
   U1269 : CLKBUF_X1 port map( A => n6624, Z => n6613);
   U1270 : INV_X1 port map( A => n5877, ZN => n6570);
   U1271 : CLKBUF_X1 port map( A => n6570, Z => n6628);
   U1272 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_31_port, B1 => 
                           n6628, B2 => REGISTERS_2_31_port, ZN => n5887);
   U1273 : INV_X1 port map( A => n5878, ZN => n6474);
   U1274 : CLKBUF_X1 port map( A => n6474, Z => n6629);
   U1275 : INV_X1 port map( A => n5879, ZN => n6541);
   U1276 : CLKBUF_X1 port map( A => n6541, Z => n6331);
   U1277 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_31_port, B1 => 
                           n6331, B2 => REGISTERS_1_31_port, ZN => n5886);
   U1278 : INV_X1 port map( A => n5880, ZN => n6626);
   U1279 : CLKBUF_X1 port map( A => n6626, Z => n6618);
   U1280 : INV_X1 port map( A => n5881, ZN => n6575);
   U1281 : CLKBUF_X1 port map( A => n6575, Z => n6617);
   U1282 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_31_port, B1 => 
                           n6617, B2 => REGISTERS_3_31_port, ZN => n5885);
   U1283 : INV_X1 port map( A => n5882, ZN => n6542);
   U1284 : CLKBUF_X1 port map( A => n6542, Z => n6332);
   U1285 : INV_X1 port map( A => n5883, ZN => n6576);
   U1286 : CLKBUF_X1 port map( A => n6576, Z => n6625);
   U1287 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_31_port, B1 => 
                           n6625, B2 => REGISTERS_0_31_port, ZN => n5884);
   U1288 : NAND4_X1 port map( A1 => n5887, A2 => n5886, A3 => n5885, A4 => 
                           n5884, ZN => n5894);
   U1289 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n5888, A3 => n6586, ZN => 
                           n6636);
   U1290 : CLKBUF_X1 port map( A => n6636, Z => n6480);
   U1291 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_31_port, B1 => 
                           n6331, B2 => REGISTERS_9_31_port, ZN => n5892);
   U1292 : CLKBUF_X1 port map( A => n6575, Z => n6623);
   U1293 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_31_port, B1 => 
                           n6623, B2 => REGISTERS_11_31_port, ZN => n5891);
   U1294 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_31_port, B1 => 
                           n6625, B2 => REGISTERS_8_31_port, ZN => n5890);
   U1295 : CLKBUF_X1 port map( A => n6626, Z => n6569);
   U1296 : CLKBUF_X1 port map( A => n6624, Z => n6577);
   U1297 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_12_31_port, B1 => 
                           n6577, B2 => REGISTERS_13_31_port, ZN => n5889);
   U1298 : NAND4_X1 port map( A1 => n5892, A2 => n5891, A3 => n5890, A4 => 
                           n5889, ZN => n5893);
   U1299 : AOI22_X1 port map( A1 => n6456, A2 => n5894, B1 => n6480, B2 => 
                           n5893, ZN => n5895);
   U1300 : OAI21_X1 port map( B1 => n6586, B2 => n5896, A => n5895, ZN => N448)
                           ;
   U1301 : CLKBUF_X1 port map( A => n6369, Z => n6606);
   U1302 : CLKBUF_X1 port map( A => n6589, Z => n6388);
   U1303 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_30_port, B1 => 
                           n6388, B2 => REGISTERS_30_30_port, ZN => n5900);
   U1304 : CLKBUF_X1 port map( A => n6439, Z => n6587);
   U1305 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_30_port, B1 => 
                           n6587, B2 => REGISTERS_25_30_port, ZN => n5899);
   U1306 : CLKBUF_X1 port map( A => n6320, Z => n6591);
   U1307 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_30_port, B1 => 
                           n6561, B2 => REGISTERS_28_30_port, ZN => n5898);
   U1308 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_30_port, B1 => 
                           n6604, B2 => REGISTERS_19_30_port, ZN => n5897);
   U1309 : NAND4_X1 port map( A1 => n5900, A2 => n5899, A3 => n5898, A4 => 
                           n5897, ZN => n5906);
   U1310 : CLKBUF_X1 port map( A => n6459, Z => n6600);
   U1311 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_30_port, B1 => 
                           n6603, B2 => REGISTERS_29_30_port, ZN => n5904);
   U1312 : CLKBUF_X1 port map( A => n6416, Z => n6599);
   U1313 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_30_port, B1 => 
                           n6599, B2 => REGISTERS_17_30_port, ZN => n5903);
   U1314 : CLKBUF_X1 port map( A => n6592, Z => n6393);
   U1315 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_30_port, B1 => 
                           n6555, B2 => REGISTERS_27_30_port, ZN => n5902);
   U1316 : CLKBUF_X1 port map( A => n6364, Z => n6593);
   U1317 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_30_port, B1 => 
                           n6593, B2 => REGISTERS_23_30_port, ZN => n5901);
   U1318 : NAND4_X1 port map( A1 => n5904, A2 => n5903, A3 => n5902, A4 => 
                           n5901, ZN => n5905);
   U1319 : NOR2_X1 port map( A1 => n5906, A2 => n5905, ZN => n5918);
   U1320 : CLKBUF_X1 port map( A => n6570, Z => n6614);
   U1321 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_5_30_port, B1 => 
                           n6614, B2 => REGISTERS_2_30_port, ZN => n5910);
   U1322 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_30_port, B1 => 
                           n6331, B2 => REGISTERS_1_30_port, ZN => n5909);
   U1323 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_30_port, B1 => 
                           n6474, B2 => REGISTERS_7_30_port, ZN => n5908);
   U1324 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_30_port, B1 => 
                           n6625, B2 => REGISTERS_0_30_port, ZN => n5907);
   U1325 : NAND4_X1 port map( A1 => n5910, A2 => n5909, A3 => n5908, A4 => 
                           n5907, ZN => n5916);
   U1326 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_30_port, B1 => 
                           n6614, B2 => REGISTERS_10_30_port, ZN => n5914);
   U1327 : CLKBUF_X1 port map( A => n6576, Z => n6615);
   U1328 : CLKBUF_X1 port map( A => n6474, Z => n6616);
   U1329 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_30_port, B1 => 
                           n6616, B2 => REGISTERS_15_30_port, ZN => n5913);
   U1330 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_30_port, B1 => 
                           n6331, B2 => REGISTERS_9_30_port, ZN => n5912);
   U1331 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_30_port, B1 => 
                           n6623, B2 => REGISTERS_11_30_port, ZN => n5911);
   U1332 : NAND4_X1 port map( A1 => n5914, A2 => n5913, A3 => n5912, A4 => 
                           n5911, ZN => n5915);
   U1333 : AOI22_X1 port map( A1 => n6456, A2 => n5916, B1 => n6480, B2 => 
                           n5915, ZN => n5917);
   U1334 : OAI21_X1 port map( B1 => n6586, B2 => n5918, A => n5917, ZN => N447)
                           ;
   U1335 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_29_port, B1 => 
                           n6364, B2 => REGISTERS_23_29_port, ZN => n5922);
   U1336 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_29_port, B1 => 
                           n6315, B2 => REGISTERS_29_29_port, ZN => n5921);
   U1337 : AOI22_X1 port map( A1 => n6587, A2 => REGISTERS_25_29_port, B1 => 
                           n6388, B2 => REGISTERS_30_29_port, ZN => n5920);
   U1338 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_29_port, B1 => 
                           n6561, B2 => REGISTERS_28_29_port, ZN => n5919);
   U1339 : NAND4_X1 port map( A1 => n5922, A2 => n5921, A3 => n5920, A4 => 
                           n5919, ZN => n5928);
   U1340 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_29_port, B1 => 
                           n6459, B2 => REGISTERS_31_29_port, ZN => n5926);
   U1341 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_29_port, B1 => 
                           n6604, B2 => REGISTERS_19_29_port, ZN => n5925);
   U1342 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_29_port, B1 => 
                           n6416, B2 => REGISTERS_17_29_port, ZN => n5924);
   U1343 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_29_port, B1 => 
                           n6590, B2 => REGISTERS_27_29_port, ZN => n5923);
   U1344 : NAND4_X1 port map( A1 => n5926, A2 => n5925, A3 => n5924, A4 => 
                           n5923, ZN => n5927);
   U1345 : NOR2_X1 port map( A1 => n5928, A2 => n5927, ZN => n5940);
   U1346 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_2_29_port, B1 => 
                           n6623, B2 => REGISTERS_3_29_port, ZN => n5932);
   U1347 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_29_port, B1 => 
                           n6331, B2 => REGISTERS_1_29_port, ZN => n5931);
   U1348 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_29_port, B1 => 
                           n6625, B2 => REGISTERS_0_29_port, ZN => n5930);
   U1349 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_29_port, B1 => 
                           n6616, B2 => REGISTERS_7_29_port, ZN => n5929);
   U1350 : NAND4_X1 port map( A1 => n5932, A2 => n5931, A3 => n5930, A4 => 
                           n5929, ZN => n5938);
   U1351 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_29_port, B1 => 
                           n6625, B2 => REGISTERS_8_29_port, ZN => n5936);
   U1352 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_29_port, B1 => 
                           n6616, B2 => REGISTERS_15_29_port, ZN => n5935);
   U1353 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_11_29_port, B1 => 
                           n6331, B2 => REGISTERS_9_29_port, ZN => n5934);
   U1354 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_29_port, B1 => 
                           n6614, B2 => REGISTERS_10_29_port, ZN => n5933);
   U1355 : NAND4_X1 port map( A1 => n5936, A2 => n5935, A3 => n5934, A4 => 
                           n5933, ZN => n5937);
   U1356 : AOI22_X1 port map( A1 => n6456, A2 => n5938, B1 => n6480, B2 => 
                           n5937, ZN => n5939);
   U1357 : OAI21_X1 port map( B1 => n6586, B2 => n5940, A => n5939, ZN => N446)
                           ;
   U1358 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_28_port, B1 => 
                           n6315, B2 => REGISTERS_29_28_port, ZN => n5944);
   U1359 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_28_port, B1 => 
                           n6601, B2 => REGISTERS_18_28_port, ZN => n5943);
   U1360 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_28_port, B1 => 
                           n6341, B2 => REGISTERS_20_28_port, ZN => n5942);
   U1361 : AOI22_X1 port map( A1 => n6459, A2 => REGISTERS_31_28_port, B1 => 
                           n6416, B2 => REGISTERS_17_28_port, ZN => n5941);
   U1362 : NAND4_X1 port map( A1 => n5944, A2 => n5943, A3 => n5942, A4 => 
                           n5941, ZN => n5950);
   U1363 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_28_port, B1 => 
                           n6439, B2 => REGISTERS_25_28_port, ZN => n5948);
   U1364 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_28_port, B1 => 
                           n6604, B2 => REGISTERS_19_28_port, ZN => n5947);
   U1365 : AOI22_X1 port map( A1 => n6364, A2 => REGISTERS_23_28_port, B1 => 
                           n6388, B2 => REGISTERS_30_28_port, ZN => n5946);
   U1366 : CLKBUF_X1 port map( A => n6561, Z => n6588);
   U1367 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_28_port, B1 => 
                           n6590, B2 => REGISTERS_27_28_port, ZN => n5945);
   U1368 : NAND4_X1 port map( A1 => n5948, A2 => n5947, A3 => n5946, A4 => 
                           n5945, ZN => n5949);
   U1369 : NOR2_X1 port map( A1 => n5950, A2 => n5949, ZN => n5962);
   U1370 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_28_port, B1 => 
                           n6614, B2 => REGISTERS_2_28_port, ZN => n5954);
   U1371 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_28_port, B1 => 
                           n6624, B2 => REGISTERS_5_28_port, ZN => n5953);
   U1372 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_28_port, B1 => 
                           n6331, B2 => REGISTERS_1_28_port, ZN => n5952);
   U1373 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_28_port, B1 => 
                           n6623, B2 => REGISTERS_3_28_port, ZN => n5951);
   U1374 : NAND4_X1 port map( A1 => n5954, A2 => n5953, A3 => n5952, A4 => 
                           n5951, ZN => n5960);
   U1375 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_28_port, B1 => 
                           n6331, B2 => REGISTERS_9_28_port, ZN => n5958);
   U1376 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_28_port, B1 => 
                           n6614, B2 => REGISTERS_10_28_port, ZN => n5957);
   U1377 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_28_port, B1 => 
                           n6623, B2 => REGISTERS_11_28_port, ZN => n5956);
   U1378 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_28_port, B1 => 
                           n6616, B2 => REGISTERS_15_28_port, ZN => n5955);
   U1379 : NAND4_X1 port map( A1 => n5958, A2 => n5957, A3 => n5956, A4 => 
                           n5955, ZN => n5959);
   U1380 : AOI22_X1 port map( A1 => n6456, A2 => n5960, B1 => n6480, B2 => 
                           n5959, ZN => n5961);
   U1381 : OAI21_X1 port map( B1 => n6586, B2 => n5962, A => n5961, ZN => N445)
                           ;
   U1382 : AOI22_X1 port map( A1 => n6555, A2 => REGISTERS_27_27_port, B1 => 
                           n6364, B2 => REGISTERS_23_27_port, ZN => n5966);
   U1383 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_27_port, B1 => 
                           n6561, B2 => REGISTERS_28_27_port, ZN => n5965);
   U1384 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_27_port, B1 => 
                           n6591, B2 => REGISTERS_16_27_port, ZN => n5964);
   U1385 : AOI22_X1 port map( A1 => n6599, A2 => REGISTERS_17_27_port, B1 => 
                           n6439, B2 => REGISTERS_25_27_port, ZN => n5963);
   U1386 : NAND4_X1 port map( A1 => n5966, A2 => n5965, A3 => n5964, A4 => 
                           n5963, ZN => n5972);
   U1387 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_27_port, B1 => 
                           n6388, B2 => REGISTERS_30_27_port, ZN => n5970);
   U1388 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_27_port, B1 => 
                           n6315, B2 => REGISTERS_29_27_port, ZN => n5969);
   U1389 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_27_port, B1 => 
                           n6459, B2 => REGISTERS_31_27_port, ZN => n5968);
   U1390 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_27_port, B1 => 
                           n6341, B2 => REGISTERS_20_27_port, ZN => n5967);
   U1391 : NAND4_X1 port map( A1 => n5970, A2 => n5969, A3 => n5968, A4 => 
                           n5967, ZN => n5971);
   U1392 : NOR2_X1 port map( A1 => n5972, A2 => n5971, ZN => n5984);
   U1393 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_27_port, B1 => 
                           n6625, B2 => REGISTERS_0_27_port, ZN => n5976);
   U1394 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_2_27_port, B1 => 
                           n6331, B2 => REGISTERS_1_27_port, ZN => n5975);
   U1395 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_27_port, B1 => 
                           n6616, B2 => REGISTERS_7_27_port, ZN => n5974);
   U1396 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_5_27_port, B1 => 
                           n6575, B2 => REGISTERS_3_27_port, ZN => n5973);
   U1397 : NAND4_X1 port map( A1 => n5976, A2 => n5975, A3 => n5974, A4 => 
                           n5973, ZN => n5982);
   U1398 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_11_27_port, B1 => 
                           n6331, B2 => REGISTERS_9_27_port, ZN => n5980);
   U1399 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_27_port, B1 => 
                           n6576, B2 => REGISTERS_8_27_port, ZN => n5979);
   U1400 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_27_port, B1 => 
                           n6474, B2 => REGISTERS_15_27_port, ZN => n5978);
   U1401 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_27_port, B1 => 
                           n6570, B2 => REGISTERS_10_27_port, ZN => n5977);
   U1402 : NAND4_X1 port map( A1 => n5980, A2 => n5979, A3 => n5978, A4 => 
                           n5977, ZN => n5981);
   U1403 : AOI22_X1 port map( A1 => n6456, A2 => n5982, B1 => n6480, B2 => 
                           n5981, ZN => n5983);
   U1404 : OAI21_X1 port map( B1 => n6586, B2 => n5984, A => n5983, ZN => N444)
                           ;
   U1405 : AOI22_X1 port map( A1 => n6599, A2 => REGISTERS_17_26_port, B1 => 
                           n6439, B2 => REGISTERS_25_26_port, ZN => n5988);
   U1406 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_26_port, B1 => 
                           n6601, B2 => REGISTERS_18_26_port, ZN => n5987);
   U1407 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_26_port, B1 => 
                           n6388, B2 => REGISTERS_30_26_port, ZN => n5986);
   U1408 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_26_port, B1 => 
                           n6590, B2 => REGISTERS_27_26_port, ZN => n5985);
   U1409 : NAND4_X1 port map( A1 => n5988, A2 => n5987, A3 => n5986, A4 => 
                           n5985, ZN => n5994);
   U1410 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_26_port, B1 => 
                           n6604, B2 => REGISTERS_19_26_port, ZN => n5992);
   U1411 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_26_port, B1 => 
                           n6315, B2 => REGISTERS_29_26_port, ZN => n5991);
   U1412 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_26_port, B1 => 
                           n6364, B2 => REGISTERS_23_26_port, ZN => n5990);
   U1413 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_26_port, B1 => 
                           n6320, B2 => REGISTERS_16_26_port, ZN => n5989);
   U1414 : NAND4_X1 port map( A1 => n5992, A2 => n5991, A3 => n5990, A4 => 
                           n5989, ZN => n5993);
   U1415 : NOR2_X1 port map( A1 => n5994, A2 => n5993, ZN => n6006);
   U1416 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_26_port, B1 => 
                           n6331, B2 => REGISTERS_1_26_port, ZN => n5998);
   U1417 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_26_port, B1 => 
                           n6577, B2 => REGISTERS_5_26_port, ZN => n5997);
   U1418 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_26_port, B1 => 
                           n6623, B2 => REGISTERS_3_26_port, ZN => n5996);
   U1419 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_26_port, B1 => 
                           n6614, B2 => REGISTERS_2_26_port, ZN => n5995);
   U1420 : NAND4_X1 port map( A1 => n5998, A2 => n5997, A3 => n5996, A4 => 
                           n5995, ZN => n6004);
   U1421 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_26_port, B1 => 
                           n6570, B2 => REGISTERS_10_26_port, ZN => n6002);
   U1422 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_26_port, B1 => 
                           n6625, B2 => REGISTERS_8_26_port, ZN => n6001);
   U1423 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_12_26_port, B1 => 
                           n6575, B2 => REGISTERS_11_26_port, ZN => n6000);
   U1424 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_26_port, B1 => 
                           n6331, B2 => REGISTERS_9_26_port, ZN => n5999);
   U1425 : NAND4_X1 port map( A1 => n6002, A2 => n6001, A3 => n6000, A4 => 
                           n5999, ZN => n6003);
   U1426 : AOI22_X1 port map( A1 => n6456, A2 => n6004, B1 => n6480, B2 => 
                           n6003, ZN => n6005);
   U1427 : OAI21_X1 port map( B1 => n6586, B2 => n6006, A => n6005, ZN => N443)
                           ;
   U1428 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_25_port, B1 => 
                           n6416, B2 => REGISTERS_17_25_port, ZN => n6010);
   U1429 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_25_port, B1 => 
                           n6439, B2 => REGISTERS_25_25_port, ZN => n6009);
   U1430 : AOI22_X1 port map( A1 => n6590, A2 => REGISTERS_27_25_port, B1 => 
                           n6388, B2 => REGISTERS_30_25_port, ZN => n6008);
   U1431 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_25_port, B1 => 
                           n6364, B2 => REGISTERS_23_25_port, ZN => n6007);
   U1432 : NAND4_X1 port map( A1 => n6010, A2 => n6009, A3 => n6008, A4 => 
                           n6007, ZN => n6016);
   U1433 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_25_port, B1 => 
                           n6315, B2 => REGISTERS_29_25_port, ZN => n6014);
   U1434 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_25_port, B1 => 
                           n6459, B2 => REGISTERS_31_25_port, ZN => n6013);
   U1435 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_25_port, B1 => 
                           n6561, B2 => REGISTERS_28_25_port, ZN => n6012);
   U1436 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_25_port, B1 => 
                           n6601, B2 => REGISTERS_18_25_port, ZN => n6011);
   U1437 : NAND4_X1 port map( A1 => n6014, A2 => n6013, A3 => n6012, A4 => 
                           n6011, ZN => n6015);
   U1438 : NOR2_X1 port map( A1 => n6016, A2 => n6015, ZN => n6028);
   U1439 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_25_port, B1 => 
                           n6614, B2 => REGISTERS_2_25_port, ZN => n6020);
   U1440 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_25_port, B1 => 
                           n6331, B2 => REGISTERS_1_25_port, ZN => n6019);
   U1441 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_25_port, B1 => 
                           n6577, B2 => REGISTERS_5_25_port, ZN => n6018);
   U1442 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_25_port, B1 => 
                           n6576, B2 => REGISTERS_0_25_port, ZN => n6017);
   U1443 : NAND4_X1 port map( A1 => n6020, A2 => n6019, A3 => n6018, A4 => 
                           n6017, ZN => n6026);
   U1444 : CLKBUF_X1 port map( A => n6541, Z => n6627);
   U1445 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_11_25_port, B1 => 
                           n6627, B2 => REGISTERS_9_25_port, ZN => n6024);
   U1446 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_25_port, B1 => 
                           n6577, B2 => REGISTERS_13_25_port, ZN => n6023);
   U1447 : CLKBUF_X1 port map( A => n6542, Z => n6630);
   U1448 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_25_port, B1 => 
                           n6625, B2 => REGISTERS_8_25_port, ZN => n6022);
   U1449 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_25_port, B1 => 
                           n6570, B2 => REGISTERS_10_25_port, ZN => n6021);
   U1450 : NAND4_X1 port map( A1 => n6024, A2 => n6023, A3 => n6022, A4 => 
                           n6021, ZN => n6025);
   U1451 : AOI22_X1 port map( A1 => n6456, A2 => n6026, B1 => n6480, B2 => 
                           n6025, ZN => n6027);
   U1452 : OAI21_X1 port map( B1 => n6586, B2 => n6028, A => n6027, ZN => N442)
                           ;
   U1453 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_24_port, B1 => 
                           n6320, B2 => REGISTERS_16_24_port, ZN => n6032);
   U1454 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_24_port, B1 => 
                           n6315, B2 => REGISTERS_29_24_port, ZN => n6031);
   U1455 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_24_port, B1 => 
                           n6605, B2 => REGISTERS_24_24_port, ZN => n6030);
   U1456 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_24_port, B1 => 
                           n6590, B2 => REGISTERS_27_24_port, ZN => n6029);
   U1457 : NAND4_X1 port map( A1 => n6032, A2 => n6031, A3 => n6030, A4 => 
                           n6029, ZN => n6038);
   U1458 : AOI22_X1 port map( A1 => n6599, A2 => REGISTERS_17_24_port, B1 => 
                           n6364, B2 => REGISTERS_23_24_port, ZN => n6036);
   U1459 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_24_port, B1 => 
                           n6388, B2 => REGISTERS_30_24_port, ZN => n6035);
   U1460 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_24_port, B1 => 
                           n6439, B2 => REGISTERS_25_24_port, ZN => n6034);
   U1461 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_24_port, B1 => 
                           n6507, B2 => REGISTERS_26_24_port, ZN => n6033);
   U1462 : NAND4_X1 port map( A1 => n6036, A2 => n6035, A3 => n6034, A4 => 
                           n6033, ZN => n6037);
   U1463 : NOR2_X1 port map( A1 => n6038, A2 => n6037, ZN => n6050);
   U1464 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_7_24_port, B1 => 
                           n6614, B2 => REGISTERS_2_24_port, ZN => n6042);
   U1465 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_24_port, B1 => 
                           n6541, B2 => REGISTERS_1_24_port, ZN => n6041);
   U1466 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_24_port, B1 => 
                           n6623, B2 => REGISTERS_3_24_port, ZN => n6040);
   U1467 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_5_24_port, B1 => 
                           n6576, B2 => REGISTERS_0_24_port, ZN => n6039);
   U1468 : NAND4_X1 port map( A1 => n6042, A2 => n6041, A3 => n6040, A4 => 
                           n6039, ZN => n6048);
   U1469 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_24_port, B1 => 
                           n6331, B2 => REGISTERS_9_24_port, ZN => n6046);
   U1470 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_24_port, B1 => 
                           n6577, B2 => REGISTERS_13_24_port, ZN => n6045);
   U1471 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_24_port, B1 => 
                           n6575, B2 => REGISTERS_11_24_port, ZN => n6044);
   U1472 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_24_port, B1 => 
                           n6616, B2 => REGISTERS_15_24_port, ZN => n6043);
   U1473 : NAND4_X1 port map( A1 => n6046, A2 => n6045, A3 => n6044, A4 => 
                           n6043, ZN => n6047);
   U1474 : AOI22_X1 port map( A1 => n6456, A2 => n6048, B1 => n6480, B2 => 
                           n6047, ZN => n6049);
   U1475 : OAI21_X1 port map( B1 => n6586, B2 => n6050, A => n6049, ZN => N441)
                           ;
   U1476 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_23_port, B1 => 
                           n6588, B2 => REGISTERS_28_23_port, ZN => n6054);
   U1477 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_23_port, B1 => 
                           n6601, B2 => REGISTERS_18_23_port, ZN => n6053);
   U1478 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_23_port, B1 => 
                           n6416, B2 => REGISTERS_17_23_port, ZN => n6052);
   U1479 : CLKBUF_X1 port map( A => n6341, Z => n6602);
   U1480 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_23_port, B1 => 
                           n6315, B2 => REGISTERS_29_23_port, ZN => n6051);
   U1481 : NAND4_X1 port map( A1 => n6054, A2 => n6053, A3 => n6052, A4 => 
                           n6051, ZN => n6060);
   U1482 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_23_port, B1 => 
                           n6439, B2 => REGISTERS_25_23_port, ZN => n6058);
   U1483 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_23_port, B1 => 
                           n6507, B2 => REGISTERS_26_23_port, ZN => n6057);
   U1484 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_23_port, B1 => 
                           n6388, B2 => REGISTERS_30_23_port, ZN => n6056);
   U1485 : AOI22_X1 port map( A1 => n6555, A2 => REGISTERS_27_23_port, B1 => 
                           n6364, B2 => REGISTERS_23_23_port, ZN => n6055);
   U1486 : NAND4_X1 port map( A1 => n6058, A2 => n6057, A3 => n6056, A4 => 
                           n6055, ZN => n6059);
   U1487 : NOR2_X1 port map( A1 => n6060, A2 => n6059, ZN => n6072);
   U1488 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_23_port, B1 => 
                           n6474, B2 => REGISTERS_7_23_port, ZN => n6064);
   U1489 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_23_port, B1 => 
                           n6623, B2 => REGISTERS_3_23_port, ZN => n6063);
   U1490 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_23_port, B1 => 
                           n6627, B2 => REGISTERS_1_23_port, ZN => n6062);
   U1491 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_23_port, B1 => 
                           n6570, B2 => REGISTERS_2_23_port, ZN => n6061);
   U1492 : NAND4_X1 port map( A1 => n6064, A2 => n6063, A3 => n6062, A4 => 
                           n6061, ZN => n6070);
   U1493 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_23_port, B1 => 
                           n6616, B2 => REGISTERS_15_23_port, ZN => n6068);
   U1494 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_23_port, B1 => 
                           n6625, B2 => REGISTERS_8_23_port, ZN => n6067);
   U1495 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_23_port, B1 => 
                           n6541, B2 => REGISTERS_9_23_port, ZN => n6066);
   U1496 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_23_port, B1 => 
                           n6575, B2 => REGISTERS_11_23_port, ZN => n6065);
   U1497 : NAND4_X1 port map( A1 => n6068, A2 => n6067, A3 => n6066, A4 => 
                           n6065, ZN => n6069);
   U1498 : AOI22_X1 port map( A1 => n6456, A2 => n6070, B1 => n6480, B2 => 
                           n6069, ZN => n6071);
   U1499 : OAI21_X1 port map( B1 => n6641, B2 => n6072, A => n6071, ZN => N440)
                           ;
   U1500 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_22_port, B1 => 
                           n6439, B2 => REGISTERS_25_22_port, ZN => n6076);
   U1501 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_22_port, B1 => 
                           n6560, B2 => REGISTERS_18_22_port, ZN => n6075);
   U1502 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_22_port, B1 => 
                           n6315, B2 => REGISTERS_29_22_port, ZN => n6074);
   U1503 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_22_port, B1 => 
                           n6590, B2 => REGISTERS_27_22_port, ZN => n6073);
   U1504 : NAND4_X1 port map( A1 => n6076, A2 => n6075, A3 => n6074, A4 => 
                           n6073, ZN => n6082);
   U1505 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_22_port, B1 => 
                           n6588, B2 => REGISTERS_28_22_port, ZN => n6080);
   U1506 : AOI22_X1 port map( A1 => n6593, A2 => REGISTERS_23_22_port, B1 => 
                           n6388, B2 => REGISTERS_30_22_port, ZN => n6079);
   U1507 : AOI22_X1 port map( A1 => n6507, A2 => REGISTERS_26_22_port, B1 => 
                           n6416, B2 => REGISTERS_17_22_port, ZN => n6078);
   U1508 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_22_port, B1 => 
                           n6562, B2 => REGISTERS_19_22_port, ZN => n6077);
   U1509 : NAND4_X1 port map( A1 => n6080, A2 => n6079, A3 => n6078, A4 => 
                           n6077, ZN => n6081);
   U1510 : NOR2_X1 port map( A1 => n6082, A2 => n6081, ZN => n6094);
   U1511 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_22_port, B1 => 
                           n6331, B2 => REGISTERS_1_22_port, ZN => n6086);
   U1512 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_22_port, B1 => 
                           n6624, B2 => REGISTERS_5_22_port, ZN => n6085);
   U1513 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_22_port, B1 => 
                           n6474, B2 => REGISTERS_7_22_port, ZN => n6084);
   U1514 : AOI22_X1 port map( A1 => n6625, A2 => REGISTERS_0_22_port, B1 => 
                           n6614, B2 => REGISTERS_2_22_port, ZN => n6083);
   U1515 : NAND4_X1 port map( A1 => n6086, A2 => n6085, A3 => n6084, A4 => 
                           n6083, ZN => n6092);
   U1516 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_22_port, B1 => 
                           n6570, B2 => REGISTERS_10_22_port, ZN => n6090);
   U1517 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_22_port, B1 => 
                           n6616, B2 => REGISTERS_15_22_port, ZN => n6089);
   U1518 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_22_port, B1 => 
                           n6613, B2 => REGISTERS_13_22_port, ZN => n6088);
   U1519 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_11_22_port, B1 => 
                           n6627, B2 => REGISTERS_9_22_port, ZN => n6087);
   U1520 : NAND4_X1 port map( A1 => n6090, A2 => n6089, A3 => n6088, A4 => 
                           n6087, ZN => n6091);
   U1521 : AOI22_X1 port map( A1 => n6456, A2 => n6092, B1 => n6480, B2 => 
                           n6091, ZN => n6093);
   U1522 : OAI21_X1 port map( B1 => n6641, B2 => n6094, A => n6093, ZN => N439)
                           ;
   U1523 : AOI22_X1 port map( A1 => n6601, A2 => REGISTERS_18_21_port, B1 => 
                           n6561, B2 => REGISTERS_28_21_port, ZN => n6098);
   U1524 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_21_port, B1 => 
                           n6507, B2 => REGISTERS_26_21_port, ZN => n6097);
   U1525 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_21_port, B1 => 
                           n6416, B2 => REGISTERS_17_21_port, ZN => n6096);
   U1526 : AOI22_X1 port map( A1 => n6555, A2 => REGISTERS_27_21_port, B1 => 
                           n6589, B2 => REGISTERS_30_21_port, ZN => n6095);
   U1527 : NAND4_X1 port map( A1 => n6098, A2 => n6097, A3 => n6096, A4 => 
                           n6095, ZN => n6104);
   U1528 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_21_port, B1 => 
                           n6364, B2 => REGISTERS_23_21_port, ZN => n6102);
   U1529 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_21_port, B1 => 
                           n6439, B2 => REGISTERS_25_21_port, ZN => n6101);
   U1530 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_21_port, B1 => 
                           n6369, B2 => REGISTERS_21_21_port, ZN => n6100);
   U1531 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_21_port, B1 => 
                           n6603, B2 => REGISTERS_29_21_port, ZN => n6099);
   U1532 : NAND4_X1 port map( A1 => n6102, A2 => n6101, A3 => n6100, A4 => 
                           n6099, ZN => n6103);
   U1533 : NOR2_X1 port map( A1 => n6104, A2 => n6103, ZN => n6116);
   U1534 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_0_21_port, B1 => 
                           n6474, B2 => REGISTERS_7_21_port, ZN => n6108);
   U1535 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_21_port, B1 => 
                           n6541, B2 => REGISTERS_1_21_port, ZN => n6107);
   U1536 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_21_port, B1 => 
                           n6614, B2 => REGISTERS_2_21_port, ZN => n6106);
   U1537 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_21_port, B1 => 
                           n6623, B2 => REGISTERS_3_21_port, ZN => n6105);
   U1538 : NAND4_X1 port map( A1 => n6108, A2 => n6107, A3 => n6106, A4 => 
                           n6105, ZN => n6114);
   U1539 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_21_port, B1 => 
                           n6331, B2 => REGISTERS_9_21_port, ZN => n6112);
   U1540 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_21_port, B1 => 
                           n6575, B2 => REGISTERS_11_21_port, ZN => n6111);
   U1541 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_21_port, B1 => 
                           n6626, B2 => REGISTERS_12_21_port, ZN => n6110);
   U1542 : AOI22_X1 port map( A1 => n6625, A2 => REGISTERS_8_21_port, B1 => 
                           n6570, B2 => REGISTERS_10_21_port, ZN => n6109);
   U1543 : NAND4_X1 port map( A1 => n6112, A2 => n6111, A3 => n6110, A4 => 
                           n6109, ZN => n6113);
   U1544 : AOI22_X1 port map( A1 => n6456, A2 => n6114, B1 => n6480, B2 => 
                           n6113, ZN => n6115);
   U1545 : OAI21_X1 port map( B1 => n6641, B2 => n6116, A => n6115, ZN => N438)
                           ;
   U1546 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_20_port, B1 => 
                           n6560, B2 => REGISTERS_18_20_port, ZN => n6120);
   U1547 : AOI22_X1 port map( A1 => n6561, A2 => REGISTERS_28_20_port, B1 => 
                           n6587, B2 => REGISTERS_25_20_port, ZN => n6119);
   U1548 : AOI22_X1 port map( A1 => n6604, A2 => REGISTERS_19_20_port, B1 => 
                           n6416, B2 => REGISTERS_17_20_port, ZN => n6118);
   U1549 : AOI22_X1 port map( A1 => n6603, A2 => REGISTERS_29_20_port, B1 => 
                           n6590, B2 => REGISTERS_27_20_port, ZN => n6117);
   U1550 : NAND4_X1 port map( A1 => n6120, A2 => n6119, A3 => n6118, A4 => 
                           n6117, ZN => n6126);
   U1551 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_20_port, B1 => 
                           n6589, B2 => REGISTERS_30_20_port, ZN => n6124);
   U1552 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_20_port, B1 => 
                           n6507, B2 => REGISTERS_26_20_port, ZN => n6123);
   U1553 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_20_port, B1 => 
                           n6320, B2 => REGISTERS_16_20_port, ZN => n6122);
   U1554 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_20_port, B1 => 
                           n6364, B2 => REGISTERS_23_20_port, ZN => n6121);
   U1555 : NAND4_X1 port map( A1 => n6124, A2 => n6123, A3 => n6122, A4 => 
                           n6121, ZN => n6125);
   U1556 : NOR2_X1 port map( A1 => n6126, A2 => n6125, ZN => n6138);
   U1557 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_20_port, B1 => 
                           n6623, B2 => REGISTERS_3_20_port, ZN => n6130);
   U1558 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_2_20_port, B1 => 
                           n6627, B2 => REGISTERS_1_20_port, ZN => n6129);
   U1559 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_20_port, B1 => 
                           n6569, B2 => REGISTERS_4_20_port, ZN => n6128);
   U1560 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_5_20_port, B1 => 
                           n6576, B2 => REGISTERS_0_20_port, ZN => n6127);
   U1561 : NAND4_X1 port map( A1 => n6130, A2 => n6129, A3 => n6128, A4 => 
                           n6127, ZN => n6136);
   U1562 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_20_port, B1 => 
                           n6575, B2 => REGISTERS_11_20_port, ZN => n6134);
   U1563 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_8_20_port, B1 => 
                           n6570, B2 => REGISTERS_10_20_port, ZN => n6133);
   U1564 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_20_port, B1 => 
                           n6577, B2 => REGISTERS_13_20_port, ZN => n6132);
   U1565 : AOI22_X1 port map( A1 => n6616, A2 => REGISTERS_15_20_port, B1 => 
                           n6541, B2 => REGISTERS_9_20_port, ZN => n6131);
   U1566 : NAND4_X1 port map( A1 => n6134, A2 => n6133, A3 => n6132, A4 => 
                           n6131, ZN => n6135);
   U1567 : AOI22_X1 port map( A1 => n6456, A2 => n6136, B1 => n6636, B2 => 
                           n6135, ZN => n6137);
   U1568 : OAI21_X1 port map( B1 => n6641, B2 => n6138, A => n6137, ZN => N437)
                           ;
   U1569 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_19_port, B1 => 
                           n6388, B2 => REGISTERS_30_19_port, ZN => n6142);
   U1570 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_19_port, B1 => 
                           n6416, B2 => REGISTERS_17_19_port, ZN => n6141);
   U1571 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_19_port, B1 => 
                           n6593, B2 => REGISTERS_23_19_port, ZN => n6140);
   U1572 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_19_port, B1 => 
                           n6562, B2 => REGISTERS_19_19_port, ZN => n6139);
   U1573 : NAND4_X1 port map( A1 => n6142, A2 => n6141, A3 => n6140, A4 => 
                           n6139, ZN => n6148);
   U1574 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_19_port, B1 => 
                           n6560, B2 => REGISTERS_18_19_port, ZN => n6146);
   U1575 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_19_port, B1 => 
                           n6603, B2 => REGISTERS_29_19_port, ZN => n6145);
   U1576 : AOI22_X1 port map( A1 => n6561, A2 => REGISTERS_28_19_port, B1 => 
                           n6590, B2 => REGISTERS_27_19_port, ZN => n6144);
   U1577 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_19_port, B1 => 
                           n6587, B2 => REGISTERS_25_19_port, ZN => n6143);
   U1578 : NAND4_X1 port map( A1 => n6146, A2 => n6145, A3 => n6144, A4 => 
                           n6143, ZN => n6147);
   U1579 : NOR2_X1 port map( A1 => n6148, A2 => n6147, ZN => n6160);
   U1580 : CLKBUF_X1 port map( A => n6638, Z => n6482);
   U1581 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_19_port, B1 => 
                           n6614, B2 => REGISTERS_2_19_port, ZN => n6152);
   U1582 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_19_port, B1 => 
                           n6616, B2 => REGISTERS_7_19_port, ZN => n6151);
   U1583 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_19_port, B1 => 
                           n6569, B2 => REGISTERS_4_19_port, ZN => n6150);
   U1584 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_19_port, B1 => 
                           n6331, B2 => REGISTERS_1_19_port, ZN => n6149);
   U1585 : NAND4_X1 port map( A1 => n6152, A2 => n6151, A3 => n6150, A4 => 
                           n6149, ZN => n6158);
   U1586 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_19_port, B1 => 
                           n6570, B2 => REGISTERS_10_19_port, ZN => n6156);
   U1587 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_19_port, B1 => 
                           n6575, B2 => REGISTERS_11_19_port, ZN => n6155);
   U1588 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_19_port, B1 => 
                           n6627, B2 => REGISTERS_9_19_port, ZN => n6154);
   U1589 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_19_port, B1 => 
                           n6474, B2 => REGISTERS_15_19_port, ZN => n6153);
   U1590 : NAND4_X1 port map( A1 => n6156, A2 => n6155, A3 => n6154, A4 => 
                           n6153, ZN => n6157);
   U1591 : AOI22_X1 port map( A1 => n6482, A2 => n6158, B1 => n6480, B2 => 
                           n6157, ZN => n6159);
   U1592 : OAI21_X1 port map( B1 => n6641, B2 => n6160, A => n6159, ZN => N436)
                           ;
   U1593 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_18_port, B1 => 
                           n6590, B2 => REGISTERS_27_18_port, ZN => n6164);
   U1594 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_18_port, B1 => 
                           n6603, B2 => REGISTERS_29_18_port, ZN => n6163);
   U1595 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_18_port, B1 => 
                           n6599, B2 => REGISTERS_17_18_port, ZN => n6162);
   U1596 : AOI22_X1 port map( A1 => n6320, A2 => REGISTERS_16_18_port, B1 => 
                           n6593, B2 => REGISTERS_23_18_port, ZN => n6161);
   U1597 : NAND4_X1 port map( A1 => n6164, A2 => n6163, A3 => n6162, A4 => 
                           n6161, ZN => n6170);
   U1598 : AOI22_X1 port map( A1 => n6605, A2 => REGISTERS_24_18_port, B1 => 
                           n6560, B2 => REGISTERS_18_18_port, ZN => n6168);
   U1599 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_18_port, B1 => 
                           n6459, B2 => REGISTERS_31_18_port, ZN => n6167);
   U1600 : AOI22_X1 port map( A1 => n6604, A2 => REGISTERS_19_18_port, B1 => 
                           n6388, B2 => REGISTERS_30_18_port, ZN => n6166);
   U1601 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_18_port, B1 => 
                           n6587, B2 => REGISTERS_25_18_port, ZN => n6165);
   U1602 : NAND4_X1 port map( A1 => n6168, A2 => n6167, A3 => n6166, A4 => 
                           n6165, ZN => n6169);
   U1603 : NOR2_X1 port map( A1 => n6170, A2 => n6169, ZN => n6182);
   U1604 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_18_port, B1 => 
                           n6625, B2 => REGISTERS_0_18_port, ZN => n6174);
   U1605 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_18_port, B1 => 
                           n6616, B2 => REGISTERS_7_18_port, ZN => n6173);
   U1606 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_18_port, B1 => 
                           n6623, B2 => REGISTERS_3_18_port, ZN => n6172);
   U1607 : AOI22_X1 port map( A1 => n6570, A2 => REGISTERS_2_18_port, B1 => 
                           n6541, B2 => REGISTERS_1_18_port, ZN => n6171);
   U1608 : NAND4_X1 port map( A1 => n6174, A2 => n6173, A3 => n6172, A4 => 
                           n6171, ZN => n6180);
   U1609 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_18_port, B1 => 
                           n6331, B2 => REGISTERS_9_18_port, ZN => n6178);
   U1610 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_18_port, B1 => 
                           n6576, B2 => REGISTERS_8_18_port, ZN => n6177);
   U1611 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_18_port, B1 => 
                           n6575, B2 => REGISTERS_11_18_port, ZN => n6176);
   U1612 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_18_port, B1 => 
                           n6474, B2 => REGISTERS_15_18_port, ZN => n6175);
   U1613 : NAND4_X1 port map( A1 => n6178, A2 => n6177, A3 => n6176, A4 => 
                           n6175, ZN => n6179);
   U1614 : AOI22_X1 port map( A1 => n6482, A2 => n6180, B1 => n6480, B2 => 
                           n6179, ZN => n6181);
   U1615 : OAI21_X1 port map( B1 => n6641, B2 => n6182, A => n6181, ZN => N435)
                           ;
   U1616 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_17_port, B1 => 
                           n6599, B2 => REGISTERS_17_17_port, ZN => n6186);
   U1617 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_17_port, B1 => 
                           n6320, B2 => REGISTERS_16_17_port, ZN => n6185);
   U1618 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_17_port, B1 => 
                           n6555, B2 => REGISTERS_27_17_port, ZN => n6184);
   U1619 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_17_port, B1 => 
                           n6388, B2 => REGISTERS_30_17_port, ZN => n6183);
   U1620 : NAND4_X1 port map( A1 => n6186, A2 => n6185, A3 => n6184, A4 => 
                           n6183, ZN => n6192);
   U1621 : AOI22_X1 port map( A1 => n6439, A2 => REGISTERS_25_17_port, B1 => 
                           n6593, B2 => REGISTERS_23_17_port, ZN => n6190);
   U1622 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_17_port, B1 => 
                           n6603, B2 => REGISTERS_29_17_port, ZN => n6189);
   U1623 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_17_port, B1 => 
                           n6507, B2 => REGISTERS_26_17_port, ZN => n6188);
   U1624 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_17_port, B1 => 
                           n6605, B2 => REGISTERS_24_17_port, ZN => n6187);
   U1625 : NAND4_X1 port map( A1 => n6190, A2 => n6189, A3 => n6188, A4 => 
                           n6187, ZN => n6191);
   U1626 : NOR2_X1 port map( A1 => n6192, A2 => n6191, ZN => n6204);
   U1627 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_17_port, B1 => 
                           n6577, B2 => REGISTERS_5_17_port, ZN => n6196);
   U1628 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_17_port, B1 => 
                           n6474, B2 => REGISTERS_7_17_port, ZN => n6195);
   U1629 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_17_port, B1 => 
                           n6331, B2 => REGISTERS_1_17_port, ZN => n6194);
   U1630 : AOI22_X1 port map( A1 => n6625, A2 => REGISTERS_0_17_port, B1 => 
                           n6614, B2 => REGISTERS_2_17_port, ZN => n6193);
   U1631 : NAND4_X1 port map( A1 => n6196, A2 => n6195, A3 => n6194, A4 => 
                           n6193, ZN => n6202);
   U1632 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_17_port, B1 => 
                           n6625, B2 => REGISTERS_8_17_port, ZN => n6200);
   U1633 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_17_port, B1 => 
                           n6570, B2 => REGISTERS_10_17_port, ZN => n6199);
   U1634 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_17_port, B1 => 
                           n6627, B2 => REGISTERS_9_17_port, ZN => n6198);
   U1635 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_17_port, B1 => 
                           n6623, B2 => REGISTERS_11_17_port, ZN => n6197);
   U1636 : NAND4_X1 port map( A1 => n6200, A2 => n6199, A3 => n6198, A4 => 
                           n6197, ZN => n6201);
   U1637 : AOI22_X1 port map( A1 => n6482, A2 => n6202, B1 => n6480, B2 => 
                           n6201, ZN => n6203);
   U1638 : OAI21_X1 port map( B1 => n6641, B2 => n6204, A => n6203, ZN => N434)
                           ;
   U1639 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_16_port, B1 => 
                           n6605, B2 => REGISTERS_24_16_port, ZN => n6208);
   U1640 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_16_port, B1 => 
                           n6593, B2 => REGISTERS_23_16_port, ZN => n6207);
   U1641 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_16_port, B1 => 
                           n6388, B2 => REGISTERS_30_16_port, ZN => n6206);
   U1642 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_16_port, B1 => 
                           n6599, B2 => REGISTERS_17_16_port, ZN => n6205);
   U1643 : NAND4_X1 port map( A1 => n6208, A2 => n6207, A3 => n6206, A4 => 
                           n6205, ZN => n6214);
   U1644 : AOI22_X1 port map( A1 => n6315, A2 => REGISTERS_29_16_port, B1 => 
                           n6587, B2 => REGISTERS_25_16_port, ZN => n6212);
   U1645 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_16_port, B1 => 
                           n6320, B2 => REGISTERS_16_16_port, ZN => n6211);
   U1646 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_16_port, B1 => 
                           n6507, B2 => REGISTERS_26_16_port, ZN => n6210);
   U1647 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_16_port, B1 => 
                           n6555, B2 => REGISTERS_27_16_port, ZN => n6209);
   U1648 : NAND4_X1 port map( A1 => n6212, A2 => n6211, A3 => n6210, A4 => 
                           n6209, ZN => n6213);
   U1649 : NOR2_X1 port map( A1 => n6214, A2 => n6213, ZN => n6226);
   U1650 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_16_port, B1 => 
                           n6541, B2 => REGISTERS_1_16_port, ZN => n6218);
   U1651 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_16_port, B1 => 
                           n6576, B2 => REGISTERS_0_16_port, ZN => n6217);
   U1652 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_16_port, B1 => 
                           n6575, B2 => REGISTERS_3_16_port, ZN => n6216);
   U1653 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_16_port, B1 => 
                           n6614, B2 => REGISTERS_2_16_port, ZN => n6215);
   U1654 : NAND4_X1 port map( A1 => n6218, A2 => n6217, A3 => n6216, A4 => 
                           n6215, ZN => n6224);
   U1655 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_16_port, B1 => 
                           n6616, B2 => REGISTERS_15_16_port, ZN => n6222);
   U1656 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_8_16_port, B1 => 
                           n6627, B2 => REGISTERS_9_16_port, ZN => n6221);
   U1657 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_12_16_port, B1 => 
                           n6570, B2 => REGISTERS_10_16_port, ZN => n6220);
   U1658 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_16_port, B1 => 
                           n6623, B2 => REGISTERS_11_16_port, ZN => n6219);
   U1659 : NAND4_X1 port map( A1 => n6222, A2 => n6221, A3 => n6220, A4 => 
                           n6219, ZN => n6223);
   U1660 : AOI22_X1 port map( A1 => n6482, A2 => n6224, B1 => n6480, B2 => 
                           n6223, ZN => n6225);
   U1661 : OAI21_X1 port map( B1 => n6641, B2 => n6226, A => n6225, ZN => N433)
                           ;
   U1662 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_15_port, B1 => 
                           n6587, B2 => REGISTERS_25_15_port, ZN => n6230);
   U1663 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_15_port, B1 => 
                           n6562, B2 => REGISTERS_19_15_port, ZN => n6229);
   U1664 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_15_port, B1 => 
                           n6588, B2 => REGISTERS_28_15_port, ZN => n6228);
   U1665 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_15_port, B1 => 
                           n6599, B2 => REGISTERS_17_15_port, ZN => n6227);
   U1666 : NAND4_X1 port map( A1 => n6230, A2 => n6229, A3 => n6228, A4 => 
                           n6227, ZN => n6236);
   U1667 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_15_port, B1 => 
                           n6593, B2 => REGISTERS_23_15_port, ZN => n6234);
   U1668 : AOI22_X1 port map( A1 => n6605, A2 => REGISTERS_24_15_port, B1 => 
                           n6320, B2 => REGISTERS_16_15_port, ZN => n6233);
   U1669 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_15_port, B1 => 
                           n6555, B2 => REGISTERS_27_15_port, ZN => n6232);
   U1670 : AOI22_X1 port map( A1 => n6315, A2 => REGISTERS_29_15_port, B1 => 
                           n6388, B2 => REGISTERS_30_15_port, ZN => n6231);
   U1671 : NAND4_X1 port map( A1 => n6234, A2 => n6233, A3 => n6232, A4 => 
                           n6231, ZN => n6235);
   U1672 : NOR2_X1 port map( A1 => n6236, A2 => n6235, ZN => n6248);
   U1673 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_15_port, B1 => 
                           n6575, B2 => REGISTERS_3_15_port, ZN => n6240);
   U1674 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_5_15_port, B1 => 
                           n6576, B2 => REGISTERS_0_15_port, ZN => n6239);
   U1675 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_15_port, B1 => 
                           n6331, B2 => REGISTERS_1_15_port, ZN => n6238);
   U1676 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_15_port, B1 => 
                           n6628, B2 => REGISTERS_2_15_port, ZN => n6237);
   U1677 : NAND4_X1 port map( A1 => n6240, A2 => n6239, A3 => n6238, A4 => 
                           n6237, ZN => n6246);
   U1678 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_15_15_port, B1 => 
                           n6627, B2 => REGISTERS_9_15_port, ZN => n6244);
   U1679 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_15_port, B1 => 
                           n6625, B2 => REGISTERS_8_15_port, ZN => n6243);
   U1680 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_13_15_port, B1 => 
                           n6617, B2 => REGISTERS_11_15_port, ZN => n6242);
   U1681 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_15_port, B1 => 
                           n6628, B2 => REGISTERS_10_15_port, ZN => n6241);
   U1682 : NAND4_X1 port map( A1 => n6244, A2 => n6243, A3 => n6242, A4 => 
                           n6241, ZN => n6245);
   U1683 : AOI22_X1 port map( A1 => n6482, A2 => n6246, B1 => n6480, B2 => 
                           n6245, ZN => n6247);
   U1684 : OAI21_X1 port map( B1 => n6586, B2 => n6248, A => n6247, ZN => N432)
                           ;
   U1685 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_14_port, B1 => 
                           n6587, B2 => REGISTERS_25_14_port, ZN => n6252);
   U1686 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_14_port, B1 => 
                           n6507, B2 => REGISTERS_26_14_port, ZN => n6251);
   U1687 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_14_port, B1 => 
                           n6588, B2 => REGISTERS_28_14_port, ZN => n6250);
   U1688 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_14_port, B1 => 
                           n6603, B2 => REGISTERS_29_14_port, ZN => n6249);
   U1689 : NAND4_X1 port map( A1 => n6252, A2 => n6251, A3 => n6250, A4 => 
                           n6249, ZN => n6258);
   U1690 : AOI22_X1 port map( A1 => n6605, A2 => REGISTERS_24_14_port, B1 => 
                           n6593, B2 => REGISTERS_23_14_port, ZN => n6256);
   U1691 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_14_port, B1 => 
                           n6320, B2 => REGISTERS_16_14_port, ZN => n6255);
   U1692 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_14_port, B1 => 
                           n6388, B2 => REGISTERS_30_14_port, ZN => n6254);
   U1693 : AOI22_X1 port map( A1 => n6599, A2 => REGISTERS_17_14_port, B1 => 
                           n6555, B2 => REGISTERS_27_14_port, ZN => n6253);
   U1694 : NAND4_X1 port map( A1 => n6256, A2 => n6255, A3 => n6254, A4 => 
                           n6253, ZN => n6257);
   U1695 : NOR2_X1 port map( A1 => n6258, A2 => n6257, ZN => n6270);
   U1696 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_0_14_port, B1 => 
                           n6541, B2 => REGISTERS_1_14_port, ZN => n6262);
   U1697 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_14_port, B1 => 
                           n6617, B2 => REGISTERS_3_14_port, ZN => n6261);
   U1698 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_5_14_port, B1 => 
                           n6570, B2 => REGISTERS_2_14_port, ZN => n6260);
   U1699 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_14_port, B1 => 
                           n6474, B2 => REGISTERS_7_14_port, ZN => n6259);
   U1700 : NAND4_X1 port map( A1 => n6262, A2 => n6261, A3 => n6260, A4 => 
                           n6259, ZN => n6268);
   U1701 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_14_port, B1 => 
                           n6575, B2 => REGISTERS_11_14_port, ZN => n6266);
   U1702 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_12_14_port, B1 => 
                           n6576, B2 => REGISTERS_8_14_port, ZN => n6265);
   U1703 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_14_port, B1 => 
                           n6541, B2 => REGISTERS_9_14_port, ZN => n6264);
   U1704 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_14_port, B1 => 
                           n6614, B2 => REGISTERS_10_14_port, ZN => n6263);
   U1705 : NAND4_X1 port map( A1 => n6266, A2 => n6265, A3 => n6264, A4 => 
                           n6263, ZN => n6267);
   U1706 : AOI22_X1 port map( A1 => n6482, A2 => n6268, B1 => n6480, B2 => 
                           n6267, ZN => n6269);
   U1707 : OAI21_X1 port map( B1 => n6641, B2 => n6270, A => n6269, ZN => N431)
                           ;
   U1708 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_13_port, B1 => 
                           n6555, B2 => REGISTERS_27_13_port, ZN => n6274);
   U1709 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_13_port, B1 => 
                           n6587, B2 => REGISTERS_25_13_port, ZN => n6273);
   U1710 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_13_port, B1 => 
                           n6388, B2 => REGISTERS_30_13_port, ZN => n6272);
   U1711 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_13_port, B1 => 
                           n6588, B2 => REGISTERS_28_13_port, ZN => n6271);
   U1712 : NAND4_X1 port map( A1 => n6274, A2 => n6273, A3 => n6272, A4 => 
                           n6271, ZN => n6280);
   U1713 : AOI22_X1 port map( A1 => n6320, A2 => REGISTERS_16_13_port, B1 => 
                           n6593, B2 => REGISTERS_23_13_port, ZN => n6278);
   U1714 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_13_port, B1 => 
                           n6603, B2 => REGISTERS_29_13_port, ZN => n6277);
   U1715 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_13_port, B1 => 
                           n6459, B2 => REGISTERS_31_13_port, ZN => n6276);
   U1716 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_13_port, B1 => 
                           n6599, B2 => REGISTERS_17_13_port, ZN => n6275);
   U1717 : NAND4_X1 port map( A1 => n6278, A2 => n6277, A3 => n6276, A4 => 
                           n6275, ZN => n6279);
   U1718 : NOR2_X1 port map( A1 => n6280, A2 => n6279, ZN => n6292);
   U1719 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_13_port, B1 => 
                           n6570, B2 => REGISTERS_2_13_port, ZN => n6284);
   U1720 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_13_port, B1 => 
                           n6624, B2 => REGISTERS_5_13_port, ZN => n6283);
   U1721 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_13_port, B1 => 
                           n6331, B2 => REGISTERS_1_13_port, ZN => n6282);
   U1722 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_6_13_port, B1 => 
                           n6616, B2 => REGISTERS_7_13_port, ZN => n6281);
   U1723 : NAND4_X1 port map( A1 => n6284, A2 => n6283, A3 => n6282, A4 => 
                           n6281, ZN => n6290);
   U1724 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_13_port, B1 => 
                           n6625, B2 => REGISTERS_8_13_port, ZN => n6288);
   U1725 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_15_13_port, B1 => 
                           n6628, B2 => REGISTERS_10_13_port, ZN => n6287);
   U1726 : AOI22_X1 port map( A1 => n6575, A2 => REGISTERS_11_13_port, B1 => 
                           n6627, B2 => REGISTERS_9_13_port, ZN => n6286);
   U1727 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_13_port, B1 => 
                           n6624, B2 => REGISTERS_13_13_port, ZN => n6285);
   U1728 : NAND4_X1 port map( A1 => n6288, A2 => n6287, A3 => n6286, A4 => 
                           n6285, ZN => n6289);
   U1729 : AOI22_X1 port map( A1 => n6482, A2 => n6290, B1 => n6480, B2 => 
                           n6289, ZN => n6291);
   U1730 : OAI21_X1 port map( B1 => n6586, B2 => n6292, A => n6291, ZN => N430)
                           ;
   U1731 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_12_port, B1 => 
                           n6562, B2 => REGISTERS_19_12_port, ZN => n6296);
   U1732 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_12_port, B1 => 
                           n6593, B2 => REGISTERS_23_12_port, ZN => n6295);
   U1733 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_12_port, B1 => 
                           n6588, B2 => REGISTERS_28_12_port, ZN => n6294);
   U1734 : AOI22_X1 port map( A1 => n6459, A2 => REGISTERS_31_12_port, B1 => 
                           n6555, B2 => REGISTERS_27_12_port, ZN => n6293);
   U1735 : NAND4_X1 port map( A1 => n6296, A2 => n6295, A3 => n6294, A4 => 
                           n6293, ZN => n6302);
   U1736 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_12_port, B1 => 
                           n6603, B2 => REGISTERS_29_12_port, ZN => n6300);
   U1737 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_12_port, B1 => 
                           n6388, B2 => REGISTERS_30_12_port, ZN => n6299);
   U1738 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_12_port, B1 => 
                           n6587, B2 => REGISTERS_25_12_port, ZN => n6298);
   U1739 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_12_port, B1 => 
                           n6599, B2 => REGISTERS_17_12_port, ZN => n6297);
   U1740 : NAND4_X1 port map( A1 => n6300, A2 => n6299, A3 => n6298, A4 => 
                           n6297, ZN => n6301);
   U1741 : NOR2_X1 port map( A1 => n6302, A2 => n6301, ZN => n6314);
   U1742 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_12_port, B1 => 
                           n6576, B2 => REGISTERS_0_12_port, ZN => n6306);
   U1743 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_12_port, B1 => 
                           n6474, B2 => REGISTERS_7_12_port, ZN => n6305);
   U1744 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_2_12_port, B1 => 
                           n6575, B2 => REGISTERS_3_12_port, ZN => n6304);
   U1745 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_12_port, B1 => 
                           n6541, B2 => REGISTERS_1_12_port, ZN => n6303);
   U1746 : NAND4_X1 port map( A1 => n6306, A2 => n6305, A3 => n6304, A4 => 
                           n6303, ZN => n6312);
   U1747 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_12_port, B1 => 
                           n6625, B2 => REGISTERS_8_12_port, ZN => n6310);
   U1748 : AOI22_X1 port map( A1 => n6570, A2 => REGISTERS_10_12_port, B1 => 
                           n6541, B2 => REGISTERS_9_12_port, ZN => n6309);
   U1749 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_12_port, B1 => 
                           n6617, B2 => REGISTERS_11_12_port, ZN => n6308);
   U1750 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_12_port, B1 => 
                           n6616, B2 => REGISTERS_15_12_port, ZN => n6307);
   U1751 : NAND4_X1 port map( A1 => n6310, A2 => n6309, A3 => n6308, A4 => 
                           n6307, ZN => n6311);
   U1752 : AOI22_X1 port map( A1 => n6482, A2 => n6312, B1 => n6480, B2 => 
                           n6311, ZN => n6313);
   U1753 : OAI21_X1 port map( B1 => n6641, B2 => n6314, A => n6313, ZN => N429)
                           ;
   U1754 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_11_port, B1 => 
                           n6594, B2 => REGISTERS_26_11_port, ZN => n6319);
   U1755 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_11_port, B1 => 
                           n6562, B2 => REGISTERS_19_11_port, ZN => n6318);
   U1756 : AOI22_X1 port map( A1 => n6315, A2 => REGISTERS_29_11_port, B1 => 
                           n6587, B2 => REGISTERS_25_11_port, ZN => n6317);
   U1757 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_11_port, B1 => 
                           n6599, B2 => REGISTERS_17_11_port, ZN => n6316);
   U1758 : NAND4_X1 port map( A1 => n6319, A2 => n6318, A3 => n6317, A4 => 
                           n6316, ZN => n6326);
   U1759 : AOI22_X1 port map( A1 => n6459, A2 => REGISTERS_31_11_port, B1 => 
                           n6588, B2 => REGISTERS_28_11_port, ZN => n6324);
   U1760 : AOI22_X1 port map( A1 => n6590, A2 => REGISTERS_27_11_port, B1 => 
                           n6388, B2 => REGISTERS_30_11_port, ZN => n6323);
   U1761 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_11_port, B1 => 
                           n6593, B2 => REGISTERS_23_11_port, ZN => n6322);
   U1762 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_11_port, B1 => 
                           n6320, B2 => REGISTERS_16_11_port, ZN => n6321);
   U1763 : NAND4_X1 port map( A1 => n6324, A2 => n6323, A3 => n6322, A4 => 
                           n6321, ZN => n6325);
   U1764 : NOR2_X1 port map( A1 => n6326, A2 => n6325, ZN => n6340);
   U1765 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_11_port, B1 => 
                           n6623, B2 => REGISTERS_3_11_port, ZN => n6330);
   U1766 : AOI22_X1 port map( A1 => n6616, A2 => REGISTERS_7_11_port, B1 => 
                           n6614, B2 => REGISTERS_2_11_port, ZN => n6329);
   U1767 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_11_port, B1 => 
                           n6541, B2 => REGISTERS_1_11_port, ZN => n6328);
   U1768 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_11_port, B1 => 
                           n6624, B2 => REGISTERS_5_11_port, ZN => n6327);
   U1769 : NAND4_X1 port map( A1 => n6330, A2 => n6329, A3 => n6328, A4 => 
                           n6327, ZN => n6338);
   U1770 : AOI22_X1 port map( A1 => n6575, A2 => REGISTERS_11_11_port, B1 => 
                           n6331, B2 => REGISTERS_9_11_port, ZN => n6336);
   U1771 : AOI22_X1 port map( A1 => n6577, A2 => REGISTERS_13_11_port, B1 => 
                           n6616, B2 => REGISTERS_15_11_port, ZN => n6335);
   U1772 : AOI22_X1 port map( A1 => n6332, A2 => REGISTERS_14_11_port, B1 => 
                           n6570, B2 => REGISTERS_10_11_port, ZN => n6334);
   U1773 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_12_11_port, B1 => 
                           n6625, B2 => REGISTERS_8_11_port, ZN => n6333);
   U1774 : NAND4_X1 port map( A1 => n6336, A2 => n6335, A3 => n6334, A4 => 
                           n6333, ZN => n6337);
   U1775 : AOI22_X1 port map( A1 => n6482, A2 => n6338, B1 => n6480, B2 => 
                           n6337, ZN => n6339);
   U1776 : OAI21_X1 port map( B1 => n6641, B2 => n6340, A => n6339, ZN => N428)
                           ;
   U1777 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_10_port, B1 => 
                           n6603, B2 => REGISTERS_29_10_port, ZN => n6345);
   U1778 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_10_port, B1 => 
                           n6591, B2 => REGISTERS_16_10_port, ZN => n6344);
   U1779 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_10_port, B1 => 
                           n6599, B2 => REGISTERS_17_10_port, ZN => n6343);
   U1780 : AOI22_X1 port map( A1 => n6341, A2 => REGISTERS_20_10_port, B1 => 
                           n6555, B2 => REGISTERS_27_10_port, ZN => n6342);
   U1781 : NAND4_X1 port map( A1 => n6345, A2 => n6344, A3 => n6343, A4 => 
                           n6342, ZN => n6351);
   U1782 : AOI22_X1 port map( A1 => n6601, A2 => REGISTERS_18_10_port, B1 => 
                           n6587, B2 => REGISTERS_25_10_port, ZN => n6349);
   U1783 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_10_port, B1 => 
                           n6562, B2 => REGISTERS_19_10_port, ZN => n6348);
   U1784 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_10_port, B1 => 
                           n6588, B2 => REGISTERS_28_10_port, ZN => n6347);
   U1785 : AOI22_X1 port map( A1 => n6593, A2 => REGISTERS_23_10_port, B1 => 
                           n6388, B2 => REGISTERS_30_10_port, ZN => n6346);
   U1786 : NAND4_X1 port map( A1 => n6349, A2 => n6348, A3 => n6347, A4 => 
                           n6346, ZN => n6350);
   U1787 : NOR2_X1 port map( A1 => n6351, A2 => n6350, ZN => n6363);
   U1788 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_10_port, B1 => 
                           n6627, B2 => REGISTERS_1_10_port, ZN => n6355);
   U1789 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_7_10_port, B1 => 
                           n6628, B2 => REGISTERS_2_10_port, ZN => n6354);
   U1790 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_0_10_port, B1 => 
                           n6617, B2 => REGISTERS_3_10_port, ZN => n6353);
   U1791 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_10_port, B1 => 
                           n6577, B2 => REGISTERS_5_10_port, ZN => n6352);
   U1792 : NAND4_X1 port map( A1 => n6355, A2 => n6354, A3 => n6353, A4 => 
                           n6352, ZN => n6361);
   U1793 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_15_10_port, B1 => 
                           n6575, B2 => REGISTERS_11_10_port, ZN => n6359);
   U1794 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_10_port, B1 => 
                           n6624, B2 => REGISTERS_13_10_port, ZN => n6358);
   U1795 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_8_10_port, B1 => 
                           n6541, B2 => REGISTERS_9_10_port, ZN => n6357);
   U1796 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_10_port, B1 => 
                           n6614, B2 => REGISTERS_10_10_port, ZN => n6356);
   U1797 : NAND4_X1 port map( A1 => n6359, A2 => n6358, A3 => n6357, A4 => 
                           n6356, ZN => n6360);
   U1798 : AOI22_X1 port map( A1 => n6482, A2 => n6361, B1 => n6480, B2 => 
                           n6360, ZN => n6362);
   U1799 : OAI21_X1 port map( B1 => n6641, B2 => n6363, A => n6362, ZN => N427)
                           ;
   U1800 : AOI22_X1 port map( A1 => n6601, A2 => REGISTERS_18_9_port, B1 => 
                           n6594, B2 => REGISTERS_26_9_port, ZN => n6368);
   U1801 : AOI22_X1 port map( A1 => n6364, A2 => REGISTERS_23_9_port, B1 => 
                           n6388, B2 => REGISTERS_30_9_port, ZN => n6367);
   U1802 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_9_port, B1 => 
                           n6591, B2 => REGISTERS_16_9_port, ZN => n6366);
   U1803 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_9_port, B1 => 
                           n6603, B2 => REGISTERS_29_9_port, ZN => n6365);
   U1804 : NAND4_X1 port map( A1 => n6368, A2 => n6367, A3 => n6366, A4 => 
                           n6365, ZN => n6375);
   U1805 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_9_port, B1 => 
                           n6605, B2 => REGISTERS_24_9_port, ZN => n6373);
   U1806 : AOI22_X1 port map( A1 => n6416, A2 => REGISTERS_17_9_port, B1 => 
                           n6555, B2 => REGISTERS_27_9_port, ZN => n6372);
   U1807 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_9_port, B1 => 
                           n6604, B2 => REGISTERS_19_9_port, ZN => n6371);
   U1808 : AOI22_X1 port map( A1 => n6369, A2 => REGISTERS_21_9_port, B1 => 
                           n6587, B2 => REGISTERS_25_9_port, ZN => n6370);
   U1809 : NAND4_X1 port map( A1 => n6373, A2 => n6372, A3 => n6371, A4 => 
                           n6370, ZN => n6374);
   U1810 : NOR2_X1 port map( A1 => n6375, A2 => n6374, ZN => n6387);
   U1811 : AOI22_X1 port map( A1 => n6616, A2 => REGISTERS_7_9_port, B1 => 
                           n6627, B2 => REGISTERS_1_9_port, ZN => n6379);
   U1812 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_4_9_port, B1 => 
                           n6617, B2 => REGISTERS_3_9_port, ZN => n6378);
   U1813 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_9_port, B1 => 
                           n6628, B2 => REGISTERS_2_9_port, ZN => n6377);
   U1814 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_9_port, B1 => 
                           n6576, B2 => REGISTERS_0_9_port, ZN => n6376);
   U1815 : NAND4_X1 port map( A1 => n6379, A2 => n6378, A3 => n6377, A4 => 
                           n6376, ZN => n6385);
   U1816 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_9_port, B1 => 
                           n6577, B2 => REGISTERS_13_9_port, ZN => n6383);
   U1817 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_15_9_port, B1 => 
                           n6541, B2 => REGISTERS_9_9_port, ZN => n6382);
   U1818 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_9_port, B1 => 
                           n6628, B2 => REGISTERS_10_9_port, ZN => n6381);
   U1819 : AOI22_X1 port map( A1 => n6625, A2 => REGISTERS_8_9_port, B1 => 
                           n6623, B2 => REGISTERS_11_9_port, ZN => n6380);
   U1820 : NAND4_X1 port map( A1 => n6383, A2 => n6382, A3 => n6381, A4 => 
                           n6380, ZN => n6384);
   U1821 : AOI22_X1 port map( A1 => n6482, A2 => n6385, B1 => n6480, B2 => 
                           n6384, ZN => n6386);
   U1822 : OAI21_X1 port map( B1 => n6586, B2 => n6387, A => n6386, ZN => N426)
                           ;
   U1823 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_8_port, B1 => 
                           n6599, B2 => REGISTERS_17_8_port, ZN => n6392);
   U1824 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_8_port, B1 => 
                           n6593, B2 => REGISTERS_23_8_port, ZN => n6391);
   U1825 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_8_port, B1 => 
                           n6594, B2 => REGISTERS_26_8_port, ZN => n6390);
   U1826 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_8_port, B1 => 
                           n6388, B2 => REGISTERS_30_8_port, ZN => n6389);
   U1827 : NAND4_X1 port map( A1 => n6392, A2 => n6391, A3 => n6390, A4 => 
                           n6389, ZN => n6399);
   U1828 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_8_port, B1 => 
                           n6555, B2 => REGISTERS_27_8_port, ZN => n6397);
   U1829 : AOI22_X1 port map( A1 => n6393, A2 => REGISTERS_22_8_port, B1 => 
                           n6459, B2 => REGISTERS_31_8_port, ZN => n6396);
   U1830 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_8_port, B1 => 
                           n6587, B2 => REGISTERS_25_8_port, ZN => n6395);
   U1831 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_8_port, B1 => 
                           n6603, B2 => REGISTERS_29_8_port, ZN => n6394);
   U1832 : NAND4_X1 port map( A1 => n6397, A2 => n6396, A3 => n6395, A4 => 
                           n6394, ZN => n6398);
   U1833 : NOR2_X1 port map( A1 => n6399, A2 => n6398, ZN => n6411);
   U1834 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_4_8_port, B1 => 
                           n6624, B2 => REGISTERS_5_8_port, ZN => n6403);
   U1835 : AOI22_X1 port map( A1 => n6625, A2 => REGISTERS_0_8_port, B1 => 
                           n6570, B2 => REGISTERS_2_8_port, ZN => n6402);
   U1836 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_7_8_port, B1 => 
                           n6575, B2 => REGISTERS_3_8_port, ZN => n6401);
   U1837 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_8_port, B1 => 
                           n6627, B2 => REGISTERS_1_8_port, ZN => n6400);
   U1838 : NAND4_X1 port map( A1 => n6403, A2 => n6402, A3 => n6401, A4 => 
                           n6400, ZN => n6409);
   U1839 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_8_port, B1 => 
                           n6617, B2 => REGISTERS_11_8_port, ZN => n6407);
   U1840 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_8_port, B1 => 
                           n6614, B2 => REGISTERS_10_8_port, ZN => n6406);
   U1841 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_14_8_port, B1 => 
                           n6541, B2 => REGISTERS_9_8_port, ZN => n6405);
   U1842 : AOI22_X1 port map( A1 => n6569, A2 => REGISTERS_12_8_port, B1 => 
                           n6616, B2 => REGISTERS_15_8_port, ZN => n6404);
   U1843 : NAND4_X1 port map( A1 => n6407, A2 => n6406, A3 => n6405, A4 => 
                           n6404, ZN => n6408);
   U1844 : AOI22_X1 port map( A1 => n6482, A2 => n6409, B1 => n6480, B2 => 
                           n6408, ZN => n6410);
   U1845 : OAI21_X1 port map( B1 => n6641, B2 => n6411, A => n6410, ZN => N425)
                           ;
   U1846 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_7_port, B1 => 
                           n6587, B2 => REGISTERS_25_7_port, ZN => n6415);
   U1847 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_7_port, B1 => 
                           n6555, B2 => REGISTERS_27_7_port, ZN => n6414);
   U1848 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_7_port, B1 => 
                           n6589, B2 => REGISTERS_30_7_port, ZN => n6413);
   U1849 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_7_port, B1 => 
                           n6593, B2 => REGISTERS_23_7_port, ZN => n6412);
   U1850 : NAND4_X1 port map( A1 => n6415, A2 => n6414, A3 => n6413, A4 => 
                           n6412, ZN => n6422);
   U1851 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_7_port, B1 => 
                           n6601, B2 => REGISTERS_18_7_port, ZN => n6420);
   U1852 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_7_port, B1 => 
                           n6591, B2 => REGISTERS_16_7_port, ZN => n6419);
   U1853 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_7_port, B1 => 
                           n6604, B2 => REGISTERS_19_7_port, ZN => n6418);
   U1854 : AOI22_X1 port map( A1 => n6416, A2 => REGISTERS_17_7_port, B1 => 
                           n6603, B2 => REGISTERS_29_7_port, ZN => n6417);
   U1855 : NAND4_X1 port map( A1 => n6420, A2 => n6419, A3 => n6418, A4 => 
                           n6417, ZN => n6421);
   U1856 : NOR2_X1 port map( A1 => n6422, A2 => n6421, ZN => n6434);
   U1857 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_7_port, B1 => 
                           n6541, B2 => REGISTERS_1_7_port, ZN => n6426);
   U1858 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_7_port, B1 => 
                           n6624, B2 => REGISTERS_5_7_port, ZN => n6425);
   U1859 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_7_port, B1 => 
                           n6628, B2 => REGISTERS_2_7_port, ZN => n6424);
   U1860 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_7_port, B1 => 
                           n6474, B2 => REGISTERS_7_7_port, ZN => n6423);
   U1861 : NAND4_X1 port map( A1 => n6426, A2 => n6425, A3 => n6424, A4 => 
                           n6423, ZN => n6432);
   U1862 : AOI22_X1 port map( A1 => n6616, A2 => REGISTERS_15_7_port, B1 => 
                           n6575, B2 => REGISTERS_11_7_port, ZN => n6430);
   U1863 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_8_7_port, B1 => 
                           n6627, B2 => REGISTERS_9_7_port, ZN => n6429);
   U1864 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_13_7_port, B1 => 
                           n6570, B2 => REGISTERS_10_7_port, ZN => n6428);
   U1865 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_7_port, B1 => 
                           n6569, B2 => REGISTERS_12_7_port, ZN => n6427);
   U1866 : NAND4_X1 port map( A1 => n6430, A2 => n6429, A3 => n6428, A4 => 
                           n6427, ZN => n6431);
   U1867 : AOI22_X1 port map( A1 => n6482, A2 => n6432, B1 => n6480, B2 => 
                           n6431, ZN => n6433);
   U1868 : OAI21_X1 port map( B1 => n6586, B2 => n6434, A => n6433, ZN => N424)
                           ;
   U1869 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_6_port, B1 => 
                           n6591, B2 => REGISTERS_16_6_port, ZN => n6438);
   U1870 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_6_port, B1 => 
                           n6561, B2 => REGISTERS_28_6_port, ZN => n6437);
   U1871 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_6_port, B1 => 
                           n6603, B2 => REGISTERS_29_6_port, ZN => n6436);
   U1872 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_6_port, B1 => 
                           n6555, B2 => REGISTERS_27_6_port, ZN => n6435);
   U1873 : NAND4_X1 port map( A1 => n6438, A2 => n6437, A3 => n6436, A4 => 
                           n6435, ZN => n6445);
   U1874 : AOI22_X1 port map( A1 => n6439, A2 => REGISTERS_25_6_port, B1 => 
                           n6593, B2 => REGISTERS_23_6_port, ZN => n6443);
   U1875 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_6_port, B1 => 
                           n6599, B2 => REGISTERS_17_6_port, ZN => n6442);
   U1876 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_6_port, B1 => 
                           n6604, B2 => REGISTERS_19_6_port, ZN => n6441);
   U1877 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_6_port, B1 => 
                           n6589, B2 => REGISTERS_30_6_port, ZN => n6440);
   U1878 : NAND4_X1 port map( A1 => n6443, A2 => n6442, A3 => n6441, A4 => 
                           n6440, ZN => n6444);
   U1879 : NOR2_X1 port map( A1 => n6445, A2 => n6444, ZN => n6458);
   U1880 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_6_port, B1 => 
                           n6541, B2 => REGISTERS_1_6_port, ZN => n6449);
   U1881 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_6_port, B1 => 
                           n6623, B2 => REGISTERS_3_6_port, ZN => n6448);
   U1882 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_6_port, B1 => 
                           n6614, B2 => REGISTERS_2_6_port, ZN => n6447);
   U1883 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_6_port, B1 => 
                           n6576, B2 => REGISTERS_0_6_port, ZN => n6446);
   U1884 : NAND4_X1 port map( A1 => n6449, A2 => n6448, A3 => n6447, A4 => 
                           n6446, ZN => n6455);
   U1885 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_6_port, B1 => 
                           n6627, B2 => REGISTERS_9_6_port, ZN => n6453);
   U1886 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_6_port, B1 => 
                           n6629, B2 => REGISTERS_15_6_port, ZN => n6452);
   U1887 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_6_port, B1 => 
                           n6623, B2 => REGISTERS_11_6_port, ZN => n6451);
   U1888 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_13_6_port, B1 => 
                           n6615, B2 => REGISTERS_8_6_port, ZN => n6450);
   U1889 : NAND4_X1 port map( A1 => n6453, A2 => n6452, A3 => n6451, A4 => 
                           n6450, ZN => n6454);
   U1890 : AOI22_X1 port map( A1 => n6456, A2 => n6455, B1 => n6480, B2 => 
                           n6454, ZN => n6457);
   U1891 : OAI21_X1 port map( B1 => n6641, B2 => n6458, A => n6457, ZN => N423)
                           ;
   U1892 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_5_port, B1 => 
                           n6591, B2 => REGISTERS_16_5_port, ZN => n6463);
   U1893 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_5_port, B1 => 
                           n6459, B2 => REGISTERS_31_5_port, ZN => n6462);
   U1894 : AOI22_X1 port map( A1 => n6603, A2 => REGISTERS_29_5_port, B1 => 
                           n6589, B2 => REGISTERS_30_5_port, ZN => n6461);
   U1895 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_5_port, B1 => 
                           n6599, B2 => REGISTERS_17_5_port, ZN => n6460);
   U1896 : NAND4_X1 port map( A1 => n6463, A2 => n6462, A3 => n6461, A4 => 
                           n6460, ZN => n6469);
   U1897 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_5_port, B1 => 
                           n6604, B2 => REGISTERS_19_5_port, ZN => n6467);
   U1898 : AOI22_X1 port map( A1 => n6587, A2 => REGISTERS_25_5_port, B1 => 
                           n6593, B2 => REGISTERS_23_5_port, ZN => n6466);
   U1899 : AOI22_X1 port map( A1 => n6507, A2 => REGISTERS_26_5_port, B1 => 
                           n6561, B2 => REGISTERS_28_5_port, ZN => n6465);
   U1900 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_5_port, B1 => 
                           n6555, B2 => REGISTERS_27_5_port, ZN => n6464);
   U1901 : NAND4_X1 port map( A1 => n6467, A2 => n6466, A3 => n6465, A4 => 
                           n6464, ZN => n6468);
   U1902 : NOR2_X1 port map( A1 => n6469, A2 => n6468, ZN => n6484);
   U1903 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_5_port, B1 => 
                           n6474, B2 => REGISTERS_7_5_port, ZN => n6473);
   U1904 : AOI22_X1 port map( A1 => n6576, A2 => REGISTERS_0_5_port, B1 => 
                           n6541, B2 => REGISTERS_1_5_port, ZN => n6472);
   U1905 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_5_port, B1 => 
                           n6617, B2 => REGISTERS_3_5_port, ZN => n6471);
   U1906 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_5_port, B1 => 
                           n6614, B2 => REGISTERS_2_5_port, ZN => n6470);
   U1907 : NAND4_X1 port map( A1 => n6473, A2 => n6472, A3 => n6471, A4 => 
                           n6470, ZN => n6481);
   U1908 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_5_port, B1 => 
                           n6615, B2 => REGISTERS_8_5_port, ZN => n6478);
   U1909 : AOI22_X1 port map( A1 => n6474, A2 => REGISTERS_15_5_port, B1 => 
                           n6623, B2 => REGISTERS_11_5_port, ZN => n6477);
   U1910 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_5_port, B1 => 
                           n6627, B2 => REGISTERS_9_5_port, ZN => n6476);
   U1911 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_13_5_port, B1 => 
                           n6614, B2 => REGISTERS_10_5_port, ZN => n6475);
   U1912 : NAND4_X1 port map( A1 => n6478, A2 => n6477, A3 => n6476, A4 => 
                           n6475, ZN => n6479);
   U1913 : AOI22_X1 port map( A1 => n6482, A2 => n6481, B1 => n6480, B2 => 
                           n6479, ZN => n6483);
   U1914 : OAI21_X1 port map( B1 => n6586, B2 => n6484, A => n6483, ZN => N422)
                           ;
   U1915 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_4_port, B1 => 
                           n6593, B2 => REGISTERS_23_4_port, ZN => n6488);
   U1916 : AOI22_X1 port map( A1 => n6507, A2 => REGISTERS_26_4_port, B1 => 
                           n6587, B2 => REGISTERS_25_4_port, ZN => n6487);
   U1917 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_4_port, B1 => 
                           n6601, B2 => REGISTERS_18_4_port, ZN => n6486);
   U1918 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_4_port, B1 => 
                           n6603, B2 => REGISTERS_29_4_port, ZN => n6485);
   U1919 : NAND4_X1 port map( A1 => n6488, A2 => n6487, A3 => n6486, A4 => 
                           n6485, ZN => n6494);
   U1920 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_4_port, B1 => 
                           n6591, B2 => REGISTERS_16_4_port, ZN => n6492);
   U1921 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_4_port, B1 => 
                           n6555, B2 => REGISTERS_27_4_port, ZN => n6491);
   U1922 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_4_port, B1 => 
                           n6605, B2 => REGISTERS_24_4_port, ZN => n6490);
   U1923 : AOI22_X1 port map( A1 => n6599, A2 => REGISTERS_17_4_port, B1 => 
                           n6589, B2 => REGISTERS_30_4_port, ZN => n6489);
   U1924 : NAND4_X1 port map( A1 => n6492, A2 => n6491, A3 => n6490, A4 => 
                           n6489, ZN => n6493);
   U1925 : NOR2_X1 port map( A1 => n6494, A2 => n6493, ZN => n6506);
   U1926 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_4_port, B1 => 
                           n6541, B2 => REGISTERS_1_4_port, ZN => n6498);
   U1927 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_4_port, B1 => 
                           n6628, B2 => REGISTERS_2_4_port, ZN => n6497);
   U1928 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_4_port, B1 => 
                           n6623, B2 => REGISTERS_3_4_port, ZN => n6496);
   U1929 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_4_port, B1 => 
                           n6629, B2 => REGISTERS_7_4_port, ZN => n6495);
   U1930 : NAND4_X1 port map( A1 => n6498, A2 => n6497, A3 => n6496, A4 => 
                           n6495, ZN => n6504);
   U1931 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_13_4_port, B1 => 
                           n6614, B2 => REGISTERS_10_4_port, ZN => n6502);
   U1932 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_4_port, B1 => 
                           n6627, B2 => REGISTERS_9_4_port, ZN => n6501);
   U1933 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_4_port, B1 => 
                           n6575, B2 => REGISTERS_11_4_port, ZN => n6500);
   U1934 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_4_port, B1 => 
                           n6576, B2 => REGISTERS_8_4_port, ZN => n6499);
   U1935 : NAND4_X1 port map( A1 => n6502, A2 => n6501, A3 => n6500, A4 => 
                           n6499, ZN => n6503);
   U1936 : AOI22_X1 port map( A1 => n6638, A2 => n6504, B1 => n6636, B2 => 
                           n6503, ZN => n6505);
   U1937 : OAI21_X1 port map( B1 => n6641, B2 => n6506, A => n6505, ZN => N421)
                           ;
   U1938 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_3_port, B1 => 
                           n6599, B2 => REGISTERS_17_3_port, ZN => n6511);
   U1939 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_3_port, B1 => 
                           n6507, B2 => REGISTERS_26_3_port, ZN => n6510);
   U1940 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_3_port, B1 => 
                           n6593, B2 => REGISTERS_23_3_port, ZN => n6509);
   U1941 : AOI22_X1 port map( A1 => n6555, A2 => REGISTERS_27_3_port, B1 => 
                           n6589, B2 => REGISTERS_30_3_port, ZN => n6508);
   U1942 : NAND4_X1 port map( A1 => n6511, A2 => n6510, A3 => n6509, A4 => 
                           n6508, ZN => n6517);
   U1943 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_3_port, B1 => 
                           n6605, B2 => REGISTERS_24_3_port, ZN => n6515);
   U1944 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_3_port, B1 => 
                           n6603, B2 => REGISTERS_29_3_port, ZN => n6514);
   U1945 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_3_port, B1 => 
                           n6587, B2 => REGISTERS_25_3_port, ZN => n6513);
   U1946 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_3_port, B1 => 
                           n6591, B2 => REGISTERS_16_3_port, ZN => n6512);
   U1947 : NAND4_X1 port map( A1 => n6515, A2 => n6514, A3 => n6513, A4 => 
                           n6512, ZN => n6516);
   U1948 : NOR2_X1 port map( A1 => n6517, A2 => n6516, ZN => n6529);
   U1949 : AOI22_X1 port map( A1 => n6616, A2 => REGISTERS_7_3_port, B1 => 
                           n6570, B2 => REGISTERS_2_3_port, ZN => n6521);
   U1950 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_3_port, B1 => 
                           n6541, B2 => REGISTERS_1_3_port, ZN => n6520);
   U1951 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_3_port, B1 => 
                           n6625, B2 => REGISTERS_0_3_port, ZN => n6519);
   U1952 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_3_port, B1 => 
                           n6623, B2 => REGISTERS_3_3_port, ZN => n6518);
   U1953 : NAND4_X1 port map( A1 => n6521, A2 => n6520, A3 => n6519, A4 => 
                           n6518, ZN => n6527);
   U1954 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_13_3_port, B1 => 
                           n6628, B2 => REGISTERS_10_3_port, ZN => n6525);
   U1955 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_3_port, B1 => 
                           n6623, B2 => REGISTERS_11_3_port, ZN => n6524);
   U1956 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_3_port, B1 => 
                           n6627, B2 => REGISTERS_9_3_port, ZN => n6523);
   U1957 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_3_port, B1 => 
                           n6569, B2 => REGISTERS_12_3_port, ZN => n6522);
   U1958 : NAND4_X1 port map( A1 => n6525, A2 => n6524, A3 => n6523, A4 => 
                           n6522, ZN => n6526);
   U1959 : AOI22_X1 port map( A1 => n6638, A2 => n6527, B1 => n6636, B2 => 
                           n6526, ZN => n6528);
   U1960 : OAI21_X1 port map( B1 => n6586, B2 => n6529, A => n6528, ZN => N420)
                           ;
   U1961 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_2_port, B1 => 
                           n6593, B2 => REGISTERS_23_2_port, ZN => n6533);
   U1962 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_2_port, B1 => 
                           n6591, B2 => REGISTERS_16_2_port, ZN => n6532);
   U1963 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_2_port, B1 => 
                           n6587, B2 => REGISTERS_25_2_port, ZN => n6531);
   U1964 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_2_port, B1 => 
                           n6589, B2 => REGISTERS_30_2_port, ZN => n6530);
   U1965 : NAND4_X1 port map( A1 => n6533, A2 => n6532, A3 => n6531, A4 => 
                           n6530, ZN => n6540);
   U1966 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_2_port, B1 => 
                           n6599, B2 => REGISTERS_17_2_port, ZN => n6538);
   U1967 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_2_port, B1 => 
                           n6555, B2 => REGISTERS_27_2_port, ZN => n6537);
   U1968 : AOI22_X1 port map( A1 => n6534, A2 => REGISTERS_24_2_port, B1 => 
                           n6601, B2 => REGISTERS_18_2_port, ZN => n6536);
   U1969 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_2_port, B1 => 
                           n6603, B2 => REGISTERS_29_2_port, ZN => n6535);
   U1970 : NAND4_X1 port map( A1 => n6538, A2 => n6537, A3 => n6536, A4 => 
                           n6535, ZN => n6539);
   U1971 : NOR2_X1 port map( A1 => n6540, A2 => n6539, ZN => n6554);
   U1972 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_2_port, B1 => 
                           n6577, B2 => REGISTERS_5_2_port, ZN => n6546);
   U1973 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_2_port, B1 => 
                           n6570, B2 => REGISTERS_2_2_port, ZN => n6545);
   U1974 : AOI22_X1 port map( A1 => n6617, A2 => REGISTERS_3_2_port, B1 => 
                           n6541, B2 => REGISTERS_1_2_port, ZN => n6544);
   U1975 : AOI22_X1 port map( A1 => n6542, A2 => REGISTERS_6_2_port, B1 => 
                           n6629, B2 => REGISTERS_7_2_port, ZN => n6543);
   U1976 : NAND4_X1 port map( A1 => n6546, A2 => n6545, A3 => n6544, A4 => 
                           n6543, ZN => n6552);
   U1977 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_2_port, B1 => 
                           n6616, B2 => REGISTERS_15_2_port, ZN => n6550);
   U1978 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_2_port, B1 => 
                           n6577, B2 => REGISTERS_13_2_port, ZN => n6549);
   U1979 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_8_2_port, B1 => 
                           n6627, B2 => REGISTERS_9_2_port, ZN => n6548);
   U1980 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_2_port, B1 => 
                           n6575, B2 => REGISTERS_11_2_port, ZN => n6547);
   U1981 : NAND4_X1 port map( A1 => n6550, A2 => n6549, A3 => n6548, A4 => 
                           n6547, ZN => n6551);
   U1982 : AOI22_X1 port map( A1 => n6638, A2 => n6552, B1 => n6636, B2 => 
                           n6551, ZN => n6553);
   U1983 : OAI21_X1 port map( B1 => n6641, B2 => n6554, A => n6553, ZN => N419)
                           ;
   U1984 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_1_port, B1 => 
                           n6587, B2 => REGISTERS_25_1_port, ZN => n6559);
   U1985 : AOI22_X1 port map( A1 => n6591, A2 => REGISTERS_16_1_port, B1 => 
                           n6603, B2 => REGISTERS_29_1_port, ZN => n6558);
   U1986 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_1_port, B1 => 
                           n6555, B2 => REGISTERS_27_1_port, ZN => n6557);
   U1987 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_1_port, B1 => 
                           n6593, B2 => REGISTERS_23_1_port, ZN => n6556);
   U1988 : NAND4_X1 port map( A1 => n6559, A2 => n6558, A3 => n6557, A4 => 
                           n6556, ZN => n6568);
   U1989 : AOI22_X1 port map( A1 => n6560, A2 => REGISTERS_18_1_port, B1 => 
                           n6589, B2 => REGISTERS_30_1_port, ZN => n6566);
   U1990 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_1_port, B1 => 
                           n6561, B2 => REGISTERS_28_1_port, ZN => n6565);
   U1991 : AOI22_X1 port map( A1 => n6562, A2 => REGISTERS_19_1_port, B1 => 
                           n6599, B2 => REGISTERS_17_1_port, ZN => n6564);
   U1992 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_1_port, B1 => 
                           n6605, B2 => REGISTERS_24_1_port, ZN => n6563);
   U1993 : NAND4_X1 port map( A1 => n6566, A2 => n6565, A3 => n6564, A4 => 
                           n6563, ZN => n6567);
   U1994 : NOR2_X1 port map( A1 => n6568, A2 => n6567, ZN => n6585);
   U1995 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_1_port, B1 => 
                           n6569, B2 => REGISTERS_4_1_port, ZN => n6574);
   U1996 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_7_1_port, B1 => 
                           n6627, B2 => REGISTERS_1_1_port, ZN => n6573);
   U1997 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_1_port, B1 => 
                           n6617, B2 => REGISTERS_3_1_port, ZN => n6572);
   U1998 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_1_port, B1 => 
                           n6570, B2 => REGISTERS_2_1_port, ZN => n6571);
   U1999 : NAND4_X1 port map( A1 => n6574, A2 => n6573, A3 => n6572, A4 => 
                           n6571, ZN => n6583);
   U2000 : AOI22_X1 port map( A1 => n6629, A2 => REGISTERS_15_1_port, B1 => 
                           n6575, B2 => REGISTERS_11_1_port, ZN => n6581);
   U2001 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_12_1_port, B1 => 
                           n6576, B2 => REGISTERS_8_1_port, ZN => n6580);
   U2002 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_1_port, B1 => 
                           n6577, B2 => REGISTERS_13_1_port, ZN => n6579);
   U2003 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_1_port, B1 => 
                           n6627, B2 => REGISTERS_9_1_port, ZN => n6578);
   U2004 : NAND4_X1 port map( A1 => n6581, A2 => n6580, A3 => n6579, A4 => 
                           n6578, ZN => n6582);
   U2005 : AOI22_X1 port map( A1 => n6638, A2 => n6583, B1 => n6636, B2 => 
                           n6582, ZN => n6584);
   U2006 : OAI21_X1 port map( B1 => n6586, B2 => n6585, A => n6584, ZN => N418)
                           ;
   U2007 : AOI22_X1 port map( A1 => n6588, A2 => REGISTERS_28_0_port, B1 => 
                           n6587, B2 => REGISTERS_25_0_port, ZN => n6598);
   U2008 : AOI22_X1 port map( A1 => n6590, A2 => REGISTERS_27_0_port, B1 => 
                           n6589, B2 => REGISTERS_30_0_port, ZN => n6597);
   U2009 : AOI22_X1 port map( A1 => n6592, A2 => REGISTERS_22_0_port, B1 => 
                           n6591, B2 => REGISTERS_16_0_port, ZN => n6596);
   U2010 : AOI22_X1 port map( A1 => n6594, A2 => REGISTERS_26_0_port, B1 => 
                           n6593, B2 => REGISTERS_23_0_port, ZN => n6595);
   U2011 : NAND4_X1 port map( A1 => n6598, A2 => n6597, A3 => n6596, A4 => 
                           n6595, ZN => n6612);
   U2012 : AOI22_X1 port map( A1 => n6600, A2 => REGISTERS_31_0_port, B1 => 
                           n6599, B2 => REGISTERS_17_0_port, ZN => n6610);
   U2013 : AOI22_X1 port map( A1 => n6602, A2 => REGISTERS_20_0_port, B1 => 
                           n6601, B2 => REGISTERS_18_0_port, ZN => n6609);
   U2014 : AOI22_X1 port map( A1 => n6604, A2 => REGISTERS_19_0_port, B1 => 
                           n6603, B2 => REGISTERS_29_0_port, ZN => n6608);
   U2015 : AOI22_X1 port map( A1 => n6606, A2 => REGISTERS_21_0_port, B1 => 
                           n6605, B2 => REGISTERS_24_0_port, ZN => n6607);
   U2016 : NAND4_X1 port map( A1 => n6610, A2 => n6609, A3 => n6608, A4 => 
                           n6607, ZN => n6611);
   U2017 : NOR2_X1 port map( A1 => n6612, A2 => n6611, ZN => n6640);
   U2018 : AOI22_X1 port map( A1 => n6613, A2 => REGISTERS_5_0_port, B1 => 
                           n6627, B2 => REGISTERS_1_0_port, ZN => n6622);
   U2019 : AOI22_X1 port map( A1 => n6615, A2 => REGISTERS_0_0_port, B1 => 
                           n6614, B2 => REGISTERS_2_0_port, ZN => n6621);
   U2020 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_6_0_port, B1 => 
                           n6616, B2 => REGISTERS_7_0_port, ZN => n6620);
   U2021 : AOI22_X1 port map( A1 => n6618, A2 => REGISTERS_4_0_port, B1 => 
                           n6617, B2 => REGISTERS_3_0_port, ZN => n6619);
   U2022 : NAND4_X1 port map( A1 => n6622, A2 => n6621, A3 => n6620, A4 => 
                           n6619, ZN => n6637);
   U2023 : AOI22_X1 port map( A1 => n6624, A2 => REGISTERS_13_0_port, B1 => 
                           n6623, B2 => REGISTERS_11_0_port, ZN => n6634);
   U2024 : AOI22_X1 port map( A1 => n6626, A2 => REGISTERS_12_0_port, B1 => 
                           n6625, B2 => REGISTERS_8_0_port, ZN => n6633);
   U2025 : AOI22_X1 port map( A1 => n6628, A2 => REGISTERS_10_0_port, B1 => 
                           n6627, B2 => REGISTERS_9_0_port, ZN => n6632);
   U2026 : AOI22_X1 port map( A1 => n6630, A2 => REGISTERS_14_0_port, B1 => 
                           n6629, B2 => REGISTERS_15_0_port, ZN => n6631);
   U2027 : NAND4_X1 port map( A1 => n6634, A2 => n6633, A3 => n6632, A4 => 
                           n6631, ZN => n6635);
   U2028 : AOI22_X1 port map( A1 => n6638, A2 => n6637, B1 => n6636, B2 => 
                           n6635, ZN => n6639);
   U2029 : OAI21_X1 port map( B1 => n6641, B2 => n6640, A => n6639, ZN => N417)
                           ;
   U2030 : NAND3_X1 port map( A1 => n5675, A2 => ENABLE, A3 => RD1, ZN => n7423
                           );
   U2031 : INV_X1 port map( A => ADD_RD1(3), ZN => n6670);
   U2032 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n6670, ZN => n6651);
   U2033 : INV_X1 port map( A => ADD_RD1(2), ZN => n6648);
   U2034 : INV_X1 port map( A => ADD_RD1(0), ZN => n6649);
   U2035 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => n6648, A3 => n6649, ZN =>
                           n6658);
   U2036 : NOR2_X1 port map( A1 => n6651, A2 => n6658, ZN => n7188);
   U2037 : CLKBUF_X1 port map( A => n7188, Z => n7381);
   U2038 : INV_X1 port map( A => ADD_RD1(1), ZN => n6642);
   U2039 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => n6642, A3 => n6649, ZN =>
                           n6663);
   U2040 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n6650);
   U2041 : NOR2_X1 port map( A1 => n6663, A2 => n6650, ZN => n7009);
   U2042 : CLKBUF_X1 port map( A => n7009, Z => n7368);
   U2043 : AOI22_X1 port map( A1 => REGISTERS_18_31_port, A2 => n7381, B1 => 
                           REGISTERS_28_31_port, B2 => n7368, ZN => n6647);
   U2044 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => n6642, 
                           ZN => n6659);
   U2045 : NOR2_X1 port map( A1 => n6650, A2 => n6659, ZN => n7380);
   U2046 : CLKBUF_X1 port map( A => n7380, Z => n7315);
   U2047 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n6643);
   U2048 : NAND2_X1 port map( A1 => n6643, A2 => ADD_RD1(0), ZN => n6662);
   U2049 : NOR2_X1 port map( A1 => n6662, A2 => n6650, ZN => n7216);
   U2050 : CLKBUF_X1 port map( A => n7216, Z => n7374);
   U2051 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n7315, B1 => 
                           REGISTERS_25_31_port, B2 => n7374, ZN => n6646);
   U2052 : NOR2_X1 port map( A1 => n6650, A2 => n6658, ZN => n7372);
   U2053 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n6664);
   U2054 : NOR2_X1 port map( A1 => n6651, A2 => n6664, ZN => n7215);
   U2055 : CLKBUF_X1 port map( A => n7215, Z => n7384);
   U2056 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n7372, B1 => 
                           REGISTERS_23_31_port, B2 => n7384, ZN => n6645);
   U2057 : NOR2_X1 port map( A1 => n6651, A2 => n6659, ZN => n7165);
   U2058 : CLKBUF_X1 port map( A => n7165, Z => n7370);
   U2059 : NAND2_X1 port map( A1 => n6643, A2 => n6649, ZN => n6661);
   U2060 : NOR2_X1 port map( A1 => n6661, A2 => n6650, ZN => n7387);
   U2061 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n7370, B1 => 
                           REGISTERS_24_31_port, B2 => n7387, ZN => n6644);
   U2062 : NAND4_X1 port map( A1 => n6647, A2 => n6646, A3 => n6645, A4 => 
                           n6644, ZN => n6657);
   U2063 : NOR2_X1 port map( A1 => n6651, A2 => n6661, ZN => n7386);
   U2064 : CLKBUF_X1 port map( A => n7386, Z => n7285);
   U2065 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => n6648, 
                           ZN => n6660);
   U2066 : NOR2_X1 port map( A1 => n6650, A2 => n6660, ZN => n7142);
   U2067 : CLKBUF_X1 port map( A => n7142, Z => n7369);
   U2068 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n7285, B1 => 
                           REGISTERS_27_31_port, B2 => n7369, ZN => n6655);
   U2069 : NOR2_X1 port map( A1 => n6651, A2 => n6663, ZN => n7314);
   U2070 : CLKBUF_X1 port map( A => n7314, Z => n7371);
   U2071 : NOR2_X1 port map( A1 => n6662, A2 => n6651, ZN => n7383);
   U2072 : CLKBUF_X1 port map( A => n7383, Z => n7335);
   U2073 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n7371, B1 => 
                           REGISTERS_17_31_port, B2 => n7335, ZN => n6654);
   U2074 : NOR2_X1 port map( A1 => n6650, A2 => n6664, ZN => n7338);
   U2075 : CLKBUF_X1 port map( A => n7338, Z => n7373);
   U2076 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), A3 => n6649, 
                           ZN => n6665);
   U2077 : NOR2_X1 port map( A1 => n6650, A2 => n6665, ZN => n7309);
   U2078 : AOI22_X1 port map( A1 => REGISTERS_31_31_port, A2 => n7373, B1 => 
                           REGISTERS_30_31_port, B2 => n7309, ZN => n6653);
   U2079 : NOR2_X1 port map( A1 => n6651, A2 => n6665, ZN => n7266);
   U2080 : CLKBUF_X1 port map( A => n7266, Z => n7382);
   U2081 : NOR2_X1 port map( A1 => n6651, A2 => n6660, ZN => n7336);
   U2082 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n7382, B1 => 
                           REGISTERS_19_31_port, B2 => n7336, ZN => n6652);
   U2083 : NAND4_X1 port map( A1 => n6655, A2 => n6654, A3 => n6653, A4 => 
                           n6652, ZN => n6656);
   U2084 : NOR2_X1 port map( A1 => n6657, A2 => n6656, ZN => n6678);
   U2085 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n7367, 
                           ZN => n7420);
   U2086 : CLKBUF_X1 port map( A => n7420, Z => n7234);
   U2087 : INV_X1 port map( A => n6658, ZN => n7405);
   U2088 : CLKBUF_X1 port map( A => n7405, Z => n7398);
   U2089 : INV_X1 port map( A => n6659, ZN => n7227);
   U2090 : AOI22_X1 port map( A1 => REGISTERS_2_31_port, A2 => n7398, B1 => 
                           REGISTERS_5_31_port, B2 => n7227, ZN => n6669);
   U2091 : INV_X1 port map( A => n6660, ZN => n7350);
   U2092 : CLKBUF_X1 port map( A => n7350, Z => n7357);
   U2093 : INV_X1 port map( A => n6661, ZN => n7406);
   U2094 : CLKBUF_X1 port map( A => n7406, Z => n7351);
   U2095 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n7357, B1 => 
                           REGISTERS_0_31_port, B2 => n7351, ZN => n6668);
   U2096 : INV_X1 port map( A => n6662, ZN => n7356);
   U2097 : CLKBUF_X1 port map( A => n7356, Z => n7395);
   U2098 : INV_X1 port map( A => n6663, ZN => n7251);
   U2099 : CLKBUF_X1 port map( A => n7251, Z => n7410);
   U2100 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n7395, B1 => 
                           REGISTERS_4_31_port, B2 => n7410, ZN => n6667);
   U2101 : INV_X1 port map( A => n6664, ZN => n7296);
   U2102 : INV_X1 port map( A => n6665, ZN => n7399);
   U2103 : CLKBUF_X1 port map( A => n7399, Z => n7411);
   U2104 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n7296, B1 => 
                           REGISTERS_6_31_port, B2 => n7411, ZN => n6666);
   U2105 : NAND4_X1 port map( A1 => n6669, A2 => n6668, A3 => n6667, A4 => 
                           n6666, ZN => n6676);
   U2106 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n6670, A3 => n7367, ZN => 
                           n7418);
   U2107 : CLKBUF_X1 port map( A => n7418, Z => n7257);
   U2108 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n7357, B1 => 
                           REGISTERS_8_31_port, B2 => n7351, ZN => n6674);
   U2109 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n7296, B1 => 
                           REGISTERS_13_31_port, B2 => n7227, ZN => n6673);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n7395, B1 => 
                           REGISTERS_12_31_port, B2 => n7251, ZN => n6672);
   U2111 : CLKBUF_X1 port map( A => n7399, Z => n7322);
   U2112 : AOI22_X1 port map( A1 => REGISTERS_10_31_port, A2 => n7398, B1 => 
                           REGISTERS_14_31_port, B2 => n7322, ZN => n6671);
   U2113 : NAND4_X1 port map( A1 => n6674, A2 => n6673, A3 => n6672, A4 => 
                           n6671, ZN => n6675);
   U2114 : AOI22_X1 port map( A1 => n7234, A2 => n6676, B1 => n7257, B2 => 
                           n6675, ZN => n6677);
   U2115 : OAI21_X1 port map( B1 => n7367, B2 => n6678, A => n6677, ZN => N416)
                           ;
   U2116 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n7315, B1 => 
                           REGISTERS_25_30_port, B2 => n7216, ZN => n6682);
   U2117 : CLKBUF_X1 port map( A => n7387, Z => n7337);
   U2118 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n7337, B1 => 
                           REGISTERS_20_30_port, B2 => n7314, ZN => n6681);
   U2119 : AOI22_X1 port map( A1 => REGISTERS_22_30_port, A2 => n7382, B1 => 
                           REGISTERS_27_30_port, B2 => n7369, ZN => n6680);
   U2120 : AOI22_X1 port map( A1 => REGISTERS_18_30_port, A2 => n7381, B1 => 
                           REGISTERS_16_30_port, B2 => n7386, ZN => n6679);
   U2121 : NAND4_X1 port map( A1 => n6682, A2 => n6681, A3 => n6680, A4 => 
                           n6679, ZN => n6688);
   U2122 : CLKBUF_X1 port map( A => n7372, Z => n7343);
   U2123 : AOI22_X1 port map( A1 => REGISTERS_26_30_port, A2 => n7343, B1 => 
                           REGISTERS_30_30_port, B2 => n7309, ZN => n6686);
   U2124 : AOI22_X1 port map( A1 => REGISTERS_31_30_port, A2 => n7338, B1 => 
                           REGISTERS_28_30_port, B2 => n7009, ZN => n6685);
   U2125 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n7384, B1 => 
                           REGISTERS_19_30_port, B2 => n7336, ZN => n6684);
   U2126 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n7335, B1 => 
                           REGISTERS_21_30_port, B2 => n7370, ZN => n6683);
   U2127 : NAND4_X1 port map( A1 => n6686, A2 => n6685, A3 => n6684, A4 => 
                           n6683, ZN => n6687);
   U2128 : NOR2_X1 port map( A1 => n6688, A2 => n6687, ZN => n6700);
   U2129 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n7395, B1 => 
                           REGISTERS_6_30_port, B2 => n7322, ZN => n6692);
   U2130 : CLKBUF_X1 port map( A => n7227, Z => n7412);
   U2131 : CLKBUF_X1 port map( A => n7251, Z => n7396);
   U2132 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n7412, B1 => 
                           REGISTERS_4_30_port, B2 => n7396, ZN => n6691);
   U2133 : CLKBUF_X1 port map( A => n7296, Z => n7400);
   U2134 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n7400, B1 => 
                           REGISTERS_0_30_port, B2 => n7351, ZN => n6690);
   U2135 : CLKBUF_X1 port map( A => n7350, Z => n7408);
   U2136 : AOI22_X1 port map( A1 => REGISTERS_2_30_port, A2 => n7398, B1 => 
                           REGISTERS_3_30_port, B2 => n7408, ZN => n6689);
   U2137 : NAND4_X1 port map( A1 => n6692, A2 => n6691, A3 => n6690, A4 => 
                           n6689, ZN => n6698);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n7296, B1 => 
                           REGISTERS_11_30_port, B2 => n7408, ZN => n6696);
   U2139 : CLKBUF_X1 port map( A => n7406, Z => n7397);
   U2140 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n7397, B1 => 
                           REGISTERS_9_30_port, B2 => n7356, ZN => n6695);
   U2141 : CLKBUF_X1 port map( A => n7227, Z => n7394);
   U2142 : AOI22_X1 port map( A1 => REGISTERS_10_30_port, A2 => n7398, B1 => 
                           REGISTERS_13_30_port, B2 => n7394, ZN => n6694);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_14_30_port, A2 => n7411, B1 => 
                           REGISTERS_12_30_port, B2 => n7396, ZN => n6693);
   U2144 : NAND4_X1 port map( A1 => n6696, A2 => n6695, A3 => n6694, A4 => 
                           n6693, ZN => n6697);
   U2145 : AOI22_X1 port map( A1 => n7234, A2 => n6698, B1 => n7257, B2 => 
                           n6697, ZN => n6699);
   U2146 : OAI21_X1 port map( B1 => n7367, B2 => n6700, A => n6699, ZN => N415)
                           ;
   U2147 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n7285, B1 => 
                           REGISTERS_25_29_port, B2 => n7216, ZN => n6704);
   U2148 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n7368, B1 => 
                           REGISTERS_30_29_port, B2 => n7309, ZN => n6703);
   U2149 : AOI22_X1 port map( A1 => REGISTERS_18_29_port, A2 => n7381, B1 => 
                           REGISTERS_29_29_port, B2 => n7380, ZN => n6702);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_22_29_port, A2 => n7382, B1 => 
                           REGISTERS_26_29_port, B2 => n7372, ZN => n6701);
   U2151 : NAND4_X1 port map( A1 => n6704, A2 => n6703, A3 => n6702, A4 => 
                           n6701, ZN => n6710);
   U2152 : AOI22_X1 port map( A1 => REGISTERS_31_29_port, A2 => n7373, B1 => 
                           REGISTERS_20_29_port, B2 => n7314, ZN => n6708);
   U2153 : CLKBUF_X1 port map( A => n7336, Z => n7375);
   U2154 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n7375, B1 => 
                           REGISTERS_27_29_port, B2 => n7142, ZN => n6707);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n7335, B1 => 
                           REGISTERS_24_29_port, B2 => n7387, ZN => n6706);
   U2156 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n7384, B1 => 
                           REGISTERS_21_29_port, B2 => n7165, ZN => n6705);
   U2157 : NAND4_X1 port map( A1 => n6708, A2 => n6707, A3 => n6706, A4 => 
                           n6705, ZN => n6709);
   U2158 : NOR2_X1 port map( A1 => n6710, A2 => n6709, ZN => n6722);
   U2159 : CLKBUF_X1 port map( A => n7356, Z => n7409);
   U2160 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n7357, B1 => 
                           REGISTERS_1_29_port, B2 => n7409, ZN => n6714);
   U2161 : CLKBUF_X1 port map( A => n7296, Z => n7407);
   U2162 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n7412, B1 => 
                           REGISTERS_7_29_port, B2 => n7407, ZN => n6713);
   U2163 : AOI22_X1 port map( A1 => REGISTERS_2_29_port, A2 => n7398, B1 => 
                           REGISTERS_6_29_port, B2 => n7322, ZN => n6712);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n7410, B1 => 
                           REGISTERS_0_29_port, B2 => n7351, ZN => n6711);
   U2165 : NAND4_X1 port map( A1 => n6714, A2 => n6713, A3 => n6712, A4 => 
                           n6711, ZN => n6720);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n7412, B1 => 
                           REGISTERS_14_29_port, B2 => n7322, ZN => n6718);
   U2167 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n7400, B1 => 
                           REGISTERS_9_29_port, B2 => n7409, ZN => n6717);
   U2168 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n7410, B1 => 
                           REGISTERS_11_29_port, B2 => n7408, ZN => n6716);
   U2169 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n7351, B1 => 
                           REGISTERS_10_29_port, B2 => n7405, ZN => n6715);
   U2170 : NAND4_X1 port map( A1 => n6718, A2 => n6717, A3 => n6716, A4 => 
                           n6715, ZN => n6719);
   U2171 : AOI22_X1 port map( A1 => n7234, A2 => n6720, B1 => n7257, B2 => 
                           n6719, ZN => n6721);
   U2172 : OAI21_X1 port map( B1 => n7367, B2 => n6722, A => n6721, ZN => N414)
                           ;
   U2173 : AOI22_X1 port map( A1 => REGISTERS_18_28_port, A2 => n7381, B1 => 
                           REGISTERS_20_28_port, B2 => n7314, ZN => n6726);
   U2174 : AOI22_X1 port map( A1 => REGISTERS_19_28_port, A2 => n7375, B1 => 
                           REGISTERS_17_28_port, B2 => n7383, ZN => n6725);
   U2175 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n7285, B1 => 
                           REGISTERS_28_28_port, B2 => n7009, ZN => n6724);
   U2176 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n7374, B1 => 
                           REGISTERS_31_28_port, B2 => n7338, ZN => n6723);
   U2177 : NAND4_X1 port map( A1 => n6726, A2 => n6725, A3 => n6724, A4 => 
                           n6723, ZN => n6732);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n7337, B1 => 
                           REGISTERS_29_28_port, B2 => n7380, ZN => n6730);
   U2179 : CLKBUF_X1 port map( A => n7309, Z => n7385);
   U2180 : AOI22_X1 port map( A1 => REGISTERS_30_28_port, A2 => n7385, B1 => 
                           REGISTERS_26_28_port, B2 => n7372, ZN => n6729);
   U2181 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n7369, B1 => 
                           REGISTERS_23_28_port, B2 => n7215, ZN => n6728);
   U2182 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n7370, B1 => 
                           REGISTERS_22_28_port, B2 => n7382, ZN => n6727);
   U2183 : NAND4_X1 port map( A1 => n6730, A2 => n6729, A3 => n6728, A4 => 
                           n6727, ZN => n6731);
   U2184 : NOR2_X1 port map( A1 => n6732, A2 => n6731, ZN => n6744);
   U2185 : AOI22_X1 port map( A1 => REGISTERS_2_28_port, A2 => n7398, B1 => 
                           REGISTERS_4_28_port, B2 => n7396, ZN => n6736);
   U2186 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n7412, B1 => 
                           REGISTERS_3_28_port, B2 => n7408, ZN => n6735);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_6_28_port, A2 => n7411, B1 => 
                           REGISTERS_1_28_port, B2 => n7409, ZN => n6734);
   U2188 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n7406, B1 => 
                           REGISTERS_7_28_port, B2 => n7407, ZN => n6733);
   U2189 : NAND4_X1 port map( A1 => n6736, A2 => n6735, A3 => n6734, A4 => 
                           n6733, ZN => n6742);
   U2190 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n7395, B1 => 
                           REGISTERS_13_28_port, B2 => n7394, ZN => n6740);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_10_28_port, A2 => n7398, B1 => 
                           REGISTERS_11_28_port, B2 => n7408, ZN => n6739);
   U2192 : AOI22_X1 port map( A1 => REGISTERS_14_28_port, A2 => n7411, B1 => 
                           REGISTERS_8_28_port, B2 => n7406, ZN => n6738);
   U2193 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n7410, B1 => 
                           REGISTERS_15_28_port, B2 => n7296, ZN => n6737);
   U2194 : NAND4_X1 port map( A1 => n6740, A2 => n6739, A3 => n6738, A4 => 
                           n6737, ZN => n6741);
   U2195 : AOI22_X1 port map( A1 => n7234, A2 => n6742, B1 => n7257, B2 => 
                           n6741, ZN => n6743);
   U2196 : OAI21_X1 port map( B1 => n7367, B2 => n6744, A => n6743, ZN => N413)
                           ;
   U2197 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n7337, B1 => 
                           REGISTERS_25_27_port, B2 => n7216, ZN => n6748);
   U2198 : AOI22_X1 port map( A1 => REGISTERS_19_27_port, A2 => n7336, B1 => 
                           REGISTERS_17_27_port, B2 => n7383, ZN => n6747);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n7338, B1 => 
                           REGISTERS_27_27_port, B2 => n7142, ZN => n6746);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n7315, B1 => 
                           REGISTERS_18_27_port, B2 => n7381, ZN => n6745);
   U2201 : NAND4_X1 port map( A1 => n6748, A2 => n6747, A3 => n6746, A4 => 
                           n6745, ZN => n6754);
   U2202 : AOI22_X1 port map( A1 => REGISTERS_30_27_port, A2 => n7385, B1 => 
                           REGISTERS_23_27_port, B2 => n7215, ZN => n6752);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n7371, B1 => 
                           REGISTERS_21_27_port, B2 => n7165, ZN => n6751);
   U2204 : AOI22_X1 port map( A1 => REGISTERS_26_27_port, A2 => n7343, B1 => 
                           REGISTERS_16_27_port, B2 => n7386, ZN => n6750);
   U2205 : AOI22_X1 port map( A1 => REGISTERS_22_27_port, A2 => n7382, B1 => 
                           REGISTERS_28_27_port, B2 => n7009, ZN => n6749);
   U2206 : NAND4_X1 port map( A1 => n6752, A2 => n6751, A3 => n6750, A4 => 
                           n6749, ZN => n6753);
   U2207 : NOR2_X1 port map( A1 => n6754, A2 => n6753, ZN => n6766);
   U2208 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n7395, B1 => 
                           REGISTERS_3_27_port, B2 => n7408, ZN => n6758);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n7410, B1 => 
                           REGISTERS_6_27_port, B2 => n7322, ZN => n6757);
   U2210 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n7400, B1 => 
                           REGISTERS_5_27_port, B2 => n7394, ZN => n6756);
   U2211 : CLKBUF_X1 port map( A => n7405, Z => n7358);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n7406, B1 => 
                           REGISTERS_2_27_port, B2 => n7358, ZN => n6755);
   U2213 : NAND4_X1 port map( A1 => n6758, A2 => n6757, A3 => n6756, A4 => 
                           n6755, ZN => n6764);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n7406, B1 => 
                           REGISTERS_13_27_port, B2 => n7394, ZN => n6762);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_15_27_port, A2 => n7407, B1 => 
                           REGISTERS_12_27_port, B2 => n7396, ZN => n6761);
   U2216 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n7357, B1 => 
                           REGISTERS_14_27_port, B2 => n7399, ZN => n6760);
   U2217 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n7395, B1 => 
                           REGISTERS_10_27_port, B2 => n7358, ZN => n6759);
   U2218 : NAND4_X1 port map( A1 => n6762, A2 => n6761, A3 => n6760, A4 => 
                           n6759, ZN => n6763);
   U2219 : AOI22_X1 port map( A1 => n7234, A2 => n6764, B1 => n7257, B2 => 
                           n6763, ZN => n6765);
   U2220 : OAI21_X1 port map( B1 => n7367, B2 => n6766, A => n6765, ZN => N412)
                           ;
   U2221 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n7374, B1 => 
                           REGISTERS_22_26_port, B2 => n7266, ZN => n6770);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n7371, B1 => 
                           REGISTERS_24_26_port, B2 => n7387, ZN => n6769);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n7315, B1 => 
                           REGISTERS_27_26_port, B2 => n7142, ZN => n6768);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_26_26_port, A2 => n7343, B1 => 
                           REGISTERS_17_26_port, B2 => n7383, ZN => n6767);
   U2225 : NAND4_X1 port map( A1 => n6770, A2 => n6769, A3 => n6768, A4 => 
                           n6767, ZN => n6776);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_31_26_port, A2 => n7373, B1 => 
                           REGISTERS_30_26_port, B2 => n7385, ZN => n6774);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n7375, B1 => 
                           REGISTERS_21_26_port, B2 => n7165, ZN => n6773);
   U2228 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n7368, B1 => 
                           REGISTERS_18_26_port, B2 => n7188, ZN => n6772);
   U2229 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n7285, B1 => 
                           REGISTERS_23_26_port, B2 => n7215, ZN => n6771);
   U2230 : NAND4_X1 port map( A1 => n6774, A2 => n6773, A3 => n6772, A4 => 
                           n6771, ZN => n6775);
   U2231 : NOR2_X1 port map( A1 => n6776, A2 => n6775, ZN => n6788);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_6_26_port, A2 => n7411, B1 => 
                           REGISTERS_0_26_port, B2 => n7406, ZN => n6780);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n7395, B1 => 
                           REGISTERS_7_26_port, B2 => n7296, ZN => n6779);
   U2234 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n7410, B1 => 
                           REGISTERS_3_26_port, B2 => n7350, ZN => n6778);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n7412, B1 => 
                           REGISTERS_2_26_port, B2 => n7358, ZN => n6777);
   U2236 : NAND4_X1 port map( A1 => n6780, A2 => n6779, A3 => n6778, A4 => 
                           n6777, ZN => n6786);
   U2237 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n7397, B1 => 
                           REGISTERS_9_26_port, B2 => n7409, ZN => n6784);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n7296, B1 => 
                           REGISTERS_12_26_port, B2 => n7396, ZN => n6783);
   U2239 : AOI22_X1 port map( A1 => REGISTERS_10_26_port, A2 => n7398, B1 => 
                           REGISTERS_14_26_port, B2 => n7322, ZN => n6782);
   U2240 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n7357, B1 => 
                           REGISTERS_13_26_port, B2 => n7394, ZN => n6781);
   U2241 : NAND4_X1 port map( A1 => n6784, A2 => n6783, A3 => n6782, A4 => 
                           n6781, ZN => n6785);
   U2242 : AOI22_X1 port map( A1 => n7234, A2 => n6786, B1 => n7257, B2 => 
                           n6785, ZN => n6787);
   U2243 : OAI21_X1 port map( B1 => n7367, B2 => n6788, A => n6787, ZN => N411)
                           ;
   U2244 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n7370, B1 => 
                           REGISTERS_17_25_port, B2 => n7383, ZN => n6792);
   U2245 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n7371, B1 => 
                           REGISTERS_26_25_port, B2 => n7343, ZN => n6791);
   U2246 : AOI22_X1 port map( A1 => REGISTERS_22_25_port, A2 => n7382, B1 => 
                           REGISTERS_16_25_port, B2 => n7285, ZN => n6790);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_18_25_port, A2 => n7381, B1 => 
                           REGISTERS_28_25_port, B2 => n7009, ZN => n6789);
   U2248 : NAND4_X1 port map( A1 => n6792, A2 => n6791, A3 => n6790, A4 => 
                           n6789, ZN => n6798);
   U2249 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n7374, B1 => 
                           REGISTERS_30_25_port, B2 => n7385, ZN => n6796);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n7338, B1 => 
                           REGISTERS_29_25_port, B2 => n7315, ZN => n6795);
   U2251 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n7375, B1 => 
                           REGISTERS_23_25_port, B2 => n7215, ZN => n6794);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n7337, B1 => 
                           REGISTERS_27_25_port, B2 => n7142, ZN => n6793);
   U2253 : NAND4_X1 port map( A1 => n6796, A2 => n6795, A3 => n6794, A4 => 
                           n6793, ZN => n6797);
   U2254 : NOR2_X1 port map( A1 => n6798, A2 => n6797, ZN => n6810);
   U2255 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n7357, B1 => 
                           REGISTERS_4_25_port, B2 => n7251, ZN => n6802);
   U2256 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n7400, B1 => 
                           REGISTERS_0_25_port, B2 => n7397, ZN => n6801);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n7412, B1 => 
                           REGISTERS_6_25_port, B2 => n7399, ZN => n6800);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_2_25_port, A2 => n7398, B1 => 
                           REGISTERS_1_25_port, B2 => n7409, ZN => n6799);
   U2259 : NAND4_X1 port map( A1 => n6802, A2 => n6801, A3 => n6800, A4 => 
                           n6799, ZN => n6808);
   U2260 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n7410, B1 => 
                           REGISTERS_10_25_port, B2 => n7358, ZN => n6806);
   U2261 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n7357, B1 => 
                           REGISTERS_14_25_port, B2 => n7322, ZN => n6805);
   U2262 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n7395, B1 => 
                           REGISTERS_13_25_port, B2 => n7227, ZN => n6804);
   U2263 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n7406, B1 => 
                           REGISTERS_15_25_port, B2 => n7407, ZN => n6803);
   U2264 : NAND4_X1 port map( A1 => n6806, A2 => n6805, A3 => n6804, A4 => 
                           n6803, ZN => n6807);
   U2265 : AOI22_X1 port map( A1 => n7234, A2 => n6808, B1 => n7257, B2 => 
                           n6807, ZN => n6809);
   U2266 : OAI21_X1 port map( B1 => n7367, B2 => n6810, A => n6809, ZN => N410)
                           ;
   U2267 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n7369, B1 => 
                           REGISTERS_28_24_port, B2 => n7009, ZN => n6814);
   U2268 : AOI22_X1 port map( A1 => REGISTERS_26_24_port, A2 => n7343, B1 => 
                           REGISTERS_25_24_port, B2 => n7216, ZN => n6813);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_19_24_port, A2 => n7336, B1 => 
                           REGISTERS_21_24_port, B2 => n7165, ZN => n6812);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n7381, B1 => 
                           REGISTERS_24_24_port, B2 => n7337, ZN => n6811);
   U2271 : NAND4_X1 port map( A1 => n6814, A2 => n6813, A3 => n6812, A4 => 
                           n6811, ZN => n6820);
   U2272 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n7335, B1 => 
                           REGISTERS_16_24_port, B2 => n7285, ZN => n6818);
   U2273 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n7384, B1 => 
                           REGISTERS_31_24_port, B2 => n7373, ZN => n6817);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_30_24_port, A2 => n7309, B1 => 
                           REGISTERS_20_24_port, B2 => n7314, ZN => n6816);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n7315, B1 => 
                           REGISTERS_22_24_port, B2 => n7266, ZN => n6815);
   U2276 : NAND4_X1 port map( A1 => n6818, A2 => n6817, A3 => n6816, A4 => 
                           n6815, ZN => n6819);
   U2277 : NOR2_X1 port map( A1 => n6820, A2 => n6819, ZN => n6832);
   U2278 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n7296, B1 => 
                           REGISTERS_4_24_port, B2 => n7396, ZN => n6824);
   U2279 : AOI22_X1 port map( A1 => REGISTERS_6_24_port, A2 => n7411, B1 => 
                           REGISTERS_3_24_port, B2 => n7408, ZN => n6823);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_2_24_port, A2 => n7405, B1 => 
                           REGISTERS_0_24_port, B2 => n7397, ZN => n6822);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n7395, B1 => 
                           REGISTERS_5_24_port, B2 => n7394, ZN => n6821);
   U2282 : NAND4_X1 port map( A1 => n6824, A2 => n6823, A3 => n6822, A4 => 
                           n6821, ZN => n6830);
   U2283 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n7351, B1 => 
                           REGISTERS_12_24_port, B2 => n7251, ZN => n6828);
   U2284 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n7409, B1 => 
                           REGISTERS_14_24_port, B2 => n7399, ZN => n6827);
   U2285 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n7357, B1 => 
                           REGISTERS_15_24_port, B2 => n7407, ZN => n6826);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n7412, B1 => 
                           REGISTERS_10_24_port, B2 => n7358, ZN => n6825);
   U2287 : NAND4_X1 port map( A1 => n6828, A2 => n6827, A3 => n6826, A4 => 
                           n6825, ZN => n6829);
   U2288 : AOI22_X1 port map( A1 => n7234, A2 => n6830, B1 => n7257, B2 => 
                           n6829, ZN => n6831);
   U2289 : OAI21_X1 port map( B1 => n7367, B2 => n6832, A => n6831, ZN => N409)
                           ;
   U2290 : AOI22_X1 port map( A1 => REGISTERS_23_23_port, A2 => n7384, B1 => 
                           REGISTERS_20_23_port, B2 => n7371, ZN => n6836);
   U2291 : AOI22_X1 port map( A1 => REGISTERS_30_23_port, A2 => n7385, B1 => 
                           REGISTERS_29_23_port, B2 => n7315, ZN => n6835);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n7374, B1 => 
                           REGISTERS_18_23_port, B2 => n7188, ZN => n6834);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_26_23_port, A2 => n7343, B1 => 
                           REGISTERS_24_23_port, B2 => n7337, ZN => n6833);
   U2294 : NAND4_X1 port map( A1 => n6836, A2 => n6835, A3 => n6834, A4 => 
                           n6833, ZN => n6842);
   U2295 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n7285, B1 => 
                           REGISTERS_21_23_port, B2 => n7165, ZN => n6840);
   U2296 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n7368, B1 => 
                           REGISTERS_17_23_port, B2 => n7383, ZN => n6839);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n7336, B1 => 
                           REGISTERS_22_23_port, B2 => n7266, ZN => n6838);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_31_23_port, A2 => n7373, B1 => 
                           REGISTERS_27_23_port, B2 => n7142, ZN => n6837);
   U2299 : NAND4_X1 port map( A1 => n6840, A2 => n6839, A3 => n6838, A4 => 
                           n6837, ZN => n6841);
   U2300 : NOR2_X1 port map( A1 => n6842, A2 => n6841, ZN => n6854);
   U2301 : AOI22_X1 port map( A1 => REGISTERS_6_23_port, A2 => n7411, B1 => 
                           REGISTERS_4_23_port, B2 => n7396, ZN => n6846);
   U2302 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n7412, B1 => 
                           REGISTERS_1_23_port, B2 => n7356, ZN => n6845);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n7407, B1 => 
                           REGISTERS_3_23_port, B2 => n7350, ZN => n6844);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n7397, B1 => 
                           REGISTERS_2_23_port, B2 => n7405, ZN => n6843);
   U2305 : NAND4_X1 port map( A1 => n6846, A2 => n6845, A3 => n6844, A4 => 
                           n6843, ZN => n6852);
   U2306 : AOI22_X1 port map( A1 => REGISTERS_14_23_port, A2 => n7411, B1 => 
                           REGISTERS_9_23_port, B2 => n7409, ZN => n6850);
   U2307 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n7407, B1 => 
                           REGISTERS_13_23_port, B2 => n7227, ZN => n6849);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n7406, B1 => 
                           REGISTERS_10_23_port, B2 => n7358, ZN => n6848);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n7251, B1 => 
                           REGISTERS_11_23_port, B2 => n7408, ZN => n6847);
   U2310 : NAND4_X1 port map( A1 => n6850, A2 => n6849, A3 => n6848, A4 => 
                           n6847, ZN => n6851);
   U2311 : AOI22_X1 port map( A1 => n7234, A2 => n6852, B1 => n7257, B2 => 
                           n6851, ZN => n6853);
   U2312 : OAI21_X1 port map( B1 => n7423, B2 => n6854, A => n6853, ZN => N408)
                           ;
   U2313 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n7374, B1 => 
                           REGISTERS_31_22_port, B2 => n7373, ZN => n6858);
   U2314 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n7384, B1 => 
                           REGISTERS_18_22_port, B2 => n7188, ZN => n6857);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_26_22_port, A2 => n7343, B1 => 
                           REGISTERS_27_22_port, B2 => n7142, ZN => n6856);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n7368, B1 => 
                           REGISTERS_21_22_port, B2 => n7165, ZN => n6855);
   U2317 : NAND4_X1 port map( A1 => n6858, A2 => n6857, A3 => n6856, A4 => 
                           n6855, ZN => n6864);
   U2318 : AOI22_X1 port map( A1 => REGISTERS_30_22_port, A2 => n7309, B1 => 
                           REGISTERS_29_22_port, B2 => n7315, ZN => n6862);
   U2319 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n7337, B1 => 
                           REGISTERS_17_22_port, B2 => n7383, ZN => n6861);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_22_22_port, A2 => n7382, B1 => 
                           REGISTERS_20_22_port, B2 => n7371, ZN => n6860);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n7375, B1 => 
                           REGISTERS_16_22_port, B2 => n7285, ZN => n6859);
   U2322 : NAND4_X1 port map( A1 => n6862, A2 => n6861, A3 => n6860, A4 => 
                           n6859, ZN => n6863);
   U2323 : NOR2_X1 port map( A1 => n6864, A2 => n6863, ZN => n6876);
   U2324 : AOI22_X1 port map( A1 => REGISTERS_2_22_port, A2 => n7398, B1 => 
                           REGISTERS_0_22_port, B2 => n7406, ZN => n6868);
   U2325 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n7357, B1 => 
                           REGISTERS_6_22_port, B2 => n7322, ZN => n6867);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n7409, B1 => 
                           REGISTERS_4_22_port, B2 => n7251, ZN => n6866);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n7227, B1 => 
                           REGISTERS_7_22_port, B2 => n7296, ZN => n6865);
   U2328 : NAND4_X1 port map( A1 => n6868, A2 => n6867, A3 => n6866, A4 => 
                           n6865, ZN => n6874);
   U2329 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n7396, B1 => 
                           REGISTERS_15_22_port, B2 => n7407, ZN => n6872);
   U2330 : AOI22_X1 port map( A1 => REGISTERS_14_22_port, A2 => n7399, B1 => 
                           REGISTERS_11_22_port, B2 => n7350, ZN => n6871);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n7397, B1 => 
                           REGISTERS_10_22_port, B2 => n7405, ZN => n6870);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n7412, B1 => 
                           REGISTERS_9_22_port, B2 => n7356, ZN => n6869);
   U2333 : NAND4_X1 port map( A1 => n6872, A2 => n6871, A3 => n6870, A4 => 
                           n6869, ZN => n6873);
   U2334 : AOI22_X1 port map( A1 => n7234, A2 => n6874, B1 => n7257, B2 => 
                           n6873, ZN => n6875);
   U2335 : OAI21_X1 port map( B1 => n7423, B2 => n6876, A => n6875, ZN => N407)
                           ;
   U2336 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n7337, B1 => 
                           REGISTERS_30_21_port, B2 => n7385, ZN => n6880);
   U2337 : AOI22_X1 port map( A1 => REGISTERS_23_21_port, A2 => n7384, B1 => 
                           REGISTERS_31_21_port, B2 => n7373, ZN => n6879);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n7374, B1 => 
                           REGISTERS_18_21_port, B2 => n7188, ZN => n6878);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n7009, B1 => 
                           REGISTERS_27_21_port, B2 => n7142, ZN => n6877);
   U2340 : NAND4_X1 port map( A1 => n6880, A2 => n6879, A3 => n6878, A4 => 
                           n6877, ZN => n6886);
   U2341 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n7285, B1 => 
                           REGISTERS_20_21_port, B2 => n7371, ZN => n6884);
   U2342 : AOI22_X1 port map( A1 => REGISTERS_26_21_port, A2 => n7343, B1 => 
                           REGISTERS_19_21_port, B2 => n7375, ZN => n6883);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n7382, B1 => 
                           REGISTERS_29_21_port, B2 => n7380, ZN => n6882);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n7370, B1 => 
                           REGISTERS_17_21_port, B2 => n7383, ZN => n6881);
   U2345 : NAND4_X1 port map( A1 => n6884, A2 => n6883, A3 => n6882, A4 => 
                           n6881, ZN => n6885);
   U2346 : NOR2_X1 port map( A1 => n6886, A2 => n6885, ZN => n6898);
   U2347 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n7394, B1 => 
                           REGISTERS_2_21_port, B2 => n7358, ZN => n6890);
   U2348 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n7395, B1 => 
                           REGISTERS_3_21_port, B2 => n7408, ZN => n6889);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n7296, B1 => 
                           REGISTERS_6_21_port, B2 => n7399, ZN => n6888);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n7351, B1 => 
                           REGISTERS_4_21_port, B2 => n7396, ZN => n6887);
   U2351 : NAND4_X1 port map( A1 => n6890, A2 => n6889, A3 => n6888, A4 => 
                           n6887, ZN => n6896);
   U2352 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n7397, B1 => 
                           REGISTERS_10_21_port, B2 => n7405, ZN => n6894);
   U2353 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n7227, B1 => 
                           REGISTERS_11_21_port, B2 => n7350, ZN => n6893);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n7407, B1 => 
                           REGISTERS_14_21_port, B2 => n7322, ZN => n6892);
   U2355 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n7395, B1 => 
                           REGISTERS_12_21_port, B2 => n7251, ZN => n6891);
   U2356 : NAND4_X1 port map( A1 => n6894, A2 => n6893, A3 => n6892, A4 => 
                           n6891, ZN => n6895);
   U2357 : AOI22_X1 port map( A1 => n7234, A2 => n6896, B1 => n7257, B2 => 
                           n6895, ZN => n6897);
   U2358 : OAI21_X1 port map( B1 => n7423, B2 => n6898, A => n6897, ZN => N406)
                           ;
   U2359 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n7285, B1 => 
                           REGISTERS_18_20_port, B2 => n7188, ZN => n6902);
   U2360 : AOI22_X1 port map( A1 => REGISTERS_22_20_port, A2 => n7266, B1 => 
                           REGISTERS_19_20_port, B2 => n7375, ZN => n6901);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n7165, B1 => 
                           REGISTERS_23_20_port, B2 => n7215, ZN => n6900);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_30_20_port, A2 => n7385, B1 => 
                           REGISTERS_20_20_port, B2 => n7371, ZN => n6899);
   U2363 : NAND4_X1 port map( A1 => n6902, A2 => n6901, A3 => n6900, A4 => 
                           n6899, ZN => n6908);
   U2364 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n7337, B1 => 
                           REGISTERS_17_20_port, B2 => n7383, ZN => n6906);
   U2365 : AOI22_X1 port map( A1 => REGISTERS_26_20_port, A2 => n7372, B1 => 
                           REGISTERS_31_20_port, B2 => n7373, ZN => n6905);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n7374, B1 => 
                           REGISTERS_27_20_port, B2 => n7142, ZN => n6904);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n7368, B1 => 
                           REGISTERS_29_20_port, B2 => n7315, ZN => n6903);
   U2368 : NAND4_X1 port map( A1 => n6906, A2 => n6905, A3 => n6904, A4 => 
                           n6903, ZN => n6907);
   U2369 : NOR2_X1 port map( A1 => n6908, A2 => n6907, ZN => n6920);
   U2370 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n7407, B1 => 
                           REGISTERS_4_20_port, B2 => n7396, ZN => n6912);
   U2371 : AOI22_X1 port map( A1 => REGISTERS_6_20_port, A2 => n7399, B1 => 
                           REGISTERS_5_20_port, B2 => n7394, ZN => n6911);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_2_20_port, A2 => n7358, B1 => 
                           REGISTERS_0_20_port, B2 => n7406, ZN => n6910);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_3_20_port, A2 => n7408, B1 => 
                           REGISTERS_1_20_port, B2 => n7409, ZN => n6909);
   U2374 : NAND4_X1 port map( A1 => n6912, A2 => n6911, A3 => n6910, A4 => 
                           n6909, ZN => n6918);
   U2375 : AOI22_X1 port map( A1 => REGISTERS_14_20_port, A2 => n7399, B1 => 
                           REGISTERS_9_20_port, B2 => n7356, ZN => n6916);
   U2376 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n7251, B1 => 
                           REGISTERS_10_20_port, B2 => n7358, ZN => n6915);
   U2377 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n7350, B1 => 
                           REGISTERS_15_20_port, B2 => n7296, ZN => n6914);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n7351, B1 => 
                           REGISTERS_13_20_port, B2 => n7227, ZN => n6913);
   U2379 : NAND4_X1 port map( A1 => n6916, A2 => n6915, A3 => n6914, A4 => 
                           n6913, ZN => n6917);
   U2380 : AOI22_X1 port map( A1 => n7234, A2 => n6918, B1 => n7418, B2 => 
                           n6917, ZN => n6919);
   U2381 : OAI21_X1 port map( B1 => n7423, B2 => n6920, A => n6919, ZN => N405)
                           ;
   U2382 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n7009, B1 => 
                           REGISTERS_23_19_port, B2 => n7215, ZN => n6924);
   U2383 : AOI22_X1 port map( A1 => REGISTERS_27_19_port, A2 => n7369, B1 => 
                           REGISTERS_21_19_port, B2 => n7165, ZN => n6923);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n7315, B1 => 
                           REGISTERS_31_19_port, B2 => n7373, ZN => n6922);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n7371, B1 => 
                           REGISTERS_19_19_port, B2 => n7375, ZN => n6921);
   U2386 : NAND4_X1 port map( A1 => n6924, A2 => n6923, A3 => n6922, A4 => 
                           n6921, ZN => n6930);
   U2387 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n7285, B1 => 
                           REGISTERS_26_19_port, B2 => n7343, ZN => n6928);
   U2388 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n7337, B1 => 
                           REGISTERS_25_19_port, B2 => n7216, ZN => n6927);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_22_19_port, A2 => n7382, B1 => 
                           REGISTERS_17_19_port, B2 => n7335, ZN => n6926);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_18_19_port, A2 => n7381, B1 => 
                           REGISTERS_30_19_port, B2 => n7385, ZN => n6925);
   U2391 : NAND4_X1 port map( A1 => n6928, A2 => n6927, A3 => n6926, A4 => 
                           n6925, ZN => n6929);
   U2392 : NOR2_X1 port map( A1 => n6930, A2 => n6929, ZN => n6942);
   U2393 : CLKBUF_X1 port map( A => n7420, Z => n7259);
   U2394 : AOI22_X1 port map( A1 => REGISTERS_2_19_port, A2 => n7398, B1 => 
                           REGISTERS_1_19_port, B2 => n7409, ZN => n6934);
   U2395 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n7397, B1 => 
                           REGISTERS_4_19_port, B2 => n7251, ZN => n6933);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n7227, B1 => 
                           REGISTERS_7_19_port, B2 => n7296, ZN => n6932);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_6_19_port, A2 => n7411, B1 => 
                           REGISTERS_3_19_port, B2 => n7408, ZN => n6931);
   U2398 : NAND4_X1 port map( A1 => n6934, A2 => n6933, A3 => n6932, A4 => 
                           n6931, ZN => n6940);
   U2399 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n7409, B1 => 
                           REGISTERS_14_19_port, B2 => n7399, ZN => n6938);
   U2400 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n7408, B1 => 
                           REGISTERS_8_19_port, B2 => n7351, ZN => n6937);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_10_19_port, A2 => n7358, B1 => 
                           REGISTERS_13_19_port, B2 => n7394, ZN => n6936);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n7396, B1 => 
                           REGISTERS_15_19_port, B2 => n7400, ZN => n6935);
   U2403 : NAND4_X1 port map( A1 => n6938, A2 => n6937, A3 => n6936, A4 => 
                           n6935, ZN => n6939);
   U2404 : AOI22_X1 port map( A1 => n7259, A2 => n6940, B1 => n7257, B2 => 
                           n6939, ZN => n6941);
   U2405 : OAI21_X1 port map( B1 => n7423, B2 => n6942, A => n6941, ZN => N404)
                           ;
   U2406 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n7386, B1 => 
                           REGISTERS_17_18_port, B2 => n7335, ZN => n6946);
   U2407 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n7387, B1 => 
                           REGISTERS_18_18_port, B2 => n7188, ZN => n6945);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_31_18_port, A2 => n7373, B1 => 
                           REGISTERS_20_18_port, B2 => n7371, ZN => n6944);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n7009, B1 => 
                           REGISTERS_27_18_port, B2 => n7369, ZN => n6943);
   U2410 : NAND4_X1 port map( A1 => n6946, A2 => n6945, A3 => n6944, A4 => 
                           n6943, ZN => n6952);
   U2411 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n7380, B1 => 
                           REGISTERS_23_18_port, B2 => n7215, ZN => n6950);
   U2412 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n7374, B1 => 
                           REGISTERS_22_18_port, B2 => n7266, ZN => n6949);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n7165, B1 => 
                           REGISTERS_30_18_port, B2 => n7385, ZN => n6948);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n7375, B1 => 
                           REGISTERS_26_18_port, B2 => n7372, ZN => n6947);
   U2415 : NAND4_X1 port map( A1 => n6950, A2 => n6949, A3 => n6948, A4 => 
                           n6947, ZN => n6951);
   U2416 : NOR2_X1 port map( A1 => n6952, A2 => n6951, ZN => n6964);
   U2417 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n7357, B1 => 
                           REGISTERS_2_18_port, B2 => n7405, ZN => n6956);
   U2418 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n7400, B1 => 
                           REGISTERS_1_18_port, B2 => n7356, ZN => n6955);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n7412, B1 => 
                           REGISTERS_6_18_port, B2 => n7322, ZN => n6954);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n7406, B1 => 
                           REGISTERS_4_18_port, B2 => n7396, ZN => n6953);
   U2421 : NAND4_X1 port map( A1 => n6956, A2 => n6955, A3 => n6954, A4 => 
                           n6953, ZN => n6962);
   U2422 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n7356, B1 => 
                           REGISTERS_8_18_port, B2 => n7351, ZN => n6960);
   U2423 : AOI22_X1 port map( A1 => REGISTERS_14_18_port, A2 => n7399, B1 => 
                           REGISTERS_11_18_port, B2 => n7350, ZN => n6959);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n7227, B1 => 
                           REGISTERS_12_18_port, B2 => n7251, ZN => n6958);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_10_18_port, A2 => n7398, B1 => 
                           REGISTERS_15_18_port, B2 => n7400, ZN => n6957);
   U2426 : NAND4_X1 port map( A1 => n6960, A2 => n6959, A3 => n6958, A4 => 
                           n6957, ZN => n6961);
   U2427 : AOI22_X1 port map( A1 => n7259, A2 => n6962, B1 => n7257, B2 => 
                           n6961, ZN => n6963);
   U2428 : OAI21_X1 port map( B1 => n7423, B2 => n6964, A => n6963, ZN => N403)
                           ;
   U2429 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n7216, B1 => 
                           REGISTERS_26_17_port, B2 => n7343, ZN => n6968);
   U2430 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n7314, B1 => 
                           REGISTERS_17_17_port, B2 => n7335, ZN => n6967);
   U2431 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n7215, B1 => 
                           REGISTERS_16_17_port, B2 => n7285, ZN => n6966);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n7387, B1 => 
                           REGISTERS_30_17_port, B2 => n7385, ZN => n6965);
   U2433 : NAND4_X1 port map( A1 => n6968, A2 => n6967, A3 => n6966, A4 => 
                           n6965, ZN => n6974);
   U2434 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n7380, B1 => 
                           REGISTERS_28_17_port, B2 => n7009, ZN => n6972);
   U2435 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n7370, B1 => 
                           REGISTERS_27_17_port, B2 => n7369, ZN => n6971);
   U2436 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n7373, B1 => 
                           REGISTERS_19_17_port, B2 => n7375, ZN => n6970);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_22_17_port, A2 => n7382, B1 => 
                           REGISTERS_18_17_port, B2 => n7188, ZN => n6969);
   U2438 : NAND4_X1 port map( A1 => n6972, A2 => n6971, A3 => n6970, A4 => 
                           n6969, ZN => n6973);
   U2439 : NOR2_X1 port map( A1 => n6974, A2 => n6973, ZN => n6986);
   U2440 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n7251, B1 => 
                           REGISTERS_0_17_port, B2 => n7351, ZN => n6978);
   U2441 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n7227, B1 => 
                           REGISTERS_3_17_port, B2 => n7408, ZN => n6977);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n7322, B1 => 
                           REGISTERS_1_17_port, B2 => n7409, ZN => n6976);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n7296, B1 => 
                           REGISTERS_2_17_port, B2 => n7358, ZN => n6975);
   U2444 : NAND4_X1 port map( A1 => n6978, A2 => n6977, A3 => n6976, A4 => 
                           n6975, ZN => n6984);
   U2445 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n7410, B1 => 
                           REGISTERS_9_17_port, B2 => n7356, ZN => n6982);
   U2446 : AOI22_X1 port map( A1 => REGISTERS_14_17_port, A2 => n7322, B1 => 
                           REGISTERS_11_17_port, B2 => n7350, ZN => n6981);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n7351, B1 => 
                           REGISTERS_15_17_port, B2 => n7407, ZN => n6980);
   U2448 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n7398, B1 => 
                           REGISTERS_13_17_port, B2 => n7227, ZN => n6979);
   U2449 : NAND4_X1 port map( A1 => n6982, A2 => n6981, A3 => n6980, A4 => 
                           n6979, ZN => n6983);
   U2450 : AOI22_X1 port map( A1 => n7259, A2 => n6984, B1 => n7257, B2 => 
                           n6983, ZN => n6985);
   U2451 : OAI21_X1 port map( B1 => n7423, B2 => n6986, A => n6985, ZN => N402)
                           ;
   U2452 : AOI22_X1 port map( A1 => REGISTERS_26_16_port, A2 => n7372, B1 => 
                           REGISTERS_22_16_port, B2 => n7266, ZN => n6990);
   U2453 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n7386, B1 => 
                           REGISTERS_19_16_port, B2 => n7336, ZN => n6989);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n7370, B1 => 
                           REGISTERS_18_16_port, B2 => n7188, ZN => n6988);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n7380, B1 => 
                           REGISTERS_27_16_port, B2 => n7369, ZN => n6987);
   U2456 : NAND4_X1 port map( A1 => n6990, A2 => n6989, A3 => n6988, A4 => 
                           n6987, ZN => n6996);
   U2457 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n7215, B1 => 
                           REGISTERS_31_16_port, B2 => n7373, ZN => n6994);
   U2458 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n7314, B1 => 
                           REGISTERS_25_16_port, B2 => n7216, ZN => n6993);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n7337, B1 => 
                           REGISTERS_28_16_port, B2 => n7009, ZN => n6992);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n7335, B1 => 
                           REGISTERS_30_16_port, B2 => n7385, ZN => n6991);
   U2461 : NAND4_X1 port map( A1 => n6994, A2 => n6993, A3 => n6992, A4 => 
                           n6991, ZN => n6995);
   U2462 : NOR2_X1 port map( A1 => n6996, A2 => n6995, ZN => n7008);
   U2463 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n7408, B1 => 
                           REGISTERS_5_16_port, B2 => n7394, ZN => n7000);
   U2464 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n7409, B1 => 
                           REGISTERS_4_16_port, B2 => n7251, ZN => n6999);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n7407, B1 => 
                           REGISTERS_0_16_port, B2 => n7406, ZN => n6998);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_6_16_port, A2 => n7411, B1 => 
                           REGISTERS_2_16_port, B2 => n7405, ZN => n6997);
   U2467 : NAND4_X1 port map( A1 => n7000, A2 => n6999, A3 => n6998, A4 => 
                           n6997, ZN => n7006);
   U2468 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n7397, B1 => 
                           REGISTERS_12_16_port, B2 => n7396, ZN => n7004);
   U2469 : AOI22_X1 port map( A1 => REGISTERS_14_16_port, A2 => n7411, B1 => 
                           REGISTERS_13_16_port, B2 => n7227, ZN => n7003);
   U2470 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n7358, B1 => 
                           REGISTERS_11_16_port, B2 => n7350, ZN => n7002);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n7400, B1 => 
                           REGISTERS_9_16_port, B2 => n7409, ZN => n7001);
   U2472 : NAND4_X1 port map( A1 => n7004, A2 => n7003, A3 => n7002, A4 => 
                           n7001, ZN => n7005);
   U2473 : AOI22_X1 port map( A1 => n7259, A2 => n7006, B1 => n7257, B2 => 
                           n7005, ZN => n7007);
   U2474 : OAI21_X1 port map( B1 => n7423, B2 => n7008, A => n7007, ZN => N401)
                           ;
   U2475 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n7142, B1 => 
                           REGISTERS_22_15_port, B2 => n7266, ZN => n7013);
   U2476 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n7386, B1 => 
                           REGISTERS_18_15_port, B2 => n7381, ZN => n7012);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_26_15_port, A2 => n7343, B1 => 
                           REGISTERS_31_15_port, B2 => n7373, ZN => n7011);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n7383, B1 => 
                           REGISTERS_28_15_port, B2 => n7009, ZN => n7010);
   U2479 : NAND4_X1 port map( A1 => n7013, A2 => n7012, A3 => n7011, A4 => 
                           n7010, ZN => n7019);
   U2480 : AOI22_X1 port map( A1 => REGISTERS_30_15_port, A2 => n7385, B1 => 
                           REGISTERS_20_15_port, B2 => n7371, ZN => n7017);
   U2481 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n7315, B1 => 
                           REGISTERS_21_15_port, B2 => n7165, ZN => n7016);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n7337, B1 => 
                           REGISTERS_25_15_port, B2 => n7216, ZN => n7015);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n7384, B1 => 
                           REGISTERS_19_15_port, B2 => n7375, ZN => n7014);
   U2484 : NAND4_X1 port map( A1 => n7017, A2 => n7016, A3 => n7015, A4 => 
                           n7014, ZN => n7018);
   U2485 : NOR2_X1 port map( A1 => n7019, A2 => n7018, ZN => n7031);
   U2486 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n7396, B1 => 
                           REGISTERS_1_15_port, B2 => n7356, ZN => n7023);
   U2487 : AOI22_X1 port map( A1 => REGISTERS_3_15_port, A2 => n7350, B1 => 
                           REGISTERS_2_15_port, B2 => n7358, ZN => n7022);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n7406, B1 => 
                           REGISTERS_5_15_port, B2 => n7394, ZN => n7021);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_6_15_port, A2 => n7411, B1 => 
                           REGISTERS_7_15_port, B2 => n7400, ZN => n7020);
   U2490 : NAND4_X1 port map( A1 => n7023, A2 => n7022, A3 => n7021, A4 => 
                           n7020, ZN => n7029);
   U2491 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n7395, B1 => 
                           REGISTERS_8_15_port, B2 => n7351, ZN => n7027);
   U2492 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n7296, B1 => 
                           REGISTERS_12_15_port, B2 => n7251, ZN => n7026);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_14_15_port, A2 => n7411, B1 => 
                           REGISTERS_13_15_port, B2 => n7227, ZN => n7025);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n7357, B1 => 
                           REGISTERS_10_15_port, B2 => n7405, ZN => n7024);
   U2495 : NAND4_X1 port map( A1 => n7027, A2 => n7026, A3 => n7025, A4 => 
                           n7024, ZN => n7028);
   U2496 : AOI22_X1 port map( A1 => n7259, A2 => n7029, B1 => n7257, B2 => 
                           n7028, ZN => n7030);
   U2497 : OAI21_X1 port map( B1 => n7367, B2 => n7031, A => n7030, ZN => N400)
                           ;
   U2498 : AOI22_X1 port map( A1 => REGISTERS_18_14_port, A2 => n7381, B1 => 
                           REGISTERS_25_14_port, B2 => n7216, ZN => n7035);
   U2499 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n7337, B1 => 
                           REGISTERS_30_14_port, B2 => n7385, ZN => n7034);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n7370, B1 => 
                           REGISTERS_19_14_port, B2 => n7375, ZN => n7033);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n7382, B1 => 
                           REGISTERS_28_14_port, B2 => n7368, ZN => n7032);
   U2502 : NAND4_X1 port map( A1 => n7035, A2 => n7034, A3 => n7033, A4 => 
                           n7032, ZN => n7041);
   U2503 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n7314, B1 => 
                           REGISTERS_29_14_port, B2 => n7315, ZN => n7039);
   U2504 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n7383, B1 => 
                           REGISTERS_31_14_port, B2 => n7373, ZN => n7038);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n7285, B1 => 
                           REGISTERS_26_14_port, B2 => n7343, ZN => n7037);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_23_14_port, A2 => n7384, B1 => 
                           REGISTERS_27_14_port, B2 => n7369, ZN => n7036);
   U2507 : NAND4_X1 port map( A1 => n7039, A2 => n7038, A3 => n7037, A4 => 
                           n7036, ZN => n7040);
   U2508 : NOR2_X1 port map( A1 => n7041, A2 => n7040, ZN => n7053);
   U2509 : AOI22_X1 port map( A1 => REGISTERS_2_14_port, A2 => n7405, B1 => 
                           REGISTERS_7_14_port, B2 => n7407, ZN => n7045);
   U2510 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n7356, B1 => 
                           REGISTERS_3_14_port, B2 => n7408, ZN => n7044);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n7351, B1 => 
                           REGISTERS_6_14_port, B2 => n7399, ZN => n7043);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n7394, B1 => 
                           REGISTERS_4_14_port, B2 => n7396, ZN => n7042);
   U2513 : NAND4_X1 port map( A1 => n7045, A2 => n7044, A3 => n7043, A4 => 
                           n7042, ZN => n7051);
   U2514 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n7251, B1 => 
                           REGISTERS_9_14_port, B2 => n7356, ZN => n7049);
   U2515 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n7408, B1 => 
                           REGISTERS_15_14_port, B2 => n7296, ZN => n7048);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n7412, B1 => 
                           REGISTERS_14_14_port, B2 => n7399, ZN => n7047);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n7397, B1 => 
                           REGISTERS_10_14_port, B2 => n7405, ZN => n7046);
   U2518 : NAND4_X1 port map( A1 => n7049, A2 => n7048, A3 => n7047, A4 => 
                           n7046, ZN => n7050);
   U2519 : AOI22_X1 port map( A1 => n7259, A2 => n7051, B1 => n7257, B2 => 
                           n7050, ZN => n7052);
   U2520 : OAI21_X1 port map( B1 => n7423, B2 => n7053, A => n7052, ZN => N399)
                           ;
   U2521 : AOI22_X1 port map( A1 => REGISTERS_26_13_port, A2 => n7343, B1 => 
                           REGISTERS_28_13_port, B2 => n7368, ZN => n7057);
   U2522 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n7285, B1 => 
                           REGISTERS_18_13_port, B2 => n7381, ZN => n7056);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n7374, B1 => 
                           REGISTERS_24_13_port, B2 => n7337, ZN => n7055);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n7371, B1 => 
                           REGISTERS_30_13_port, B2 => n7385, ZN => n7054);
   U2525 : NAND4_X1 port map( A1 => n7057, A2 => n7056, A3 => n7055, A4 => 
                           n7054, ZN => n7063);
   U2526 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n7384, B1 => 
                           REGISTERS_22_13_port, B2 => n7266, ZN => n7061);
   U2527 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n7375, B1 => 
                           REGISTERS_17_13_port, B2 => n7335, ZN => n7060);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n7315, B1 => 
                           REGISTERS_27_13_port, B2 => n7369, ZN => n7059);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n7370, B1 => 
                           REGISTERS_31_13_port, B2 => n7373, ZN => n7058);
   U2530 : NAND4_X1 port map( A1 => n7061, A2 => n7060, A3 => n7059, A4 => 
                           n7058, ZN => n7062);
   U2531 : NOR2_X1 port map( A1 => n7063, A2 => n7062, ZN => n7075);
   U2532 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n7410, B1 => 
                           REGISTERS_7_13_port, B2 => n7407, ZN => n7067);
   U2533 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n7406, B1 => 
                           REGISTERS_1_13_port, B2 => n7409, ZN => n7066);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_2_13_port, A2 => n7405, B1 => 
                           REGISTERS_6_13_port, B2 => n7322, ZN => n7065);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n7394, B1 => 
                           REGISTERS_3_13_port, B2 => n7350, ZN => n7064);
   U2536 : NAND4_X1 port map( A1 => n7067, A2 => n7066, A3 => n7065, A4 => 
                           n7064, ZN => n7073);
   U2537 : AOI22_X1 port map( A1 => REGISTERS_11_13_port, A2 => n7357, B1 => 
                           REGISTERS_12_13_port, B2 => n7251, ZN => n7071);
   U2538 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n7356, B1 => 
                           REGISTERS_13_13_port, B2 => n7227, ZN => n7070);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n7397, B1 => 
                           REGISTERS_14_13_port, B2 => n7399, ZN => n7069);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_10_13_port, A2 => n7398, B1 => 
                           REGISTERS_15_13_port, B2 => n7296, ZN => n7068);
   U2541 : NAND4_X1 port map( A1 => n7071, A2 => n7070, A3 => n7069, A4 => 
                           n7068, ZN => n7072);
   U2542 : AOI22_X1 port map( A1 => n7259, A2 => n7073, B1 => n7257, B2 => 
                           n7072, ZN => n7074);
   U2543 : OAI21_X1 port map( B1 => n7367, B2 => n7075, A => n7074, ZN => N398)
                           ;
   U2544 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n7285, B1 => 
                           REGISTERS_21_12_port, B2 => n7370, ZN => n7079);
   U2545 : AOI22_X1 port map( A1 => REGISTERS_18_12_port, A2 => n7381, B1 => 
                           REGISTERS_23_12_port, B2 => n7215, ZN => n7078);
   U2546 : AOI22_X1 port map( A1 => REGISTERS_26_12_port, A2 => n7343, B1 => 
                           REGISTERS_27_12_port, B2 => n7369, ZN => n7077);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_30_12_port, A2 => n7385, B1 => 
                           REGISTERS_28_12_port, B2 => n7368, ZN => n7076);
   U2548 : NAND4_X1 port map( A1 => n7079, A2 => n7078, A3 => n7077, A4 => 
                           n7076, ZN => n7085);
   U2549 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n7374, B1 => 
                           REGISTERS_31_12_port, B2 => n7338, ZN => n7083);
   U2550 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n7337, B1 => 
                           REGISTERS_20_12_port, B2 => n7314, ZN => n7082);
   U2551 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n7335, B1 => 
                           REGISTERS_22_12_port, B2 => n7266, ZN => n7081);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n7315, B1 => 
                           REGISTERS_19_12_port, B2 => n7336, ZN => n7080);
   U2553 : NAND4_X1 port map( A1 => n7083, A2 => n7082, A3 => n7081, A4 => 
                           n7080, ZN => n7084);
   U2554 : NOR2_X1 port map( A1 => n7085, A2 => n7084, ZN => n7097);
   U2555 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n7397, B1 => 
                           REGISTERS_4_12_port, B2 => n7396, ZN => n7089);
   U2556 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n7412, B1 => 
                           REGISTERS_2_12_port, B2 => n7358, ZN => n7088);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n7407, B1 => 
                           REGISTERS_6_12_port, B2 => n7322, ZN => n7087);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n7357, B1 => 
                           REGISTERS_1_12_port, B2 => n7356, ZN => n7086);
   U2559 : NAND4_X1 port map( A1 => n7089, A2 => n7088, A3 => n7087, A4 => 
                           n7086, ZN => n7095);
   U2560 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n7350, B1 => 
                           REGISTERS_13_12_port, B2 => n7394, ZN => n7093);
   U2561 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n7399, B1 => 
                           REGISTERS_9_12_port, B2 => n7409, ZN => n7092);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n7400, B1 => 
                           REGISTERS_12_12_port, B2 => n7410, ZN => n7091);
   U2563 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n7397, B1 => 
                           REGISTERS_10_12_port, B2 => n7405, ZN => n7090);
   U2564 : NAND4_X1 port map( A1 => n7093, A2 => n7092, A3 => n7091, A4 => 
                           n7090, ZN => n7094);
   U2565 : AOI22_X1 port map( A1 => n7259, A2 => n7095, B1 => n7257, B2 => 
                           n7094, ZN => n7096);
   U2566 : OAI21_X1 port map( B1 => n7423, B2 => n7097, A => n7096, ZN => N397)
                           ;
   U2567 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n7384, B1 => 
                           REGISTERS_22_11_port, B2 => n7382, ZN => n7101);
   U2568 : AOI22_X1 port map( A1 => REGISTERS_31_11_port, A2 => n7373, B1 => 
                           REGISTERS_24_11_port, B2 => n7387, ZN => n7100);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_18_11_port, A2 => n7188, B1 => 
                           REGISTERS_17_11_port, B2 => n7335, ZN => n7099);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n7285, B1 => 
                           REGISTERS_19_11_port, B2 => n7375, ZN => n7098);
   U2571 : NAND4_X1 port map( A1 => n7101, A2 => n7100, A3 => n7099, A4 => 
                           n7098, ZN => n7107);
   U2572 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n7370, B1 => 
                           REGISTERS_26_11_port, B2 => n7343, ZN => n7105);
   U2573 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n7315, B1 => 
                           REGISTERS_25_11_port, B2 => n7374, ZN => n7104);
   U2574 : AOI22_X1 port map( A1 => REGISTERS_27_11_port, A2 => n7142, B1 => 
                           REGISTERS_28_11_port, B2 => n7368, ZN => n7103);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_30_11_port, A2 => n7385, B1 => 
                           REGISTERS_20_11_port, B2 => n7371, ZN => n7102);
   U2576 : NAND4_X1 port map( A1 => n7105, A2 => n7104, A3 => n7103, A4 => 
                           n7102, ZN => n7106);
   U2577 : NOR2_X1 port map( A1 => n7107, A2 => n7106, ZN => n7119);
   U2578 : AOI22_X1 port map( A1 => REGISTERS_2_11_port, A2 => n7405, B1 => 
                           REGISTERS_5_11_port, B2 => n7227, ZN => n7111);
   U2579 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n7296, B1 => 
                           REGISTERS_1_11_port, B2 => n7356, ZN => n7110);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n7397, B1 => 
                           REGISTERS_6_11_port, B2 => n7399, ZN => n7109);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n7350, B1 => 
                           REGISTERS_4_11_port, B2 => n7251, ZN => n7108);
   U2582 : NAND4_X1 port map( A1 => n7111, A2 => n7110, A3 => n7109, A4 => 
                           n7108, ZN => n7117);
   U2583 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n7227, B1 => 
                           REGISTERS_14_11_port, B2 => n7322, ZN => n7115);
   U2584 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n7405, B1 => 
                           REGISTERS_12_11_port, B2 => n7251, ZN => n7114);
   U2585 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n7395, B1 => 
                           REGISTERS_15_11_port, B2 => n7296, ZN => n7113);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n7350, B1 => 
                           REGISTERS_8_11_port, B2 => n7351, ZN => n7112);
   U2587 : NAND4_X1 port map( A1 => n7115, A2 => n7114, A3 => n7113, A4 => 
                           n7112, ZN => n7116);
   U2588 : AOI22_X1 port map( A1 => n7259, A2 => n7117, B1 => n7257, B2 => 
                           n7116, ZN => n7118);
   U2589 : OAI21_X1 port map( B1 => n7423, B2 => n7119, A => n7118, ZN => N396)
                           ;
   U2590 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n7371, B1 => 
                           REGISTERS_17_10_port, B2 => n7335, ZN => n7123);
   U2591 : AOI22_X1 port map( A1 => REGISTERS_30_10_port, A2 => n7385, B1 => 
                           REGISTERS_31_10_port, B2 => n7338, ZN => n7122);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n7216, B1 => 
                           REGISTERS_22_10_port, B2 => n7382, ZN => n7121);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_26_10_port, A2 => n7343, B1 => 
                           REGISTERS_19_10_port, B2 => n7375, ZN => n7120);
   U2594 : NAND4_X1 port map( A1 => n7123, A2 => n7122, A3 => n7121, A4 => 
                           n7120, ZN => n7129);
   U2595 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n7285, B1 => 
                           REGISTERS_21_10_port, B2 => n7370, ZN => n7127);
   U2596 : AOI22_X1 port map( A1 => REGISTERS_18_10_port, A2 => n7381, B1 => 
                           REGISTERS_23_10_port, B2 => n7384, ZN => n7126);
   U2597 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n7337, B1 => 
                           REGISTERS_27_10_port, B2 => n7369, ZN => n7125);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n7368, B1 => 
                           REGISTERS_29_10_port, B2 => n7315, ZN => n7124);
   U2599 : NAND4_X1 port map( A1 => n7127, A2 => n7126, A3 => n7125, A4 => 
                           n7124, ZN => n7128);
   U2600 : NOR2_X1 port map( A1 => n7129, A2 => n7128, ZN => n7141);
   U2601 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n7407, B1 => 
                           REGISTERS_5_10_port, B2 => n7394, ZN => n7133);
   U2602 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n7397, B1 => 
                           REGISTERS_6_10_port, B2 => n7411, ZN => n7132);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n7251, B1 => 
                           REGISTERS_1_10_port, B2 => n7395, ZN => n7131);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_2_10_port, A2 => n7405, B1 => 
                           REGISTERS_3_10_port, B2 => n7408, ZN => n7130);
   U2605 : NAND4_X1 port map( A1 => n7133, A2 => n7132, A3 => n7131, A4 => 
                           n7130, ZN => n7139);
   U2606 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n7357, B1 => 
                           REGISTERS_14_10_port, B2 => n7399, ZN => n7137);
   U2607 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n7400, B1 => 
                           REGISTERS_9_10_port, B2 => n7356, ZN => n7136);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n7394, B1 => 
                           REGISTERS_8_10_port, B2 => n7351, ZN => n7135);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n7410, B1 => 
                           REGISTERS_10_10_port, B2 => n7358, ZN => n7134);
   U2610 : NAND4_X1 port map( A1 => n7137, A2 => n7136, A3 => n7135, A4 => 
                           n7134, ZN => n7138);
   U2611 : AOI22_X1 port map( A1 => n7259, A2 => n7139, B1 => n7257, B2 => 
                           n7138, ZN => n7140);
   U2612 : OAI21_X1 port map( B1 => n7423, B2 => n7141, A => n7140, ZN => N395)
                           ;
   U2613 : AOI22_X1 port map( A1 => REGISTERS_27_9_port, A2 => n7142, B1 => 
                           REGISTERS_22_9_port, B2 => n7382, ZN => n7146);
   U2614 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n7335, B1 => 
                           REGISTERS_24_9_port, B2 => n7387, ZN => n7145);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n7374, B1 => 
                           REGISTERS_29_9_port, B2 => n7315, ZN => n7144);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_26_9_port, A2 => n7343, B1 => 
                           REGISTERS_31_9_port, B2 => n7373, ZN => n7143);
   U2617 : NAND4_X1 port map( A1 => n7146, A2 => n7145, A3 => n7144, A4 => 
                           n7143, ZN => n7152);
   U2618 : AOI22_X1 port map( A1 => REGISTERS_19_9_port, A2 => n7375, B1 => 
                           REGISTERS_20_9_port, B2 => n7314, ZN => n7150);
   U2619 : AOI22_X1 port map( A1 => REGISTERS_18_9_port, A2 => n7188, B1 => 
                           REGISTERS_16_9_port, B2 => n7386, ZN => n7149);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_30_9_port, A2 => n7385, B1 => 
                           REGISTERS_28_9_port, B2 => n7368, ZN => n7148);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n7370, B1 => 
                           REGISTERS_23_9_port, B2 => n7384, ZN => n7147);
   U2622 : NAND4_X1 port map( A1 => n7150, A2 => n7149, A3 => n7148, A4 => 
                           n7147, ZN => n7151);
   U2623 : NOR2_X1 port map( A1 => n7152, A2 => n7151, ZN => n7164);
   U2624 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n7357, B1 => 
                           REGISTERS_0_9_port, B2 => n7406, ZN => n7156);
   U2625 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n7227, B1 => 
                           REGISTERS_2_9_port, B2 => n7398, ZN => n7155);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n7400, B1 => 
                           REGISTERS_4_9_port, B2 => n7396, ZN => n7154);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n7356, B1 => 
                           REGISTERS_6_9_port, B2 => n7399, ZN => n7153);
   U2628 : NAND4_X1 port map( A1 => n7156, A2 => n7155, A3 => n7154, A4 => 
                           n7153, ZN => n7162);
   U2629 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n7397, B1 => 
                           REGISTERS_11_9_port, B2 => n7408, ZN => n7160);
   U2630 : AOI22_X1 port map( A1 => REGISTERS_10_9_port, A2 => n7398, B1 => 
                           REGISTERS_12_9_port, B2 => n7396, ZN => n7159);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_14_9_port, A2 => n7399, B1 => 
                           REGISTERS_15_9_port, B2 => n7296, ZN => n7158);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n7227, B1 => 
                           REGISTERS_9_9_port, B2 => n7409, ZN => n7157);
   U2633 : NAND4_X1 port map( A1 => n7160, A2 => n7159, A3 => n7158, A4 => 
                           n7157, ZN => n7161);
   U2634 : AOI22_X1 port map( A1 => n7259, A2 => n7162, B1 => n7257, B2 => 
                           n7161, ZN => n7163);
   U2635 : OAI21_X1 port map( B1 => n7367, B2 => n7164, A => n7163, ZN => N394)
                           ;
   U2636 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n7165, B1 => 
                           REGISTERS_26_8_port, B2 => n7372, ZN => n7169);
   U2637 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n7337, B1 => 
                           REGISTERS_18_8_port, B2 => n7381, ZN => n7168);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n7369, B1 => 
                           REGISTERS_30_8_port, B2 => n7309, ZN => n7167);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n7368, B1 => 
                           REGISTERS_16_8_port, B2 => n7386, ZN => n7166);
   U2640 : NAND4_X1 port map( A1 => n7169, A2 => n7168, A3 => n7167, A4 => 
                           n7166, ZN => n7175);
   U2641 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n7315, B1 => 
                           REGISTERS_25_8_port, B2 => n7374, ZN => n7173);
   U2642 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n7375, B1 => 
                           REGISTERS_17_8_port, B2 => n7335, ZN => n7172);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_31_8_port, A2 => n7373, B1 => 
                           REGISTERS_22_8_port, B2 => n7382, ZN => n7171);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n7371, B1 => 
                           REGISTERS_23_8_port, B2 => n7384, ZN => n7170);
   U2645 : NAND4_X1 port map( A1 => n7173, A2 => n7172, A3 => n7171, A4 => 
                           n7170, ZN => n7174);
   U2646 : NOR2_X1 port map( A1 => n7175, A2 => n7174, ZN => n7187);
   U2647 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n7410, B1 => 
                           REGISTERS_5_8_port, B2 => n7412, ZN => n7179);
   U2648 : AOI22_X1 port map( A1 => REGISTERS_3_8_port, A2 => n7350, B1 => 
                           REGISTERS_1_8_port, B2 => n7356, ZN => n7178);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n7397, B1 => 
                           REGISTERS_2_8_port, B2 => n7358, ZN => n7177);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n7400, B1 => 
                           REGISTERS_6_8_port, B2 => n7322, ZN => n7176);
   U2651 : NAND4_X1 port map( A1 => n7179, A2 => n7178, A3 => n7177, A4 => 
                           n7176, ZN => n7185);
   U2652 : AOI22_X1 port map( A1 => REGISTERS_10_8_port, A2 => n7358, B1 => 
                           REGISTERS_9_8_port, B2 => n7409, ZN => n7183);
   U2653 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n7394, B1 => 
                           REGISTERS_12_8_port, B2 => n7396, ZN => n7182);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n7397, B1 => 
                           REGISTERS_11_8_port, B2 => n7350, ZN => n7181);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_14_8_port, A2 => n7399, B1 => 
                           REGISTERS_15_8_port, B2 => n7407, ZN => n7180);
   U2656 : NAND4_X1 port map( A1 => n7183, A2 => n7182, A3 => n7181, A4 => 
                           n7180, ZN => n7184);
   U2657 : AOI22_X1 port map( A1 => n7259, A2 => n7185, B1 => n7257, B2 => 
                           n7184, ZN => n7186);
   U2658 : OAI21_X1 port map( B1 => n7423, B2 => n7187, A => n7186, ZN => N393)
                           ;
   U2659 : AOI22_X1 port map( A1 => REGISTERS_18_7_port, A2 => n7188, B1 => 
                           REGISTERS_17_7_port, B2 => n7335, ZN => n7192);
   U2660 : AOI22_X1 port map( A1 => REGISTERS_31_7_port, A2 => n7373, B1 => 
                           REGISTERS_19_7_port, B2 => n7336, ZN => n7191);
   U2661 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n7315, B1 => 
                           REGISTERS_25_7_port, B2 => n7374, ZN => n7190);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n7370, B1 => 
                           REGISTERS_28_7_port, B2 => n7368, ZN => n7189);
   U2663 : NAND4_X1 port map( A1 => n7192, A2 => n7191, A3 => n7190, A4 => 
                           n7189, ZN => n7198);
   U2664 : AOI22_X1 port map( A1 => REGISTERS_30_7_port, A2 => n7385, B1 => 
                           REGISTERS_20_7_port, B2 => n7314, ZN => n7196);
   U2665 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n7337, B1 => 
                           REGISTERS_27_7_port, B2 => n7369, ZN => n7195);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n7285, B1 => 
                           REGISTERS_26_7_port, B2 => n7372, ZN => n7194);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n7382, B1 => 
                           REGISTERS_23_7_port, B2 => n7384, ZN => n7193);
   U2668 : NAND4_X1 port map( A1 => n7196, A2 => n7195, A3 => n7194, A4 => 
                           n7193, ZN => n7197);
   U2669 : NOR2_X1 port map( A1 => n7198, A2 => n7197, ZN => n7210);
   U2670 : AOI22_X1 port map( A1 => REGISTERS_6_7_port, A2 => n7322, B1 => 
                           REGISTERS_2_7_port, B2 => n7398, ZN => n7202);
   U2671 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n7357, B1 => 
                           REGISTERS_7_7_port, B2 => n7407, ZN => n7201);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n7412, B1 => 
                           REGISTERS_0_7_port, B2 => n7351, ZN => n7200);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n7395, B1 => 
                           REGISTERS_4_7_port, B2 => n7251, ZN => n7199);
   U2674 : NAND4_X1 port map( A1 => n7202, A2 => n7201, A3 => n7200, A4 => 
                           n7199, ZN => n7208);
   U2675 : AOI22_X1 port map( A1 => REGISTERS_15_7_port, A2 => n7400, B1 => 
                           REGISTERS_8_7_port, B2 => n7351, ZN => n7206);
   U2676 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n7227, B1 => 
                           REGISTERS_12_7_port, B2 => n7410, ZN => n7205);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_10_7_port, A2 => n7398, B1 => 
                           REGISTERS_14_7_port, B2 => n7322, ZN => n7204);
   U2678 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n7357, B1 => 
                           REGISTERS_9_7_port, B2 => n7409, ZN => n7203);
   U2679 : NAND4_X1 port map( A1 => n7206, A2 => n7205, A3 => n7204, A4 => 
                           n7203, ZN => n7207);
   U2680 : AOI22_X1 port map( A1 => n7259, A2 => n7208, B1 => n7257, B2 => 
                           n7207, ZN => n7209);
   U2681 : OAI21_X1 port map( B1 => n7367, B2 => n7210, A => n7209, ZN => N392)
                           ;
   U2682 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n7285, B1 => 
                           REGISTERS_29_6_port, B2 => n7380, ZN => n7214);
   U2683 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n7368, B1 => 
                           REGISTERS_27_6_port, B2 => n7369, ZN => n7213);
   U2684 : AOI22_X1 port map( A1 => REGISTERS_22_6_port, A2 => n7266, B1 => 
                           REGISTERS_24_6_port, B2 => n7387, ZN => n7212);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n7371, B1 => 
                           REGISTERS_26_6_port, B2 => n7372, ZN => n7211);
   U2686 : NAND4_X1 port map( A1 => n7214, A2 => n7213, A3 => n7212, A4 => 
                           n7211, ZN => n7222);
   U2687 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n7215, B1 => 
                           REGISTERS_30_6_port, B2 => n7309, ZN => n7220);
   U2688 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n7335, B1 => 
                           REGISTERS_31_6_port, B2 => n7338, ZN => n7219);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n7216, B1 => 
                           REGISTERS_19_6_port, B2 => n7336, ZN => n7218);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n7370, B1 => 
                           REGISTERS_18_6_port, B2 => n7381, ZN => n7217);
   U2691 : NAND4_X1 port map( A1 => n7220, A2 => n7219, A3 => n7218, A4 => 
                           n7217, ZN => n7221);
   U2692 : NOR2_X1 port map( A1 => n7222, A2 => n7221, ZN => n7236);
   U2693 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n7400, B1 => 
                           REGISTERS_6_6_port, B2 => n7411, ZN => n7226);
   U2694 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n7356, B1 => 
                           REGISTERS_3_6_port, B2 => n7357, ZN => n7225);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_2_6_port, A2 => n7405, B1 => 
                           REGISTERS_0_6_port, B2 => n7406, ZN => n7224);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n7396, B1 => 
                           REGISTERS_5_6_port, B2 => n7412, ZN => n7223);
   U2697 : NAND4_X1 port map( A1 => n7226, A2 => n7225, A3 => n7224, A4 => 
                           n7223, ZN => n7233);
   U2698 : AOI22_X1 port map( A1 => REGISTERS_10_6_port, A2 => n7398, B1 => 
                           REGISTERS_8_6_port, B2 => n7406, ZN => n7231);
   U2699 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n7356, B1 => 
                           REGISTERS_15_6_port, B2 => n7296, ZN => n7230);
   U2700 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n7410, B1 => 
                           REGISTERS_13_6_port, B2 => n7227, ZN => n7229);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_14_6_port, A2 => n7411, B1 => 
                           REGISTERS_11_6_port, B2 => n7357, ZN => n7228);
   U2702 : NAND4_X1 port map( A1 => n7231, A2 => n7230, A3 => n7229, A4 => 
                           n7228, ZN => n7232);
   U2703 : AOI22_X1 port map( A1 => n7234, A2 => n7233, B1 => n7257, B2 => 
                           n7232, ZN => n7235);
   U2704 : OAI21_X1 port map( B1 => n7423, B2 => n7236, A => n7235, ZN => N391)
                           ;
   U2705 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n7371, B1 => 
                           REGISTERS_18_5_port, B2 => n7381, ZN => n7240);
   U2706 : AOI22_X1 port map( A1 => REGISTERS_26_5_port, A2 => n7343, B1 => 
                           REGISTERS_31_5_port, B2 => n7338, ZN => n7239);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n7370, B1 => 
                           REGISTERS_16_5_port, B2 => n7386, ZN => n7238);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n7384, B1 => 
                           REGISTERS_24_5_port, B2 => n7387, ZN => n7237);
   U2709 : NAND4_X1 port map( A1 => n7240, A2 => n7239, A3 => n7238, A4 => 
                           n7237, ZN => n7246);
   U2710 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n7368, B1 => 
                           REGISTERS_17_5_port, B2 => n7335, ZN => n7244);
   U2711 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n7369, B1 => 
                           REGISTERS_30_5_port, B2 => n7309, ZN => n7243);
   U2712 : AOI22_X1 port map( A1 => REGISTERS_22_5_port, A2 => n7382, B1 => 
                           REGISTERS_29_5_port, B2 => n7380, ZN => n7242);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n7374, B1 => 
                           REGISTERS_19_5_port, B2 => n7336, ZN => n7241);
   U2714 : NAND4_X1 port map( A1 => n7244, A2 => n7243, A3 => n7242, A4 => 
                           n7241, ZN => n7245);
   U2715 : NOR2_X1 port map( A1 => n7246, A2 => n7245, ZN => n7261);
   U2716 : AOI22_X1 port map( A1 => REGISTERS_6_5_port, A2 => n7322, B1 => 
                           REGISTERS_5_5_port, B2 => n7394, ZN => n7250);
   U2717 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n7400, B1 => 
                           REGISTERS_3_5_port, B2 => n7408, ZN => n7249);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n7395, B1 => 
                           REGISTERS_0_5_port, B2 => n7406, ZN => n7248);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n7251, B1 => 
                           REGISTERS_2_5_port, B2 => n7358, ZN => n7247);
   U2720 : NAND4_X1 port map( A1 => n7250, A2 => n7249, A3 => n7248, A4 => 
                           n7247, ZN => n7258);
   U2721 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n7397, B1 => 
                           REGISTERS_9_5_port, B2 => n7395, ZN => n7255);
   U2722 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n7350, B1 => 
                           REGISTERS_12_5_port, B2 => n7251, ZN => n7254);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n7400, B1 => 
                           REGISTERS_13_5_port, B2 => n7394, ZN => n7253);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_14_5_port, A2 => n7322, B1 => 
                           REGISTERS_10_5_port, B2 => n7398, ZN => n7252);
   U2725 : NAND4_X1 port map( A1 => n7255, A2 => n7254, A3 => n7253, A4 => 
                           n7252, ZN => n7256);
   U2726 : AOI22_X1 port map( A1 => n7259, A2 => n7258, B1 => n7257, B2 => 
                           n7256, ZN => n7260);
   U2727 : OAI21_X1 port map( B1 => n7367, B2 => n7261, A => n7260, ZN => N390)
                           ;
   U2728 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n7371, B1 => 
                           REGISTERS_23_4_port, B2 => n7384, ZN => n7265);
   U2729 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n7375, B1 => 
                           REGISTERS_18_4_port, B2 => n7381, ZN => n7264);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n7369, B1 => 
                           REGISTERS_17_4_port, B2 => n7335, ZN => n7263);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n7285, B1 => 
                           REGISTERS_25_4_port, B2 => n7374, ZN => n7262);
   U2732 : NAND4_X1 port map( A1 => n7265, A2 => n7264, A3 => n7263, A4 => 
                           n7262, ZN => n7272);
   U2733 : AOI22_X1 port map( A1 => REGISTERS_30_4_port, A2 => n7309, B1 => 
                           REGISTERS_21_4_port, B2 => n7370, ZN => n7270);
   U2734 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n7266, B1 => 
                           REGISTERS_26_4_port, B2 => n7372, ZN => n7269);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n7337, B1 => 
                           REGISTERS_31_4_port, B2 => n7338, ZN => n7268);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n7368, B1 => 
                           REGISTERS_29_4_port, B2 => n7380, ZN => n7267);
   U2737 : NAND4_X1 port map( A1 => n7270, A2 => n7269, A3 => n7268, A4 => 
                           n7267, ZN => n7271);
   U2738 : NOR2_X1 port map( A1 => n7272, A2 => n7271, ZN => n7284);
   U2739 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n7409, B1 => 
                           REGISTERS_3_4_port, B2 => n7350, ZN => n7276);
   U2740 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n7412, B1 => 
                           REGISTERS_4_4_port, B2 => n7410, ZN => n7275);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_6_4_port, A2 => n7411, B1 => 
                           REGISTERS_7_4_port, B2 => n7407, ZN => n7274);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_2_4_port, A2 => n7405, B1 => 
                           REGISTERS_0_4_port, B2 => n7351, ZN => n7273);
   U2743 : NAND4_X1 port map( A1 => n7276, A2 => n7275, A3 => n7274, A4 => 
                           n7273, ZN => n7282);
   U2744 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n7410, B1 => 
                           REGISTERS_14_4_port, B2 => n7322, ZN => n7280);
   U2745 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n7400, B1 => 
                           REGISTERS_11_4_port, B2 => n7357, ZN => n7279);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n7394, B1 => 
                           REGISTERS_9_4_port, B2 => n7395, ZN => n7278);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_10_4_port, A2 => n7358, B1 => 
                           REGISTERS_8_4_port, B2 => n7351, ZN => n7277);
   U2748 : NAND4_X1 port map( A1 => n7280, A2 => n7279, A3 => n7278, A4 => 
                           n7277, ZN => n7281);
   U2749 : AOI22_X1 port map( A1 => n7420, A2 => n7282, B1 => n7418, B2 => 
                           n7281, ZN => n7283);
   U2750 : OAI21_X1 port map( B1 => n7423, B2 => n7284, A => n7283, ZN => N389)
                           ;
   U2751 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n7315, B1 => 
                           REGISTERS_31_3_port, B2 => n7338, ZN => n7289);
   U2752 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n7285, B1 => 
                           REGISTERS_25_3_port, B2 => n7374, ZN => n7288);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n7368, B1 => 
                           REGISTERS_18_3_port, B2 => n7381, ZN => n7287);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n7375, B1 => 
                           REGISTERS_23_3_port, B2 => n7384, ZN => n7286);
   U2755 : NAND4_X1 port map( A1 => n7289, A2 => n7288, A3 => n7287, A4 => 
                           n7286, ZN => n7295);
   U2756 : AOI22_X1 port map( A1 => REGISTERS_26_3_port, A2 => n7343, B1 => 
                           REGISTERS_17_3_port, B2 => n7335, ZN => n7293);
   U2757 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n7371, B1 => 
                           REGISTERS_24_3_port, B2 => n7387, ZN => n7292);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_27_3_port, A2 => n7369, B1 => 
                           REGISTERS_22_3_port, B2 => n7382, ZN => n7291);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n7370, B1 => 
                           REGISTERS_30_3_port, B2 => n7309, ZN => n7290);
   U2760 : NAND4_X1 port map( A1 => n7293, A2 => n7292, A3 => n7291, A4 => 
                           n7290, ZN => n7294);
   U2761 : NOR2_X1 port map( A1 => n7295, A2 => n7294, ZN => n7308);
   U2762 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n7395, B1 => 
                           REGISTERS_4_3_port, B2 => n7410, ZN => n7300);
   U2763 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n7412, B1 => 
                           REGISTERS_3_3_port, B2 => n7357, ZN => n7299);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_6_3_port, A2 => n7411, B1 => 
                           REGISTERS_0_3_port, B2 => n7406, ZN => n7298);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n7405, B1 => 
                           REGISTERS_7_3_port, B2 => n7296, ZN => n7297);
   U2766 : NAND4_X1 port map( A1 => n7300, A2 => n7299, A3 => n7298, A4 => 
                           n7297, ZN => n7306);
   U2767 : AOI22_X1 port map( A1 => REGISTERS_10_3_port, A2 => n7358, B1 => 
                           REGISTERS_14_3_port, B2 => n7399, ZN => n7304);
   U2768 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n7397, B1 => 
                           REGISTERS_12_3_port, B2 => n7396, ZN => n7303);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n7412, B1 => 
                           REGISTERS_11_3_port, B2 => n7350, ZN => n7302);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n7356, B1 => 
                           REGISTERS_15_3_port, B2 => n7407, ZN => n7301);
   U2771 : NAND4_X1 port map( A1 => n7304, A2 => n7303, A3 => n7302, A4 => 
                           n7301, ZN => n7305);
   U2772 : AOI22_X1 port map( A1 => n7420, A2 => n7306, B1 => n7418, B2 => 
                           n7305, ZN => n7307);
   U2773 : OAI21_X1 port map( B1 => n7367, B2 => n7308, A => n7307, ZN => N388)
                           ;
   U2774 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n7373, B1 => 
                           REGISTERS_17_2_port, B2 => n7335, ZN => n7313);
   U2775 : AOI22_X1 port map( A1 => REGISTERS_26_2_port, A2 => n7343, B1 => 
                           REGISTERS_25_2_port, B2 => n7374, ZN => n7312);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n7337, B1 => 
                           REGISTERS_16_2_port, B2 => n7386, ZN => n7311);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_19_2_port, A2 => n7375, B1 => 
                           REGISTERS_30_2_port, B2 => n7309, ZN => n7310);
   U2778 : NAND4_X1 port map( A1 => n7313, A2 => n7312, A3 => n7311, A4 => 
                           n7310, ZN => n7321);
   U2779 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n7315, B1 => 
                           REGISTERS_20_2_port, B2 => n7314, ZN => n7319);
   U2780 : AOI22_X1 port map( A1 => REGISTERS_18_2_port, A2 => n7381, B1 => 
                           REGISTERS_21_2_port, B2 => n7370, ZN => n7318);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_22_2_port, A2 => n7382, B1 => 
                           REGISTERS_23_2_port, B2 => n7384, ZN => n7317);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n7369, B1 => 
                           REGISTERS_28_2_port, B2 => n7368, ZN => n7316);
   U2783 : NAND4_X1 port map( A1 => n7319, A2 => n7318, A3 => n7317, A4 => 
                           n7316, ZN => n7320);
   U2784 : NOR2_X1 port map( A1 => n7321, A2 => n7320, ZN => n7334);
   U2785 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n7410, B1 => 
                           REGISTERS_1_2_port, B2 => n7409, ZN => n7326);
   U2786 : AOI22_X1 port map( A1 => REGISTERS_2_2_port, A2 => n7398, B1 => 
                           REGISTERS_0_2_port, B2 => n7406, ZN => n7325);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n7400, B1 => 
                           REGISTERS_6_2_port, B2 => n7322, ZN => n7324);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n7412, B1 => 
                           REGISTERS_3_2_port, B2 => n7408, ZN => n7323);
   U2789 : NAND4_X1 port map( A1 => n7326, A2 => n7325, A3 => n7324, A4 => 
                           n7323, ZN => n7332);
   U2790 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n7410, B1 => 
                           REGISTERS_11_2_port, B2 => n7350, ZN => n7330);
   U2791 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n7400, B1 => 
                           REGISTERS_9_2_port, B2 => n7395, ZN => n7329);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_14_2_port, A2 => n7411, B1 => 
                           REGISTERS_10_2_port, B2 => n7358, ZN => n7328);
   U2793 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n7412, B1 => 
                           REGISTERS_8_2_port, B2 => n7351, ZN => n7327);
   U2794 : NAND4_X1 port map( A1 => n7330, A2 => n7329, A3 => n7328, A4 => 
                           n7327, ZN => n7331);
   U2795 : AOI22_X1 port map( A1 => n7420, A2 => n7332, B1 => n7418, B2 => 
                           n7331, ZN => n7333);
   U2796 : OAI21_X1 port map( B1 => n7423, B2 => n7334, A => n7333, ZN => N387)
                           ;
   U2797 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n7381, B1 => 
                           REGISTERS_17_1_port, B2 => n7335, ZN => n7342);
   U2798 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n7337, B1 => 
                           REGISTERS_19_1_port, B2 => n7336, ZN => n7341);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n7371, B1 => 
                           REGISTERS_31_1_port, B2 => n7338, ZN => n7340);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n7370, B1 => 
                           REGISTERS_29_1_port, B2 => n7380, ZN => n7339);
   U2801 : NAND4_X1 port map( A1 => n7342, A2 => n7341, A3 => n7340, A4 => 
                           n7339, ZN => n7349);
   U2802 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n7368, B1 => 
                           REGISTERS_25_1_port, B2 => n7374, ZN => n7347);
   U2803 : AOI22_X1 port map( A1 => REGISTERS_30_1_port, A2 => n7385, B1 => 
                           REGISTERS_22_1_port, B2 => n7382, ZN => n7346);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_23_1_port, A2 => n7384, B1 => 
                           REGISTERS_27_1_port, B2 => n7369, ZN => n7345);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_26_1_port, A2 => n7343, B1 => 
                           REGISTERS_16_1_port, B2 => n7386, ZN => n7344);
   U2806 : NAND4_X1 port map( A1 => n7347, A2 => n7346, A3 => n7345, A4 => 
                           n7344, ZN => n7348);
   U2807 : NOR2_X1 port map( A1 => n7349, A2 => n7348, ZN => n7366);
   U2808 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n7395, B1 => 
                           REGISTERS_3_1_port, B2 => n7350, ZN => n7355);
   U2809 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n7410, B1 => 
                           REGISTERS_2_1_port, B2 => n7405, ZN => n7354);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n7400, B1 => 
                           REGISTERS_0_1_port, B2 => n7351, ZN => n7353);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n7411, B1 => 
                           REGISTERS_5_1_port, B2 => n7412, ZN => n7352);
   U2812 : NAND4_X1 port map( A1 => n7355, A2 => n7354, A3 => n7353, A4 => 
                           n7352, ZN => n7364);
   U2813 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n7410, B1 => 
                           REGISTERS_9_1_port, B2 => n7356, ZN => n7362);
   U2814 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n7397, B1 => 
                           REGISTERS_13_1_port, B2 => n7394, ZN => n7361);
   U2815 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n7357, B1 => 
                           REGISTERS_15_1_port, B2 => n7407, ZN => n7360);
   U2816 : AOI22_X1 port map( A1 => REGISTERS_14_1_port, A2 => n7411, B1 => 
                           REGISTERS_10_1_port, B2 => n7358, ZN => n7359);
   U2817 : NAND4_X1 port map( A1 => n7362, A2 => n7361, A3 => n7360, A4 => 
                           n7359, ZN => n7363);
   U2818 : AOI22_X1 port map( A1 => n7420, A2 => n7364, B1 => n7418, B2 => 
                           n7363, ZN => n7365);
   U2819 : OAI21_X1 port map( B1 => n7367, B2 => n7366, A => n7365, ZN => N386)
                           ;
   U2820 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n7369, B1 => 
                           REGISTERS_28_0_port, B2 => n7368, ZN => n7379);
   U2821 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n7371, B1 => 
                           REGISTERS_21_0_port, B2 => n7370, ZN => n7378);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_31_0_port, A2 => n7373, B1 => 
                           REGISTERS_26_0_port, B2 => n7372, ZN => n7377);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_19_0_port, A2 => n7375, B1 => 
                           REGISTERS_25_0_port, B2 => n7374, ZN => n7376);
   U2824 : NAND4_X1 port map( A1 => n7379, A2 => n7378, A3 => n7377, A4 => 
                           n7376, ZN => n7393);
   U2825 : AOI22_X1 port map( A1 => REGISTERS_18_0_port, A2 => n7381, B1 => 
                           REGISTERS_29_0_port, B2 => n7380, ZN => n7391);
   U2826 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n7383, B1 => 
                           REGISTERS_22_0_port, B2 => n7382, ZN => n7390);
   U2827 : AOI22_X1 port map( A1 => REGISTERS_30_0_port, A2 => n7385, B1 => 
                           REGISTERS_23_0_port, B2 => n7384, ZN => n7389);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n7387, B1 => 
                           REGISTERS_16_0_port, B2 => n7386, ZN => n7388);
   U2829 : NAND4_X1 port map( A1 => n7391, A2 => n7390, A3 => n7389, A4 => 
                           n7388, ZN => n7392);
   U2830 : NOR2_X1 port map( A1 => n7393, A2 => n7392, ZN => n7422);
   U2831 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n7395, B1 => 
                           REGISTERS_5_0_port, B2 => n7394, ZN => n7404);
   U2832 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n7397, B1 => 
                           REGISTERS_4_0_port, B2 => n7396, ZN => n7403);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n7398, B1 => 
                           REGISTERS_3_0_port, B2 => n7408, ZN => n7402);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n7400, B1 => 
                           REGISTERS_6_0_port, B2 => n7399, ZN => n7401);
   U2835 : NAND4_X1 port map( A1 => n7404, A2 => n7403, A3 => n7402, A4 => 
                           n7401, ZN => n7419);
   U2836 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n7406, B1 => 
                           REGISTERS_10_0_port, B2 => n7405, ZN => n7416);
   U2837 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n7408, B1 => 
                           REGISTERS_15_0_port, B2 => n7407, ZN => n7415);
   U2838 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n7410, B1 => 
                           REGISTERS_9_0_port, B2 => n7409, ZN => n7414);
   U2839 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n7412, B1 => 
                           REGISTERS_14_0_port, B2 => n7411, ZN => n7413);
   U2840 : NAND4_X1 port map( A1 => n7416, A2 => n7415, A3 => n7414, A4 => 
                           n7413, ZN => n7417);
   U2841 : AOI22_X1 port map( A1 => n7420, A2 => n7419, B1 => n7418, B2 => 
                           n7417, ZN => n7421);
   U2842 : OAI21_X1 port map( B1 => n7423, B2 => n7422, A => n7421, ZN => N385)
                           ;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ENABLE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_28_port, 
      curr_instruction_to_cu_i_27_port, curr_instruction_to_cu_i_26_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_5_port, curr_instruction_to_cu_i_4_port, 
      curr_instruction_to_cu_i_3_port, curr_instruction_to_cu_i_2_port, 
      curr_instruction_to_cu_i_1_port, curr_instruction_to_cu_i_0_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n131, cu_i_n127, 
      cu_i_n126, cu_i_n125, cu_i_n124, cu_i_n123, cu_i_n210, cu_i_n209, 
      cu_i_n145, cu_i_n26, cu_i_n25, cu_i_n23, cu_i_cw1_i_4_port, 
      cu_i_cw1_i_7_port, cu_i_cw1_i_8_port, cu_i_cw3_6_port, cu_i_cw2_5_port, 
      cu_i_cw2_6_port, cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_0_port, 
      cu_i_cw1_1_port, cu_i_cw1_2_port, cu_i_cw1_3_port, cu_i_cw1_4_port, 
      cu_i_cw1_5_port, cu_i_cw1_6_port, cu_i_cw1_7_port, cu_i_cw1_8_port, 
      cu_i_cw1_10_port, cu_i_cw1_11_port, cu_i_cw1_12_port, cu_i_cw1_13_port, 
      cu_i_N279, cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, 
      cu_i_N273, cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, 
      cu_i_cmd_alu_op_type_0_port, cu_i_cmd_alu_op_type_1_port, 
      cu_i_cmd_alu_op_type_2_port, cu_i_cmd_alu_op_type_3_port, 
      cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, cu_i_cmd_word_4_port, 
      cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, cu_i_cmd_word_8_port, 
      cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n78, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_n12, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_decode_stage_dp_enable_sign_extension_logic, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n309, n310, n311, n691, n697,
      n699, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n737, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n756, n758, n759, n760, n761, n762, n763, n764, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1155, n1156, n1157, n1158, n1159, n1160, n1161, 
      n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, 
      n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, 
      n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, 
      n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, 
      n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, 
      n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, 
      n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
      n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, 
      n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
      n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, 
      n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, 
      n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, 
      n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, 
      n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
      n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, 
      n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, 
      n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
      n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, 
      n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, 
      n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, 
      n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, 
      n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
      n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, 
      n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, 
      n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, 
      n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, 
      n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
      n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
      n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, 
      n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1546, DRAM_ENABLE_port, n1548, n1549, n_1413
      , n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422,
      n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, 
      n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, 
      n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, 
      n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, 
      n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, 
      n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, 
      n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, 
      n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, 
      n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, 
      n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, 
      n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, 
      n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, 
      n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, 
      n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, 
      n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, 
      n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, 
      n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, 
      n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, 
      n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, 
      n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, 
      n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, 
      n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, 
      n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, 
      n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, 
      n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, 
      n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, 
      n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, 
      n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, 
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, 
      n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, 
      n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, 
      n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, 
      n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, 
      n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, 
      n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, 
      n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, 
      n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, 
      n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, 
      n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => n1542, QN => cu_i_n25);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => n1539, QN => cu_i_n124);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => n1532, QN => cu_i_n125);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => n_1413, QN => cu_i_n123);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n12, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n43, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1414, mul_exeception => 
                           n_1415, FUNC(0) => n1147, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1416, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n1546, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n309, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n1546, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n309, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n1546, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n309, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n1546, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n309, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n1546, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n309, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n309, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n309, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n1546, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n1546, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n1546, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n1546, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n1546, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n1546, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n1546, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n1546, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n1546, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n1546, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n309, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n309, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n1546, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n1546, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n1546, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n1546, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n1546, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n1546, Z 
                           => DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n1548, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n1548, Z =>
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n1548, Z =>
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n1548, Z =>
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n1548, Z =>
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n1548, Z =>
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n1548, Z =>
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n1548, Z =>
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n1548, Z =>
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n1548, Z =>
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n1548, Z =>
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n1548, Z =>
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => n1548, Z =>
                           DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => n1548, Z =>
                           DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => n1548, Z =>
                           DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => n1548, Z =>
                           DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => n1548, Z =>
                           DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1417);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n1545, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n1545, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n1545, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n310, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n1545, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n1545, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n310, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n18, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n1549, D => datapath_i_n17, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n1549, D => datapath_i_n16, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n15, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n1549, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n1549, D => 
                           curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n1549, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n12, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n11, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n1549, D => datapath_i_n10, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n1549, D => datapath_i_n9, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n1155, CK => CLK, RN => RST
                           , Q => cu_i_cw3_6_port, QN => n_1418);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n131, CK => CLK, RN =>
                           RST, Q => n_1419, QN => n699);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1420);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1421);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1422);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n126, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n1544);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => n_1423, QN => n756);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n310, CK => CLK, RN => RST,
                           Q => cu_i_cw1_13_port, QN => n_1424);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1425)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1426)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1427)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1428);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1429);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n311, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1430);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1431);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => n1152, CK => CLK, RN => RST,
                           Q => cu_i_cw1_4_port, QN => n_1432);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1433);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1434);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1435);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1436);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1437);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1438);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1439);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1440);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1441);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1442);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1443);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1444);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1445);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1446);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1447);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1448);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1449);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1450);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1451);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1452);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1453);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1454);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1455);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1456);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1457);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1458);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1459);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1460);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1461);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1462);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1463);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1464);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1465);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1466);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1467);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1468)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1469)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1470)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1471)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1472)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1473)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1474)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1475)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1476)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1477)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1478)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1479)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1480)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1481)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1482)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1483)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1484)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1485)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1486)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1487)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1488)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1489)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1490);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1491);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1492);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1493);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1494);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1495);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1496);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1497);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1498);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1499);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1500);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1501);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1502);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1503);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1504);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1505);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1506);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1507);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1508);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1509);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1510);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1511);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1512);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1513);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1514);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1515);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1516);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1517);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1518);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1519);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1520);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1521);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1522);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1523);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1524);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1525);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1526);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1527);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1528);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1529);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1530);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1531);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1532);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1533);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1534);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1535);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1536);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1537);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1538);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1539);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1540);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1541);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1542);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1543);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1544);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1545);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1546);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1547);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1548);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1549);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1550);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1551);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1552);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1553);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1554);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1555);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1556);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1557);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1558);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1559);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1560);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1561);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1562);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1563);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1564, QN => n703);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1565, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1566, QN => n726);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1567, QN => n725);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1568, QN => n724);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1569, QN => n691);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1570, QN => n723);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1571, QN => n722);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1572, QN => n721);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1573, QN => n720);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1574, QN => n719);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1575, QN => n718);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1576, QN => n717);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1577, QN => n716);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1578, QN => n715);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1579, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1580, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1581, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1582, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1583, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1584, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1585, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1586, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1587, QN => n706);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1588, QN => n705);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1589, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1590, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1591, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1592, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1593, QN => n728);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1594, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1595, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1596);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1597);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1598);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1599);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1600);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1601);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1602);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1603);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1604);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1605);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1606);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1607);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1608);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1609);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1610);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1611);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1612);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1613);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1614);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1615);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1616);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1617);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1618);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1619);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1620);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1621);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1622);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1623);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1624);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1625);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1626);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1627);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1628);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1629);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1630);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1631);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1632);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1633);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1634);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1635);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1636);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1637);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1638);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1639);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1640);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1641);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1642);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1643);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1644);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1645);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1646);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1647);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1648);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1649);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1650);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1651);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1652);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1653);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1654);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n764);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n763);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n762);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n761);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n760);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n759);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n758);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1655);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1656);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1657);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1658);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1659);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1660);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1661);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1662);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1663);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1664);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1665);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1666);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1667);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1668);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1669);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1670);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1671);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1672);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1673);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1674);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1675);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1676);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1677);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1678);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1679);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1680);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1681);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1682);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1683);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1684);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1685);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1686);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1687);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1688);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1689);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1690);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1691);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1692);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1693);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1694);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1695);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1696);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1697);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1698);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1699);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1700);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1701);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1702);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1703);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1704);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1705);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1706);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1707);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1708);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1709);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1710);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1711);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1712);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1713);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1714);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1715);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1716);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1717);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1718);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1719);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1720);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1721);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => n1148, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1722);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => n1149, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1723);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1724);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => n1150, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1725);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n1151, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1726);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n1537);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n1531);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => n1528, QN => n737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n1533);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n1541);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n1526);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1727);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1728);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1729);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1730);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1731);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1732);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1733);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n697);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1734);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1735);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1736);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1738);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1741);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1742);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1743);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1744);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n1543);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n_1745);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n1536);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n_1746);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n1527);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n1530);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1747
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1748
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1749
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1750
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1751
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1752
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1753
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1754
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1755
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1756
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1757
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1758
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1759
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1760
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1761
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1762
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1763
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1764
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1765
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1766
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1767
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1768
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1769)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1770)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1771)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1772)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1773)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1774)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1775)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1776)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1777)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1778)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1779);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_30_port, QN => 
                           n_1780);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n753);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_28_port, QN => 
                           n_1781);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n751);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_26_port, QN => 
                           n_1782);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n750);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_24_port, QN => 
                           n_1783);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n749);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_22_port, QN => 
                           n_1784);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n748);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_20_port, QN => 
                           n_1785);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n747);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_18_port, QN => 
                           n_1786);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n746);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_16_port, QN => 
                           n_1787);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n745);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_14_port, QN => 
                           n_1788);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n752);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_12_port, QN => 
                           n_1789);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n744);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_10_port, QN => 
                           n_1790);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n743
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_8_port, QN => 
                           n_1791);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n742
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_6_port, QN => 
                           n_1792);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n741
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_1793);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_1794);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_1795);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1796);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1797);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => n1529, QN => n1534);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1798);
   U1244 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(0), ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   U1245 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(10), ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U1246 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(11), ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U1247 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(12), ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U1248 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(13), ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U1249 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(14), ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U1250 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(15), ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U1251 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U1252 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U1253 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U1254 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U1255 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U1256 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U1257 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(21), ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U1258 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(22), ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U1259 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(23), ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U1260 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(24), ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U1261 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(25), ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U1262 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(26), ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U1263 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(27), ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U1264 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(28), ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U1265 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(29), ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U1266 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U1267 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(30), ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U1268 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(31), ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U1269 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U1270 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U1271 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U1272 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U1273 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U1274 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(8), ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U1275 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => n1538, QN => cu_i_n26);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => n1540, QN => cu_i_n23);
   cu_i_stall_reg : DFFR_X2 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n704, QN => n1535);
   U1276 : NOR2_X1 port map( A1 => n1528, A2 => 
                           curr_instruction_to_cu_i_31_port, ZN => n1158);
   U1277 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           curr_instruction_to_cu_i_30_port, A3 => n1160, A4 =>
                           n1289, ZN => n1296);
   U1278 : NOR3_X1 port map( A1 => n1537, A2 => n1156, A3 => n1526, ZN => 
                           cu_i_cmd_word_4_port);
   U1279 : AOI21_X1 port map( B1 => n1415, B2 => n1414, A => cu_i_cw3_6_port, 
                           ZN => n1416);
   U1280 : OAI21_X1 port map( B1 => n1281, B2 => n1282, A => n699, ZN => 
                           write_rf_i);
   U1281 : NAND2_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, ZN => n1161);
   U1282 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U1283 : NAND2_X1 port map( A1 => n1161, A2 => n1539, ZN => n1281);
   U1284 : NOR2_X1 port map( A1 => cu_i_n123, A2 => n1540, ZN => n1284);
   U1285 : AOI22_X1 port map( A1 => n704, A2 => n310, B1 => cu_i_cw1_13_port, 
                           B2 => n1535, ZN => n1488);
   U1286 : CLKBUF_X1 port map( A => n1525, Z => n1514);
   U1287 : CLKBUF_X1 port map( A => n1403, Z => n1223);
   U1288 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n1534, ZN => n1403);
   U1289 : CLKBUF_X1 port map( A => n1360, Z => n1409);
   U1290 : AOI21_X1 port map( B1 => n1171, B2 => n1249, A => n1240, ZN => n1412
                           );
   U1291 : NOR3_X1 port map( A1 => n1527, A2 => n1530, A3 => n1162, ZN => n1249
                           );
   U1292 : INV_X1 port map( A => n704, ZN => n1306);
   U1293 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n1284, A3 => n1533, A4 => n1531, ZN => n1156);
   U1294 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n1533, ZN => n1157);
   U1295 : NAND4_X1 port map( A1 => n1158, A2 => n1284, A3 => n1157, A4 => 
                           n1531, ZN => n1456);
   U1296 : NOR2_X1 port map( A1 => n1456, A2 => n1526, ZN => 
                           cu_i_cmd_word_7_port);
   U1297 : INV_X1 port map( A => n1158, ZN => n1160);
   U1298 : NOR2_X1 port map( A1 => n1160, A2 => n1156, ZN => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic);
   U1299 : NAND2_X1 port map( A1 => n1157, A2 => n1526, ZN => n1266);
   U1300 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => n737
                           , A3 => curr_instruction_to_cu_i_27_port, A4 => 
                           n1531, ZN => n1241);
   U1301 : NAND2_X1 port map( A1 => n1533, A2 => n1526, ZN => n1289);
   U1302 : NAND2_X1 port map( A1 => n1241, A2 => n1289, ZN => n1259);
   U1303 : NAND3_X1 port map( A1 => n1537, A2 => n1528, A3 => n1531, ZN => 
                           n1271);
   U1304 : INV_X1 port map( A => n1271, ZN => n1283);
   U1305 : OAI21_X1 port map( B1 => n1157, B2 => n1526, A => n1283, ZN => n1159
                           );
   U1306 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n1158, A3 => curr_instruction_to_cu_i_30_port, A4 =>
                           n1526, ZN => n1276);
   U1307 : AND3_X1 port map( A1 => n1259, A2 => n1159, A3 => n1276, ZN => n1293
                           );
   U1308 : OAI21_X1 port map( B1 => n1160, B2 => n1266, A => n1293, ZN => n1291
                           );
   U1309 : AOI211_X1 port map( C1 => n1284, C2 => n1291, A => 
                           cu_i_cmd_word_4_port, B => cu_i_cmd_word_7_port, ZN 
                           => n1248);
   U1310 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n1455);
   U1311 : NAND2_X1 port map( A1 => n1248, A2 => n1455, ZN => n310);
   U1312 : NAND2_X1 port map( A1 => n1284, A2 => n1296, ZN => n1240);
   U1313 : INV_X1 port map( A => n1240, ZN => n1286);
   U1314 : OR2_X1 port map( A1 => n310, A2 => n1286, ZN => cu_i_N278);
   U1315 : OAI22_X1 port map( A1 => n1535, A2 => cu_i_cmd_word_4_port, B1 => 
                           cu_i_cw2_8_port, B2 => n704, ZN => n309);
   U1316 : INV_X1 port map( A => n309, ZN => DRAM_ENABLE_port);
   U1317 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n1546);
   U1318 : INV_X1 port map( A => cu_i_cmd_word_4_port, ZN => n1410);
   U1319 : NOR2_X1 port map( A1 => n1528, A2 => n1410, ZN => 
                           cu_i_cmd_word_3_port);
   U1320 : OAI22_X1 port map( A1 => n1535, A2 => cu_i_cmd_word_3_port, B1 => 
                           cu_i_cw2_7_port, B2 => n704, ZN => n1250);
   U1321 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n1250, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U1322 : CLKBUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n1548);
   U1323 : NAND4_X1 port map( A1 => cu_i_n26, A2 => cu_i_n25, A3 => n1532, A4 
                           => n1539, ZN => cu_i_n145);
   U1324 : INV_X1 port map( A => n1455, ZN => n1549);
   U1325 : NAND2_X1 port map( A1 => cu_i_n145, A2 => n1281, ZN => n1171);
   U1326 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => 
                           curr_instruction_to_cu_i_5_port, A3 => 
                           curr_instruction_to_cu_i_2_port, A4 => 
                           curr_instruction_to_cu_i_3_port, ZN => n1162);
   U1327 : INV_X1 port map( A => n1412, ZN => n1411);
   U1328 : AOI221_X1 port map( B1 => n1411, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n1412, C2 =>
                           curr_instruction_to_cu_i_11_port, A => n1549, ZN => 
                           n1163);
   U1329 : INV_X1 port map( A => n1163, ZN => n1151);
   U1330 : AOI221_X1 port map( B1 => n1411, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n1412, C2 =>
                           curr_instruction_to_cu_i_12_port, A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n1164);
   U1331 : INV_X1 port map( A => n1164, ZN => n1150);
   U1332 : AOI221_X1 port map( B1 => n1411, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n1412, C2 =>
                           curr_instruction_to_cu_i_14_port, A => n1549, ZN => 
                           n1165);
   U1333 : INV_X1 port map( A => n1165, ZN => n1149);
   U1334 : AOI221_X1 port map( B1 => n1411, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n1412, C2 =>
                           curr_instruction_to_cu_i_15_port, A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n1166);
   U1335 : INV_X1 port map( A => n1166, ZN => n1148);
   U1336 : NOR2_X1 port map( A1 => n1529, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n1400);
   U1337 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_2_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_2_port, ZN => 
                           n1167);
   U1338 : OAI21_X1 port map( B1 => n728, B2 => n1403, A => n1167, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U1339 : INV_X1 port map( A => n1534, ZN => n1401);
   U1340 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_3_port, ZN => 
                           n1168);
   U1341 : OAI21_X1 port map( B1 => n729, B2 => n1223, A => n1168, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U1342 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_5_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_5_port, ZN => 
                           n1169);
   U1343 : OAI21_X1 port map( B1 => n731, B2 => n1403, A => n1169, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U1344 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_4_port, ZN => 
                           n1170);
   U1345 : OAI21_X1 port map( B1 => n730, B2 => n1223, A => n1170, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U1346 : NAND2_X1 port map( A1 => n1455, A2 => n1456, ZN => n1152);
   U1347 : NAND2_X1 port map( A1 => n1249, A2 => n1296, ZN => n1243);
   U1348 : OAI21_X1 port map( B1 => n1171, B2 => n1243, A => n1284, ZN => n1172
                           );
   U1349 : NAND2_X1 port map( A1 => cu_i_n123, A2 => n1540, ZN => n1300);
   U1350 : AOI21_X1 port map( B1 => n1172, B2 => n1300, A => n704, ZN => 
                           IRAM_ENABLE_port);
   U1351 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN
                           => n1173);
   U1352 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_3_port, ZN =>
                           n1315);
   U1353 : INV_X1 port map( A => n1152, ZN => n1301);
   U1354 : OAI221_X1 port map( B1 => n1535, B2 => n1301, C1 => n704, C2 => n756
                           , A => n1534, ZN => n1312);
   U1355 : INV_X1 port map( A => n1312, ZN => n1360);
   U1356 : NOR2_X1 port map( A1 => n1173, A2 => n1315, ZN => n1322);
   U1357 : AOI211_X1 port map( C1 => n1173, C2 => n1315, A => n1360, B => n1322
                           , ZN => n1175);
   U1358 : NAND2_X1 port map( A1 => IRAM_ENABLE_port, A2 => IRAM_ADDRESS_2_port
                           , ZN => n1309);
   U1359 : INV_X1 port map( A => n1309, ZN => n1311);
   U1360 : AND2_X1 port map( A1 => n1311, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n1318);
   U1361 : NAND2_X1 port map( A1 => n1318, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n1317);
   U1362 : NOR2_X1 port map( A1 => n741, A2 => n1317, ZN => n1324);
   U1363 : AOI211_X1 port map( C1 => n741, C2 => n1317, A => n1324, B => n1312,
                           ZN => n1174);
   U1364 : OR2_X1 port map( A1 => n1175, A2 => n1174, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U1365 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_7_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_7_port, ZN => 
                           n1176);
   U1366 : OAI21_X1 port map( B1 => n705, B2 => n1223, A => n1176, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U1367 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_6_port, ZN => 
                           n1177);
   U1368 : OAI21_X1 port map( B1 => n732, B2 => n1403, A => n1177, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U1369 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN
                           => n1178);
   U1370 : NAND2_X1 port map( A1 => n1322, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n1321);
   U1371 : NOR2_X1 port map( A1 => n1178, A2 => n1321, ZN => n1328);
   U1372 : AOI211_X1 port map( C1 => n1178, C2 => n1321, A => n1360, B => n1328
                           , ZN => n1180);
   U1373 : NAND2_X1 port map( A1 => n1324, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n1323);
   U1374 : NOR2_X1 port map( A1 => n742, A2 => n1323, ZN => n1330);
   U1375 : INV_X1 port map( A => n1409, ZN => n1406);
   U1376 : AOI211_X1 port map( C1 => n742, C2 => n1323, A => n1330, B => n1406,
                           ZN => n1179);
   U1377 : OR2_X1 port map( A1 => n1180, A2 => n1179, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U1378 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_9_port, B1 => n1400, B2 
                           => datapath_i_new_pc_value_decode_9_port, ZN => 
                           n1181);
   U1379 : OAI21_X1 port map( B1 => n707, B2 => n1403, A => n1181, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U1380 : CLKBUF_X1 port map( A => n1400, Z => n1394);
   U1381 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_8_port, B1 => n1394, B2 
                           => datapath_i_new_pc_value_decode_8_port, ZN => 
                           n1182);
   U1382 : OAI21_X1 port map( B1 => n706, B2 => n1223, A => n1182, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U1383 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN
                           => n1183);
   U1384 : NAND2_X1 port map( A1 => n1328, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n1327);
   U1385 : NOR2_X1 port map( A1 => n1183, A2 => n1327, ZN => n1334);
   U1386 : AOI211_X1 port map( C1 => n1183, C2 => n1327, A => n1360, B => n1334
                           , ZN => n1185);
   U1387 : NAND2_X1 port map( A1 => n1330, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n1329);
   U1388 : NOR2_X1 port map( A1 => n743, A2 => n1329, ZN => n1336);
   U1389 : AOI211_X1 port map( C1 => n743, C2 => n1329, A => n1336, B => n1406,
                           ZN => n1184);
   U1390 : OR2_X1 port map( A1 => n1185, A2 => n1184, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U1391 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_11_port, B1 => n1400, B2
                           => datapath_i_new_pc_value_decode_11_port, ZN => 
                           n1186);
   U1392 : OAI21_X1 port map( B1 => n709, B2 => n1223, A => n1186, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U1393 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_10_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_10_port, ZN => 
                           n1187);
   U1394 : OAI21_X1 port map( B1 => n708, B2 => n1403, A => n1187, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U1395 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, 
                           ZN => n1188);
   U1396 : NAND2_X1 port map( A1 => n1334, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n1333);
   U1397 : NOR2_X1 port map( A1 => n1188, A2 => n1333, ZN => n1340);
   U1398 : AOI211_X1 port map( C1 => n1188, C2 => n1333, A => n1360, B => n1340
                           , ZN => n1190);
   U1399 : NAND2_X1 port map( A1 => n1336, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n1335);
   U1400 : NOR2_X1 port map( A1 => n744, A2 => n1335, ZN => n1342);
   U1401 : AOI211_X1 port map( C1 => n744, C2 => n1335, A => n1342, B => n1312,
                           ZN => n1189);
   U1402 : OR2_X1 port map( A1 => n1190, A2 => n1189, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U1403 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_13_port, ZN => 
                           n1191);
   U1404 : OAI21_X1 port map( B1 => n711, B2 => n1403, A => n1191, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U1405 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_12_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_12_port, ZN => 
                           n1192);
   U1406 : OAI21_X1 port map( B1 => n710, B2 => n1403, A => n1192, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U1407 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, 
                           ZN => n1193);
   U1408 : NAND2_X1 port map( A1 => n1340, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n1339);
   U1409 : NOR2_X1 port map( A1 => n1193, A2 => n1339, ZN => n1346);
   U1410 : AOI211_X1 port map( C1 => n1193, C2 => n1339, A => n1409, B => n1346
                           , ZN => n1195);
   U1411 : NAND2_X1 port map( A1 => n1342, A2 => IRAM_ADDRESS_12_port, ZN => 
                           n1341);
   U1412 : NOR2_X1 port map( A1 => n752, A2 => n1341, ZN => n1348);
   U1413 : AOI211_X1 port map( C1 => n752, C2 => n1341, A => n1348, B => n1312,
                           ZN => n1194);
   U1414 : OR2_X1 port map( A1 => n1195, A2 => n1194, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U1415 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_15_port, ZN => 
                           n1196);
   U1416 : OAI21_X1 port map( B1 => n713, B2 => n1223, A => n1196, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U1417 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_14_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_14_port, ZN => 
                           n1197);
   U1418 : OAI21_X1 port map( B1 => n712, B2 => n1223, A => n1197, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U1419 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, 
                           ZN => n1198);
   U1420 : NAND2_X1 port map( A1 => n1346, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n1345);
   U1421 : NOR2_X1 port map( A1 => n1198, A2 => n1345, ZN => n1352);
   U1422 : AOI211_X1 port map( C1 => n1198, C2 => n1345, A => n1360, B => n1352
                           , ZN => n1200);
   U1423 : NAND2_X1 port map( A1 => n1348, A2 => IRAM_ADDRESS_14_port, ZN => 
                           n1347);
   U1424 : NOR2_X1 port map( A1 => n745, A2 => n1347, ZN => n1354);
   U1425 : AOI211_X1 port map( C1 => n745, C2 => n1347, A => n1354, B => n1406,
                           ZN => n1199);
   U1426 : OR2_X1 port map( A1 => n1200, A2 => n1199, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U1427 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_17_port, ZN => 
                           n1201);
   U1428 : OAI21_X1 port map( B1 => n715, B2 => n1223, A => n1201, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U1429 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_16_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_16_port, ZN => 
                           n1202);
   U1430 : OAI21_X1 port map( B1 => n714, B2 => n1223, A => n1202, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U1431 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, 
                           ZN => n1203);
   U1432 : NAND2_X1 port map( A1 => n1352, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n1351);
   U1433 : NOR2_X1 port map( A1 => n1203, A2 => n1351, ZN => n1358);
   U1434 : AOI211_X1 port map( C1 => n1203, C2 => n1351, A => n1360, B => n1358
                           , ZN => n1205);
   U1435 : NAND2_X1 port map( A1 => n1354, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n1353);
   U1436 : NOR2_X1 port map( A1 => n746, A2 => n1353, ZN => n1361);
   U1437 : AOI211_X1 port map( C1 => n746, C2 => n1353, A => n1361, B => n1406,
                           ZN => n1204);
   U1438 : OR2_X1 port map( A1 => n1205, A2 => n1204, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U1439 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_19_port, ZN => 
                           n1206);
   U1440 : OAI21_X1 port map( B1 => n717, B2 => n1223, A => n1206, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U1441 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_18_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_18_port, ZN => 
                           n1207);
   U1442 : OAI21_X1 port map( B1 => n716, B2 => n1223, A => n1207, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U1443 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, 
                           ZN => n1208);
   U1444 : NAND2_X1 port map( A1 => n1358, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n1357);
   U1445 : NOR2_X1 port map( A1 => n1208, A2 => n1357, ZN => n1365);
   U1446 : AOI211_X1 port map( C1 => n1208, C2 => n1357, A => n1360, B => n1365
                           , ZN => n1210);
   U1447 : NAND2_X1 port map( A1 => n1361, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n1359);
   U1448 : NOR2_X1 port map( A1 => n747, A2 => n1359, ZN => n1367);
   U1449 : AOI211_X1 port map( C1 => n747, C2 => n1359, A => n1367, B => n1406,
                           ZN => n1209);
   U1450 : OR2_X1 port map( A1 => n1210, A2 => n1209, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U1451 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_21_port, ZN => 
                           n1211);
   U1452 : OAI21_X1 port map( B1 => n719, B2 => n1223, A => n1211, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U1453 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_20_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_20_port, ZN => 
                           n1212);
   U1454 : OAI21_X1 port map( B1 => n718, B2 => n1223, A => n1212, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U1455 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, 
                           ZN => n1213);
   U1456 : NAND2_X1 port map( A1 => n1365, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n1364);
   U1457 : NOR2_X1 port map( A1 => n1213, A2 => n1364, ZN => n1371);
   U1458 : AOI211_X1 port map( C1 => n1213, C2 => n1364, A => n1360, B => n1371
                           , ZN => n1215);
   U1459 : NAND2_X1 port map( A1 => n1367, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n1366);
   U1460 : NOR2_X1 port map( A1 => n748, A2 => n1366, ZN => n1373);
   U1461 : AOI211_X1 port map( C1 => n748, C2 => n1366, A => n1373, B => n1406,
                           ZN => n1214);
   U1462 : OR2_X1 port map( A1 => n1215, A2 => n1214, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U1463 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n1400, B2
                           => datapath_i_new_pc_value_decode_23_port, ZN => 
                           n1216);
   U1464 : OAI21_X1 port map( B1 => n721, B2 => n1223, A => n1216, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U1465 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_22_port, B1 => n1400, B2
                           => datapath_i_new_pc_value_decode_22_port, ZN => 
                           n1217);
   U1466 : OAI21_X1 port map( B1 => n720, B2 => n1223, A => n1217, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U1467 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, 
                           ZN => n1218);
   U1468 : NAND2_X1 port map( A1 => n1371, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n1370);
   U1469 : NOR2_X1 port map( A1 => n1218, A2 => n1370, ZN => n1377);
   U1470 : AOI211_X1 port map( C1 => n1218, C2 => n1370, A => n1360, B => n1377
                           , ZN => n1220);
   U1471 : NAND2_X1 port map( A1 => n1373, A2 => IRAM_ADDRESS_22_port, ZN => 
                           n1372);
   U1472 : NOR2_X1 port map( A1 => n749, A2 => n1372, ZN => n1379);
   U1473 : AOI211_X1 port map( C1 => n749, C2 => n1372, A => n1379, B => n1312,
                           ZN => n1219);
   U1474 : OR2_X1 port map( A1 => n1220, A2 => n1219, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U1475 : AOI22_X1 port map( A1 => n1529, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_25_port, ZN => 
                           n1221);
   U1476 : OAI21_X1 port map( B1 => n723, B2 => n1223, A => n1221, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U1477 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_24_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_24_port, ZN => 
                           n1222);
   U1478 : OAI21_X1 port map( B1 => n722, B2 => n1223, A => n1222, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U1479 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, 
                           ZN => n1224);
   U1480 : NAND2_X1 port map( A1 => n1377, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n1376);
   U1481 : NOR2_X1 port map( A1 => n1224, A2 => n1376, ZN => n1383);
   U1482 : AOI211_X1 port map( C1 => n1224, C2 => n1376, A => n1409, B => n1383
                           , ZN => n1226);
   U1483 : NAND2_X1 port map( A1 => n1379, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n1378);
   U1484 : NOR2_X1 port map( A1 => n750, A2 => n1378, ZN => n1385);
   U1485 : AOI211_X1 port map( C1 => n750, C2 => n1378, A => n1385, B => n1312,
                           ZN => n1225);
   U1486 : OR2_X1 port map( A1 => n1226, A2 => n1225, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U1487 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_27_port, ZN => 
                           n1227);
   U1488 : OAI21_X1 port map( B1 => n724, B2 => n1403, A => n1227, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U1489 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_26_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_26_port, ZN => 
                           n1228);
   U1490 : OAI21_X1 port map( B1 => n691, B2 => n1403, A => n1228, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U1491 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, 
                           ZN => n1229);
   U1492 : NAND2_X1 port map( A1 => n1383, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n1382);
   U1493 : NOR2_X1 port map( A1 => n1229, A2 => n1382, ZN => n1389);
   U1494 : AOI211_X1 port map( C1 => n1229, C2 => n1382, A => n1409, B => n1389
                           , ZN => n1231);
   U1495 : NAND2_X1 port map( A1 => n1385, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n1384);
   U1496 : NOR2_X1 port map( A1 => n751, A2 => n1384, ZN => n1391);
   U1497 : AOI211_X1 port map( C1 => n751, C2 => n1384, A => n1391, B => n1312,
                           ZN => n1230);
   U1498 : OR2_X1 port map( A1 => n1231, A2 => n1230, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U1499 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_29_port, ZN => 
                           n1232);
   U1500 : OAI21_X1 port map( B1 => n726, B2 => n1403, A => n1232, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U1501 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_28_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_28_port, ZN => 
                           n1233);
   U1502 : OAI21_X1 port map( B1 => n725, B2 => n1403, A => n1233, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U1503 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, 
                           ZN => n1234);
   U1504 : NAND2_X1 port map( A1 => n1389, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n1388);
   U1505 : NOR2_X1 port map( A1 => n1234, A2 => n1388, ZN => n1396);
   U1506 : AOI211_X1 port map( C1 => n1234, C2 => n1388, A => n1409, B => n1396
                           , ZN => n1236);
   U1507 : NAND2_X1 port map( A1 => n1391, A2 => IRAM_ADDRESS_28_port, ZN => 
                           n1390);
   U1508 : NOR2_X1 port map( A1 => n753, A2 => n1390, ZN => n1397);
   U1509 : AOI211_X1 port map( C1 => n753, C2 => n1390, A => n1397, B => n1406,
                           ZN => n1235);
   U1510 : OR2_X1 port map( A1 => n1236, A2 => n1235, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U1511 : OAI22_X1 port map( A1 => n1535, A2 => cu_i_cw3_6_port, B1 => 
                           cu_i_cw2_6_port, B2 => n704, ZN => n1237);
   U1512 : INV_X1 port map( A => n1237, ZN => n1155);
   U1513 : CLKBUF_X1 port map( A => n310, Z => n1545);
   U1514 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_0_port, B1
                           => cu_i_cw1_0_port, B2 => n1535, ZN => n1252);
   U1515 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_1_port, B1
                           => cu_i_cw1_1_port, B2 => n1535, ZN => n1254);
   U1516 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_3_port, B1
                           => cu_i_cw1_3_port, B2 => n1535, ZN => n1251);
   U1517 : INV_X1 port map( A => n1251, ZN => n1471);
   U1518 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_2_port, B1
                           => cu_i_cw1_2_port, B2 => n1306, ZN => n1472);
   U1519 : OAI211_X1 port map( C1 => n1252, C2 => n1254, A => n1471, B => n1472
                           , ZN => n1238);
   U1520 : INV_X1 port map( A => n1238, ZN => n1147);
   U1521 : AOI21_X1 port map( B1 => n1472, B2 => n1254, A => n1251, ZN => n1239
                           );
   U1522 : NOR2_X1 port map( A1 => n1252, A2 => n1239, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U1523 : INV_X1 port map( A => n1284, ZN => n1302);
   U1524 : OAI222_X1 port map( A1 => n1526, A2 => n1455, B1 => n1240, B2 => 
                           n1249, C1 => n1302, C2 => n1293, ZN => n311);
   U1525 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n311, ZN => 
                           cu_i_cmd_word_1_port);
   U1526 : INV_X1 port map( A => n1296, ZN => n1298);
   U1527 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => n1543
                           , A3 => n1298, ZN => n1274);
   U1528 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           n1274, A3 => n1527, ZN => n1260);
   U1529 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n1530
                           , A3 => n1260, ZN => n1247);
   U1530 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => 
                           n1241, A3 => n1533, ZN => n1242);
   U1531 : OAI211_X1 port map( C1 => n1266, C2 => n1271, A => n1243, B => n1242
                           , ZN => n1246);
   U1532 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => n1298
                           , ZN => n1244);
   U1533 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => 
                           n1244, A3 => n1530, A4 => n1536, ZN => n1278);
   U1534 : OAI221_X1 port map( B1 => n1278, B2 => 
                           curr_instruction_to_cu_i_5_port, C1 => n1278, C2 => 
                           curr_instruction_to_cu_i_1_port, A => n1276, ZN => 
                           n1245);
   U1535 : OR3_X1 port map( A1 => n1247, A2 => n1246, A3 => n1245, ZN => 
                           cu_i_N265);
   U1536 : NAND2_X1 port map( A1 => n1248, A2 => n1411, ZN => enable_rf_i);
   U1537 : NAND2_X1 port map( A1 => n1249, A2 => n1286, ZN => n1282);
   U1538 : AND2_X1 port map( A1 => n310, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U1539 : INV_X1 port map( A => n1250, ZN => DRAM_READNOTWRITE);
   U1540 : MUX2_X1 port map( A => datapath_i_val_immediate_i_3_port, B => 
                           datapath_i_val_b_i_3_port, S => n1488, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U1541 : AOI21_X1 port map( B1 => n1472, B2 => n1252, A => n1251, ZN => n1253
                           );
   U1542 : NOR2_X1 port map( A1 => n1254, A2 => n1253, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U1543 : NOR2_X1 port map( A1 => n1532, A2 => n1282, ZN => cu_i_N273);
   U1544 : INV_X1 port map( A => n1282, ZN => n1414);
   U1545 : AOI221_X1 port map( B1 => cu_i_n25, B2 => n1414, C1 => cu_i_n26, C2 
                           => n1414, A => cu_i_N273, ZN => n1255);
   U1546 : INV_X1 port map( A => n1255, ZN => n1258);
   U1547 : NOR2_X1 port map( A1 => cu_i_n125, A2 => n1282, ZN => n1256);
   U1548 : NAND2_X1 port map( A1 => n1256, A2 => n1538, ZN => n1280);
   U1549 : NOR2_X1 port map( A1 => cu_i_n25, A2 => n1280, ZN => n1257);
   U1550 : MUX2_X1 port map( A => n1258, B => n1257, S => cu_i_n124, Z => 
                           cu_i_N277);
   U1551 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           curr_instruction_to_cu_i_2_port, ZN => n1261);
   U1552 : OAI21_X1 port map( B1 => n1261, B2 => n1260, A => n1259, ZN => 
                           cu_i_N267);
   datapath_i_execute_stage_dp_n9 <= '0';
   U1554 : NOR2_X1 port map( A1 => n1535, A2 => n1152, ZN => n1262);
   U1555 : NOR2_X1 port map( A1 => n704, A2 => cu_i_cw1_4_port, ZN => n1290);
   U1556 : NOR2_X1 port map( A1 => n1262, A2 => n1290, ZN => n1263);
   U1557 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n1263, ZN => n1525);
   U1558 : INV_X1 port map( A => n1263, ZN => n1510);
   U1559 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n1510, ZN => n1523);
   U1560 : CLKBUF_X1 port map( A => n1523, Z => n1512);
   U1561 : CLKBUF_X1 port map( A => n1510, Z => n1522);
   U1562 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n1522, ZN => n1264);
   U1563 : OAI21_X1 port map( B1 => n691, B2 => n1514, A => n1264, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U1564 : INV_X1 port map( A => n1488, ZN => n1485);
   U1565 : CLKBUF_X1 port map( A => n1485, Z => n1487);
   U1566 : MUX2_X1 port map( A => datapath_i_val_b_i_0_port, B => 
                           datapath_i_val_immediate_i_0_port, S => n1487, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U1567 : MUX2_X1 port map( A => datapath_i_val_b_i_2_port, B => 
                           datapath_i_val_immediate_i_2_port, S => n1485, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U1568 : OAI221_X1 port map( B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           curr_instruction_to_cu_i_2_port, C1 => n1527, C2 => 
                           n1536, A => n1274, ZN => n1270);
   U1569 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n1271, A => n1276, ZN => n1268);
   U1570 : NAND2_X1 port map( A1 => n1537, A2 => n1528, ZN => n1265);
   U1571 : OAI22_X1 port map( A1 => n1527, A2 => n1278, B1 => n1266, B2 => 
                           n1265, ZN => n1267);
   U1572 : AOI21_X1 port map( B1 => curr_instruction_to_cu_i_27_port, B2 => 
                           n1268, A => n1267, ZN => n1269);
   U1573 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_0_port, B2 => 
                           n1270, A => n1269, ZN => cu_i_N264);
   U1574 : AOI221_X1 port map( B1 => curr_instruction_to_cu_i_27_port, B2 => 
                           curr_instruction_to_cu_i_26_port, C1 => n1541, C2 =>
                           n1526, A => n1271, ZN => n1275);
   U1575 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => 
                           n1536, ZN => n1272);
   U1576 : AOI221_X1 port map( B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           curr_instruction_to_cu_i_0_port, C1 => n1527, C2 => 
                           n1530, A => n1272, ZN => n1273);
   U1577 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n1275, B1 => n1274, B2 => n1273, ZN => n1277);
   U1578 : OAI211_X1 port map( C1 => curr_instruction_to_cu_i_5_port, C2 => 
                           n1278, A => n1277, B => n1276, ZN => cu_i_N266);
   U1579 : NAND2_X1 port map( A1 => n704, A2 => n1282, ZN => cu_i_N274);
   U1580 : AOI221_X1 port map( B1 => cu_i_n125, B2 => cu_i_n26, C1 => n1532, C2
                           => n1538, A => n1282, ZN => cu_i_N275);
   U1581 : OAI21_X1 port map( B1 => cu_i_n26, B2 => cu_i_n125, A => n1414, ZN 
                           => n1279);
   U1582 : AOI22_X1 port map( A1 => cu_i_n25, A2 => n1280, B1 => n1279, B2 => 
                           n1542, ZN => cu_i_N276);
   U1583 : INV_X1 port map( A => n1281, ZN => n1415);
   U1584 : AOI211_X1 port map( C1 => n704, C2 => cu_i_n145, A => n1415, B => 
                           n1282, ZN => cu_i_N279);
   U1585 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n1284, A3 => n1283, ZN => n1288);
   U1586 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => 
                           curr_instruction_to_cu_i_0_port, A3 => 
                           curr_instruction_to_cu_i_2_port, A4 => 
                           curr_instruction_to_cu_i_3_port, ZN => n1285);
   U1587 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => 
                           curr_instruction_to_cu_i_5_port, A3 => n1286, A4 => 
                           n1285, ZN => n1287);
   U1588 : OAI21_X1 port map( B1 => n1289, B2 => n1288, A => n1287, ZN => 
                           cu_i_cmd_word_8_port);
   U1589 : MUX2_X1 port map( A => cu_i_cmd_word_8_port, B => cu_i_cw1_12_port, 
                           S => n1306, Z => alu_cin_i);
   U1590 : AOI21_X1 port map( B1 => n756, B2 => n704, A => n1290, ZN => 
                           cu_i_cw1_i_4_port);
   U1591 : MUX2_X1 port map( A => cu_i_cw2_7_port, B => cu_i_cw1_7_port, S => 
                           n1535, Z => cu_i_cw1_i_7_port);
   U1592 : MUX2_X1 port map( A => cu_i_cw2_8_port, B => cu_i_cw1_8_port, S => 
                           n1535, Z => cu_i_cw1_i_8_port);
   U1593 : INV_X1 port map( A => n1291, ZN => n1299);
   U1594 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_12_port, A2 => 
                           curr_instruction_to_cu_i_11_port, A3 => 
                           curr_instruction_to_cu_i_15_port, A4 => 
                           curr_instruction_to_cu_i_14_port, ZN => n1292);
   U1595 : NAND2_X1 port map( A1 => n740, A2 => n1292, ZN => n1297);
   U1596 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_17_port, A2 => 
                           curr_instruction_to_cu_i_16_port, A3 => 
                           curr_instruction_to_cu_i_20_port, A4 => 
                           curr_instruction_to_cu_i_19_port, ZN => n1294);
   U1597 : AOI21_X1 port map( B1 => n697, B2 => n1294, A => n1293, ZN => n1295)
                           ;
   U1598 : AOI221_X1 port map( B1 => n1299, B2 => n1298, C1 => n1297, C2 => 
                           n1296, A => n1295, ZN => n1303);
   U1599 : OAI211_X1 port map( C1 => n1303, C2 => n1302, A => n1301, B => n1300
                           , ZN => cu_i_n209);
   U1600 : NOR2_X1 port map( A1 => cu_i_n123, A2 => cu_i_n23, ZN => cu_i_n210);
   U1601 : AOI22_X1 port map( A1 => n704, A2 => n699, B1 => n1544, B2 => n1306,
                           ZN => cu_i_n131);
   U1602 : MUX2_X1 port map( A => cu_i_cw2_6_port, B => cu_i_cw1_6_port, S => 
                           n1306, Z => cu_i_n127);
   U1603 : MUX2_X1 port map( A => cu_i_cw2_5_port, B => cu_i_cw1_5_port, S => 
                           n1306, Z => cu_i_n126);
   U1604 : MUX2_X1 port map( A => curr_instruction_to_cu_i_31_port, B => 
                           IRAM_DATA(31), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U1605 : MUX2_X1 port map( A => curr_instruction_to_cu_i_30_port, B => 
                           IRAM_DATA(30), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U1606 : MUX2_X1 port map( A => n1528, B => IRAM_DATA(29), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U1607 : MUX2_X1 port map( A => curr_instruction_to_cu_i_28_port, B => 
                           IRAM_DATA(28), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U1608 : MUX2_X1 port map( A => curr_instruction_to_cu_i_27_port, B => 
                           IRAM_DATA(27), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U1609 : MUX2_X1 port map( A => curr_instruction_to_cu_i_26_port, B => 
                           IRAM_DATA(26), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U1610 : MUX2_X1 port map( A => datapath_i_n9, B => IRAM_DATA(25), S => n1306
                           , Z => datapath_i_fetch_stage_dp_n63);
   U1611 : MUX2_X1 port map( A => datapath_i_n10, B => IRAM_DATA(24), S => 
                           n1306, Z => datapath_i_fetch_stage_dp_n62);
   U1612 : MUX2_X1 port map( A => datapath_i_n11, B => IRAM_DATA(23), S => 
                           n1306, Z => datapath_i_fetch_stage_dp_n61);
   U1613 : MUX2_X1 port map( A => datapath_i_n12, B => IRAM_DATA(22), S => 
                           n1535, Z => datapath_i_fetch_stage_dp_n60);
   U1614 : MUX2_X1 port map( A => datapath_i_n13, B => IRAM_DATA(21), S => 
                           n1535, Z => datapath_i_fetch_stage_dp_n59);
   U1615 : MUX2_X1 port map( A => curr_instruction_to_cu_i_20_port, B => 
                           IRAM_DATA(20), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U1616 : MUX2_X1 port map( A => curr_instruction_to_cu_i_19_port, B => 
                           IRAM_DATA(19), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U1617 : NAND2_X1 port map( A1 => n1535, A2 => IRAM_DATA(18), ZN => n1304);
   U1618 : OAI21_X1 port map( B1 => n1535, B2 => n697, A => n1304, ZN => 
                           datapath_i_fetch_stage_dp_n56);
   U1619 : MUX2_X1 port map( A => curr_instruction_to_cu_i_17_port, B => 
                           IRAM_DATA(17), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U1620 : MUX2_X1 port map( A => curr_instruction_to_cu_i_16_port, B => 
                           IRAM_DATA(16), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U1621 : MUX2_X1 port map( A => curr_instruction_to_cu_i_15_port, B => 
                           IRAM_DATA(15), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U1622 : MUX2_X1 port map( A => curr_instruction_to_cu_i_14_port, B => 
                           IRAM_DATA(14), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U1623 : NAND2_X1 port map( A1 => n1535, A2 => IRAM_DATA(13), ZN => n1305);
   U1624 : OAI21_X1 port map( B1 => n1306, B2 => n740, A => n1305, ZN => 
                           datapath_i_fetch_stage_dp_n51);
   U1625 : MUX2_X1 port map( A => curr_instruction_to_cu_i_12_port, B => 
                           IRAM_DATA(12), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U1626 : MUX2_X1 port map( A => curr_instruction_to_cu_i_11_port, B => 
                           IRAM_DATA(11), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U1627 : MUX2_X1 port map( A => datapath_i_n14, B => IRAM_DATA(10), S => 
                           n1306, Z => datapath_i_fetch_stage_dp_n48);
   U1628 : MUX2_X1 port map( A => datapath_i_n15, B => IRAM_DATA(9), S => n1306
                           , Z => datapath_i_fetch_stage_dp_n47);
   U1629 : MUX2_X1 port map( A => datapath_i_n16, B => IRAM_DATA(8), S => n1535
                           , Z => datapath_i_fetch_stage_dp_n46);
   U1630 : MUX2_X1 port map( A => datapath_i_n17, B => IRAM_DATA(7), S => n1306
                           , Z => datapath_i_fetch_stage_dp_n45);
   U1631 : MUX2_X1 port map( A => datapath_i_n18, B => IRAM_DATA(6), S => n1306
                           , Z => datapath_i_fetch_stage_dp_n44);
   U1632 : MUX2_X1 port map( A => curr_instruction_to_cu_i_5_port, B => 
                           IRAM_DATA(5), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U1633 : MUX2_X1 port map( A => curr_instruction_to_cu_i_4_port, B => 
                           IRAM_DATA(4), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U1634 : MUX2_X1 port map( A => curr_instruction_to_cu_i_3_port, B => 
                           IRAM_DATA(3), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U1635 : MUX2_X1 port map( A => curr_instruction_to_cu_i_2_port, B => 
                           IRAM_DATA(2), S => n1535, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U1636 : MUX2_X1 port map( A => curr_instruction_to_cu_i_1_port, B => 
                           IRAM_DATA(1), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U1637 : MUX2_X1 port map( A => curr_instruction_to_cu_i_0_port, B => 
                           IRAM_DATA(0), S => n1306, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U1638 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n1394, B2 
                           => datapath_i_new_pc_value_decode_0_port, ZN => 
                           n1307);
   U1639 : OAI21_X1 port map( B1 => n733, B2 => n1403, A => n1307, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U1640 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N39_port, B => 
                           datapath_i_fetch_stage_dp_N5, S => n1312, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U1641 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_1_port, B1 => n1394, B2 
                           => datapath_i_new_pc_value_decode_1_port, ZN => 
                           n1308);
   U1642 : OAI21_X1 port map( B1 => n734, B2 => n1403, A => n1308, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U1643 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N40_port, B => 
                           datapath_i_fetch_stage_dp_N6, S => n1312, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U1644 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n1309, ZN => n1310);
   U1645 : AOI22_X1 port map( A1 => n1409, A2 => n1310, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n1406, ZN => datapath_i_fetch_stage_dp_n35);
   U1646 : OAI21_X1 port map( B1 => n1311, B2 => IRAM_ADDRESS_3_port, A => 
                           n1360, ZN => n1314);
   U1647 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n1316);
   U1648 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           B2 => datapath_i_new_pc_value_mem_stage_i_3_port, A 
                           => n1312, ZN => n1313);
   U1649 : OAI22_X1 port map( A1 => n1318, A2 => n1314, B1 => n1316, B2 => 
                           n1313, ZN => datapath_i_fetch_stage_dp_n34);
   U1650 : OAI211_X1 port map( C1 => n1316, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n1406, B => n1315, ZN => n1320);
   U1651 : OAI211_X1 port map( C1 => n1318, C2 => IRAM_ADDRESS_4_port, A => 
                           n1409, B => n1317, ZN => n1319);
   U1652 : NAND2_X1 port map( A1 => n1320, A2 => n1319, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U1653 : OAI211_X1 port map( C1 => n1322, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n1406, B => n1321, ZN => n1326);
   U1654 : OAI211_X1 port map( C1 => n1324, C2 => IRAM_ADDRESS_6_port, A => 
                           n1409, B => n1323, ZN => n1325);
   U1655 : NAND2_X1 port map( A1 => n1326, A2 => n1325, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U1656 : OAI211_X1 port map( C1 => n1328, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n1406, B => n1327, ZN => n1332);
   U1657 : OAI211_X1 port map( C1 => n1330, C2 => IRAM_ADDRESS_8_port, A => 
                           n1409, B => n1329, ZN => n1331);
   U1658 : NAND2_X1 port map( A1 => n1332, A2 => n1331, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U1659 : OAI211_X1 port map( C1 => n1334, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n1406, B => n1333, ZN => n1338);
   U1660 : OAI211_X1 port map( C1 => n1336, C2 => IRAM_ADDRESS_10_port, A => 
                           n1409, B => n1335, ZN => n1337);
   U1661 : NAND2_X1 port map( A1 => n1338, A2 => n1337, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U1662 : OAI211_X1 port map( C1 => n1340, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n1406, B => n1339, ZN => n1344);
   U1663 : OAI211_X1 port map( C1 => n1342, C2 => IRAM_ADDRESS_12_port, A => 
                           n1360, B => n1341, ZN => n1343);
   U1664 : NAND2_X1 port map( A1 => n1344, A2 => n1343, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U1665 : OAI211_X1 port map( C1 => n1346, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n1406, B => n1345, ZN => n1350);
   U1666 : OAI211_X1 port map( C1 => n1348, C2 => IRAM_ADDRESS_14_port, A => 
                           n1360, B => n1347, ZN => n1349);
   U1667 : NAND2_X1 port map( A1 => n1350, A2 => n1349, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U1668 : OAI211_X1 port map( C1 => n1352, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n1406, B => n1351, ZN => n1356);
   U1669 : OAI211_X1 port map( C1 => n1354, C2 => IRAM_ADDRESS_16_port, A => 
                           n1360, B => n1353, ZN => n1355);
   U1670 : NAND2_X1 port map( A1 => n1356, A2 => n1355, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U1671 : OAI211_X1 port map( C1 => n1358, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n1406, B => n1357, ZN => n1363);
   U1672 : OAI211_X1 port map( C1 => n1361, C2 => IRAM_ADDRESS_18_port, A => 
                           n1360, B => n1359, ZN => n1362);
   U1673 : NAND2_X1 port map( A1 => n1363, A2 => n1362, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U1674 : OAI211_X1 port map( C1 => n1365, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n1406, B => n1364, ZN => n1369);
   U1675 : OAI211_X1 port map( C1 => n1367, C2 => IRAM_ADDRESS_20_port, A => 
                           n1409, B => n1366, ZN => n1368);
   U1676 : NAND2_X1 port map( A1 => n1369, A2 => n1368, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U1677 : OAI211_X1 port map( C1 => n1371, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n1406, B => n1370, ZN => n1375);
   U1678 : OAI211_X1 port map( C1 => n1373, C2 => IRAM_ADDRESS_22_port, A => 
                           n1409, B => n1372, ZN => n1374);
   U1679 : NAND2_X1 port map( A1 => n1375, A2 => n1374, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U1680 : OAI211_X1 port map( C1 => n1377, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n1406, B => n1376, ZN => n1381);
   U1681 : OAI211_X1 port map( C1 => n1379, C2 => IRAM_ADDRESS_24_port, A => 
                           n1409, B => n1378, ZN => n1380);
   U1682 : NAND2_X1 port map( A1 => n1381, A2 => n1380, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U1683 : OAI211_X1 port map( C1 => n1383, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n1406, B => n1382, ZN => n1387);
   U1684 : OAI211_X1 port map( C1 => n1385, C2 => IRAM_ADDRESS_26_port, A => 
                           n1409, B => n1384, ZN => n1386);
   U1685 : NAND2_X1 port map( A1 => n1387, A2 => n1386, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U1686 : OAI211_X1 port map( C1 => n1389, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n1406, B => n1388, ZN => n1393);
   U1687 : OAI211_X1 port map( C1 => n1391, C2 => IRAM_ADDRESS_28_port, A => 
                           n1409, B => n1390, ZN => n1392);
   U1688 : NAND2_X1 port map( A1 => n1393, A2 => n1392, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U1689 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_30_port, B1 => n1394, B2
                           => datapath_i_new_pc_value_decode_30_port, ZN => 
                           n1395);
   U1690 : OAI21_X1 port map( B1 => n727, B2 => n1403, A => n1395, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   U1691 : NAND2_X1 port map( A1 => n1396, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n1405);
   U1692 : OAI211_X1 port map( C1 => n1396, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n1406, B => n1405, ZN => n1399);
   U1693 : NAND2_X1 port map( A1 => n1397, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n1404);
   U1694 : OAI211_X1 port map( C1 => n1397, C2 => IRAM_ADDRESS_30_port, A => 
                           n1409, B => n1404, ZN => n1398);
   U1695 : NAND2_X1 port map( A1 => n1399, A2 => n1398, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U1696 : AOI22_X1 port map( A1 => n1401, A2 => 
                           datapath_i_alu_output_val_i_31_port, B1 => 
                           datapath_i_new_pc_value_decode_31_port, B2 => n1400,
                           ZN => n1402);
   U1697 : OAI21_X1 port map( B1 => n703, B2 => n1403, A => n1402, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U1698 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n1404, Z => n1408)
                           ;
   U1699 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n1405, Z => n1407);
   U1700 : AOI22_X1 port map( A1 => n1409, A2 => n1408, B1 => n1407, B2 => 
                           n1406, ZN => datapath_i_fetch_stage_dp_n2);
   U1701 : OAI21_X1 port map( B1 => n737, B2 => n1410, A => n1411, ZN => 
                           read_rf_p2_i);
   U1702 : OAI221_X1 port map( B1 => n1412, B2 => n697, C1 => n1411, C2 => n740
                           , A => n1455, ZN => datapath_i_decode_stage_dp_n78);
   U1703 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ZN => n1413);
   U1704 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n1413, ZN => n1429);
   U1705 : INV_X1 port map( A => n1429, ZN => n1438);
   U1706 : AND2_X2 port map( A1 => n1438, A2 => n1416, ZN => n1452);
   U1707 : NOR2_X1 port map( A1 => n1429, A2 => n1416, ZN => n1451);
   U1708 : CLKBUF_X1 port map( A => n1451, Z => n1442);
   U1709 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_0_port, ZN => n1417
                           );
   U1710 : OAI21_X1 port map( B1 => n733, B2 => n1438, A => n1417, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U1711 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_1_port, ZN => n1418
                           );
   U1712 : OAI21_X1 port map( B1 => n734, B2 => n1438, A => n1418, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U1713 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_2_port, ZN => n1419
                           );
   U1714 : OAI21_X1 port map( B1 => n728, B2 => n1438, A => n1419, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U1715 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_3_port, ZN => n1420
                           );
   U1716 : OAI21_X1 port map( B1 => n729, B2 => n1438, A => n1420, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U1717 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_4_port, ZN => n1421
                           );
   U1718 : OAI21_X1 port map( B1 => n730, B2 => n1438, A => n1421, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U1719 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_5_port, ZN => n1422
                           );
   U1720 : OAI21_X1 port map( B1 => n731, B2 => n1438, A => n1422, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U1721 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_6_port, ZN => n1423
                           );
   U1722 : OAI21_X1 port map( B1 => n732, B2 => n1438, A => n1423, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U1723 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_7_port, ZN => n1424
                           );
   U1724 : OAI21_X1 port map( B1 => n705, B2 => n1438, A => n1424, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U1725 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_8_port, ZN => n1425
                           );
   U1726 : OAI21_X1 port map( B1 => n706, B2 => n1438, A => n1425, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U1727 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_9_port, ZN => n1426
                           );
   U1728 : OAI21_X1 port map( B1 => n707, B2 => n1438, A => n1426, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U1729 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => 
                           n1427);
   U1730 : OAI21_X1 port map( B1 => n708, B2 => n1438, A => n1427, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U1731 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => 
                           n1428);
   U1732 : OAI21_X1 port map( B1 => n709, B2 => n1438, A => n1428, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U1733 : INV_X1 port map( A => n1429, ZN => n1454);
   U1734 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => 
                           n1430);
   U1735 : OAI21_X1 port map( B1 => n710, B2 => n1454, A => n1430, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U1736 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => 
                           n1431);
   U1737 : OAI21_X1 port map( B1 => n711, B2 => n1438, A => n1431, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U1738 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => 
                           n1432);
   U1739 : OAI21_X1 port map( B1 => n712, B2 => n1454, A => n1432, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U1740 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => 
                           n1433);
   U1741 : OAI21_X1 port map( B1 => n713, B2 => n1438, A => n1433, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U1742 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => 
                           n1434);
   U1743 : OAI21_X1 port map( B1 => n714, B2 => n1454, A => n1434, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U1744 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => 
                           n1435);
   U1745 : OAI21_X1 port map( B1 => n715, B2 => n1438, A => n1435, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U1746 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => 
                           n1436);
   U1747 : OAI21_X1 port map( B1 => n716, B2 => n1454, A => n1436, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U1748 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => 
                           n1437);
   U1749 : OAI21_X1 port map( B1 => n717, B2 => n1438, A => n1437, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U1750 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => 
                           n1439);
   U1751 : OAI21_X1 port map( B1 => n718, B2 => n1454, A => n1439, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U1752 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => 
                           n1440);
   U1753 : OAI21_X1 port map( B1 => n719, B2 => n1454, A => n1440, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U1754 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => 
                           n1441);
   U1755 : OAI21_X1 port map( B1 => n720, B2 => n1454, A => n1441, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U1756 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n1442, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => 
                           n1443);
   U1757 : OAI21_X1 port map( B1 => n721, B2 => n1454, A => n1443, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U1758 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => 
                           n1444);
   U1759 : OAI21_X1 port map( B1 => n722, B2 => n1454, A => n1444, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U1760 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => 
                           n1445);
   U1761 : OAI21_X1 port map( B1 => n723, B2 => n1454, A => n1445, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U1762 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => 
                           n1446);
   U1763 : OAI21_X1 port map( B1 => n691, B2 => n1454, A => n1446, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U1764 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => 
                           n1447);
   U1765 : OAI21_X1 port map( B1 => n724, B2 => n1454, A => n1447, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U1766 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => 
                           n1448);
   U1767 : OAI21_X1 port map( B1 => n725, B2 => n1454, A => n1448, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U1768 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => 
                           n1449);
   U1769 : OAI21_X1 port map( B1 => n726, B2 => n1454, A => n1449, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U1770 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => 
                           n1450);
   U1771 : OAI21_X1 port map( B1 => n727, B2 => n1454, A => n1450, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U1772 : AOI22_X1 port map( A1 => n1452, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n1451, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => 
                           n1453);
   U1773 : OAI21_X1 port map( B1 => n703, B2 => n1454, A => n1453, ZN => 
                           datapath_i_decode_stage_dp_n12);
   U1774 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n1456, A => n1455, ZN => cu_i_cmd_word_6_port);
   U1775 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_6_port, B1 => 
                           cu_i_cw1_10_port, B2 => n1535, ZN => n1470);
   U1776 : NOR4_X1 port map( A1 => datapath_i_val_a_i_14_port, A2 => 
                           datapath_i_val_a_i_15_port, A3 => 
                           datapath_i_val_a_i_16_port, A4 => 
                           datapath_i_val_a_i_17_port, ZN => n1460);
   U1777 : NOR4_X1 port map( A1 => datapath_i_val_a_i_18_port, A2 => 
                           datapath_i_val_a_i_19_port, A3 => 
                           datapath_i_val_a_i_20_port, A4 => 
                           datapath_i_val_a_i_21_port, ZN => n1459);
   U1778 : NOR4_X1 port map( A1 => datapath_i_val_a_i_26_port, A2 => 
                           datapath_i_val_a_i_7_port, A3 => 
                           datapath_i_val_a_i_8_port, A4 => 
                           datapath_i_val_a_i_9_port, ZN => n1458);
   U1779 : NOR4_X1 port map( A1 => datapath_i_val_a_i_10_port, A2 => 
                           datapath_i_val_a_i_11_port, A3 => 
                           datapath_i_val_a_i_12_port, A4 => 
                           datapath_i_val_a_i_13_port, ZN => n1457);
   U1780 : NAND4_X1 port map( A1 => n1460, A2 => n1459, A3 => n1458, A4 => 
                           n1457, ZN => n1466);
   U1781 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n1464);
   U1782 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n1463);
   U1783 : NOR4_X1 port map( A1 => datapath_i_val_a_i_22_port, A2 => 
                           datapath_i_val_a_i_23_port, A3 => 
                           datapath_i_val_a_i_24_port, A4 => 
                           datapath_i_val_a_i_25_port, ZN => n1462);
   U1784 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n1461);
   U1785 : NAND4_X1 port map( A1 => n1464, A2 => n1463, A3 => n1462, A4 => 
                           n1461, ZN => n1465);
   U1786 : NOR2_X1 port map( A1 => n1466, A2 => n1465, ZN => n1468);
   U1787 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_7_port, B1 => 
                           cu_i_cw1_11_port, B2 => n1535, ZN => n1467);
   U1788 : NAND2_X1 port map( A1 => n1468, A2 => n1467, ZN => n1469);
   U1789 : OAI22_X1 port map( A1 => n1470, A2 => n1469, B1 => n1468, B2 => 
                           n1467, ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U1790 : NOR2_X1 port map( A1 => n1472, A2 => n1471, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U1791 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U1792 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U1793 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U1794 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U1795 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U1796 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U1797 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U1798 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U1799 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
                           ZN => n1473);
   U1800 : NAND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
                           A2 => n310, ZN => n1483);
   U1801 : OAI21_X1 port map( B1 => n310, B2 => n1473, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U1802 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
                           ZN => n1474);
   U1803 : OAI21_X1 port map( B1 => n310, B2 => n1474, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U1804 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
                           ZN => n1475);
   U1805 : OAI21_X1 port map( B1 => n310, B2 => n1475, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U1806 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
                           ZN => n1476);
   U1807 : OAI21_X1 port map( B1 => n1545, B2 => n1476, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U1808 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
                           ZN => n1477);
   U1809 : OAI21_X1 port map( B1 => n310, B2 => n1477, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U1810 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
                           ZN => n1478);
   U1811 : OAI21_X1 port map( B1 => n1545, B2 => n1478, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U1812 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
                           ZN => n1479);
   U1813 : OAI21_X1 port map( B1 => n310, B2 => n1479, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U1814 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
                           ZN => n1480);
   U1815 : OAI21_X1 port map( B1 => n1545, B2 => n1480, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U1816 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
                           ZN => n1481);
   U1817 : OAI21_X1 port map( B1 => n1545, B2 => n1481, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U1818 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
                           ZN => n1482);
   U1819 : OAI21_X1 port map( B1 => n310, B2 => n1482, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U1820 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, S 
                           => n310, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U1821 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
                           ZN => n1484);
   U1822 : OAI21_X1 port map( B1 => n310, B2 => n1484, A => n1483, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U1823 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, S 
                           => n310, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U1824 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U1825 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U1826 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U1827 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U1828 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, S 
                           => n1545, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U1829 : MUX2_X1 port map( A => datapath_i_val_b_i_7_port, B => 
                           datapath_i_val_immediate_i_7_port, S => n1485, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U1830 : MUX2_X1 port map( A => datapath_i_val_b_i_8_port, B => 
                           datapath_i_val_immediate_i_8_port, S => n1485, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U1831 : MUX2_X1 port map( A => datapath_i_val_b_i_9_port, B => 
                           datapath_i_val_immediate_i_9_port, S => n1485, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U1832 : MUX2_X1 port map( A => datapath_i_val_b_i_10_port, B => 
                           datapath_i_val_immediate_i_10_port, S => n1485, Z =>
                           datapath_i_execute_stage_dp_opb_10_port);
   U1833 : MUX2_X1 port map( A => datapath_i_val_b_i_11_port, B => 
                           datapath_i_val_immediate_i_11_port, S => n1485, Z =>
                           datapath_i_execute_stage_dp_opb_11_port);
   U1834 : MUX2_X1 port map( A => datapath_i_val_b_i_12_port, B => 
                           datapath_i_val_immediate_i_12_port, S => n1485, Z =>
                           datapath_i_execute_stage_dp_opb_12_port);
   U1835 : MUX2_X1 port map( A => datapath_i_val_b_i_13_port, B => 
                           datapath_i_val_immediate_i_13_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_13_port);
   U1836 : MUX2_X1 port map( A => datapath_i_val_b_i_14_port, B => 
                           datapath_i_val_immediate_i_14_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_14_port);
   U1837 : MUX2_X1 port map( A => datapath_i_val_b_i_15_port, B => 
                           datapath_i_val_immediate_i_15_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_15_port);
   U1838 : MUX2_X1 port map( A => datapath_i_val_b_i_16_port, B => 
                           datapath_i_val_immediate_i_16_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_16_port);
   U1839 : MUX2_X1 port map( A => datapath_i_val_b_i_17_port, B => 
                           datapath_i_val_immediate_i_17_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_17_port);
   U1840 : MUX2_X1 port map( A => datapath_i_val_b_i_18_port, B => 
                           datapath_i_val_immediate_i_18_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_18_port);
   U1841 : MUX2_X1 port map( A => datapath_i_val_b_i_19_port, B => 
                           datapath_i_val_immediate_i_19_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_19_port);
   U1842 : MUX2_X1 port map( A => datapath_i_val_b_i_20_port, B => 
                           datapath_i_val_immediate_i_20_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_20_port);
   U1843 : MUX2_X1 port map( A => datapath_i_val_b_i_21_port, B => 
                           datapath_i_val_immediate_i_21_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_21_port);
   U1844 : MUX2_X1 port map( A => datapath_i_val_b_i_22_port, B => 
                           datapath_i_val_immediate_i_22_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_22_port);
   U1845 : MUX2_X1 port map( A => datapath_i_val_b_i_23_port, B => 
                           datapath_i_val_immediate_i_23_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_23_port);
   U1846 : MUX2_X1 port map( A => datapath_i_val_b_i_24_port, B => 
                           datapath_i_val_immediate_i_24_port, S => n1487, Z =>
                           datapath_i_execute_stage_dp_opb_24_port);
   U1847 : NAND2_X1 port map( A1 => n1485, A2 => 
                           datapath_i_val_immediate_i_25_port, ZN => n1486);
   U1848 : OAI21_X1 port map( B1 => n1485, B2 => n758, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U1849 : OAI21_X1 port map( B1 => n1487, B2 => n759, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U1850 : OAI21_X1 port map( B1 => n1485, B2 => n760, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U1851 : OAI21_X1 port map( B1 => n1485, B2 => n761, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U1852 : OAI21_X1 port map( B1 => n1485, B2 => n762, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U1853 : OAI21_X1 port map( B1 => n1485, B2 => n763, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U1854 : OAI21_X1 port map( B1 => n1487, B2 => n764, A => n1486, ZN => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U1855 : MUX2_X1 port map( A => datapath_i_val_immediate_i_1_port, B => 
                           datapath_i_val_b_i_1_port, S => n1488, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U1856 : MUX2_X1 port map( A => datapath_i_val_immediate_i_4_port, B => 
                           datapath_i_val_b_i_4_port, S => n1488, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U1857 : MUX2_X1 port map( A => datapath_i_val_immediate_i_5_port, B => 
                           datapath_i_val_b_i_5_port, S => n1488, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U1858 : MUX2_X1 port map( A => datapath_i_val_immediate_i_6_port, B => 
                           datapath_i_val_b_i_6_port, S => n1488, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U1859 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_7_port, B2 => 
                           n1510, ZN => n1489);
   U1860 : OAI21_X1 port map( B1 => n705, B2 => n1525, A => n1489, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U1861 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_8_port, B2 => 
                           n1522, ZN => n1490);
   U1862 : OAI21_X1 port map( B1 => n706, B2 => n1514, A => n1490, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U1863 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_9_port, B2 => 
                           n1510, ZN => n1491);
   U1864 : OAI21_X1 port map( B1 => n707, B2 => n1525, A => n1491, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U1865 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n1522, ZN => n1492);
   U1866 : OAI21_X1 port map( B1 => n708, B2 => n1514, A => n1492, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U1867 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n1510, ZN => n1493);
   U1868 : OAI21_X1 port map( B1 => n709, B2 => n1525, A => n1493, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U1869 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n1522, ZN => n1494);
   U1870 : OAI21_X1 port map( B1 => n710, B2 => n1514, A => n1494, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U1871 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n1510, ZN => n1495);
   U1872 : OAI21_X1 port map( B1 => n711, B2 => n1525, A => n1495, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U1873 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n1522, ZN => n1496);
   U1874 : OAI21_X1 port map( B1 => n712, B2 => n1514, A => n1496, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U1875 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n1510, ZN => n1497);
   U1876 : OAI21_X1 port map( B1 => n713, B2 => n1525, A => n1497, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U1877 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n1510, ZN => n1498);
   U1878 : OAI21_X1 port map( B1 => n714, B2 => n1525, A => n1498, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U1879 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n1522, ZN => n1499);
   U1880 : OAI21_X1 port map( B1 => n715, B2 => n1525, A => n1499, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U1881 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n1510, ZN => n1500);
   U1882 : OAI21_X1 port map( B1 => n716, B2 => n1514, A => n1500, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U1883 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n1522, ZN => n1501);
   U1884 : OAI21_X1 port map( B1 => n717, B2 => n1514, A => n1501, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U1885 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n1510, ZN => n1502);
   U1886 : OAI21_X1 port map( B1 => n718, B2 => n1514, A => n1502, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U1887 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n1522, ZN => n1503);
   U1888 : OAI21_X1 port map( B1 => n719, B2 => n1514, A => n1503, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U1889 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n1510, ZN => n1504);
   U1890 : OAI21_X1 port map( B1 => n720, B2 => n1514, A => n1504, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U1891 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n1510, ZN => n1505);
   U1892 : OAI21_X1 port map( B1 => n721, B2 => n1514, A => n1505, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U1893 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n1510, ZN => n1506);
   U1894 : OAI21_X1 port map( B1 => n722, B2 => n1514, A => n1506, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U1895 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n1510, ZN => n1507);
   U1896 : OAI21_X1 port map( B1 => n723, B2 => n1514, A => n1507, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U1897 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_0_port, B2 => 
                           n1510, ZN => n1508);
   U1898 : OAI21_X1 port map( B1 => n733, B2 => n1514, A => n1508, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U1899 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n1510, ZN => n1509);
   U1900 : OAI21_X1 port map( B1 => n724, B2 => n1514, A => n1509, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U1901 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n1510, ZN => n1511);
   U1902 : OAI21_X1 port map( B1 => n725, B2 => n1514, A => n1511, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U1903 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n1512, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n1522, ZN => n1513);
   U1904 : OAI21_X1 port map( B1 => n726, B2 => n1514, A => n1513, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U1905 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n1522, ZN => n1515);
   U1906 : OAI21_X1 port map( B1 => n727, B2 => n1525, A => n1515, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U1907 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n1522, ZN => n1516);
   U1908 : OAI21_X1 port map( B1 => n703, B2 => n1525, A => n1516, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U1909 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_1_port, B2 => 
                           n1522, ZN => n1517);
   U1910 : OAI21_X1 port map( B1 => n734, B2 => n1525, A => n1517, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U1911 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_2_port, B2 => 
                           n1522, ZN => n1518);
   U1912 : OAI21_X1 port map( B1 => n728, B2 => n1525, A => n1518, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U1913 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_3_port, B2 => 
                           n1522, ZN => n1519);
   U1914 : OAI21_X1 port map( B1 => n729, B2 => n1525, A => n1519, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U1915 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_4_port, B2 => 
                           n1522, ZN => n1520);
   U1916 : OAI21_X1 port map( B1 => n730, B2 => n1525, A => n1520, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U1917 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_5_port, B2 => 
                           n1522, ZN => n1521);
   U1918 : OAI21_X1 port map( B1 => n731, B2 => n1525, A => n1521, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U1919 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n1523, B1 => datapath_i_val_a_i_6_port, B2 => 
                           n1522, ZN => n1524);
   U1920 : OAI21_X1 port map( B1 => n732, B2 => n1525, A => n1524, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);

end SYN_dlx_rtl;
