
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n3076, 
      n3077, n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n1995, n1996, 
      n1997, n5121, n5122, n5123, n5124, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n1991, n1992, n7164, n7165, n1993, n1994, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n9196, n9197, n9198, 
      n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, 
      n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, 
      n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, 
      n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, 
      n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, 
      n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, 
      n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, 
      n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, 
      n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, 
      n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, 
      n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, 
      n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, 
      n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, 
      n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, 
      n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, 
      n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, 
      n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, 
      n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, 
      n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, 
      n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, 
      n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, 
      n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, 
      n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, 
      n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, 
      n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, 
      n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, 
      n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, 
      n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, 
      n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, 
      n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, 
      n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, 
      n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, 
      n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, 
      n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, 
      n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, 
      n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, 
      n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, 
      n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, 
      n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, 
      n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, 
      n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, 
      n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, 
      n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, 
      n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, 
      n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, 
      n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, 
      n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, 
      n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, 
      n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, 
      n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, 
      n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, 
      n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, 
      n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, 
      n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, 
      n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, 
      n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, 
      n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, 
      n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, 
      n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, 
      n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, 
      n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, 
      n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, 
      n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, 
      n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, 
      n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, 
      n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, 
      n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, 
      n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, 
      n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, 
      n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, 
      n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, 
      n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, 
      n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, 
      n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, 
      n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, 
      n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, 
      n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, 
      n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, 
      n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, 
      n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, 
      n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, 
      n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, 
      n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, 
      n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, 
      n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, 
      n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, 
      n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, 
      n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, 
      n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, 
      n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, 
      n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, 
      n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, 
      n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, 
      n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, 
      n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, 
      n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, 
      n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, 
      n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, 
      n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, 
      n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, 
      n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, 
      n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, 
      n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, 
      n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, 
      n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, 
      n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, 
      n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, 
      n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, 
      n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, 
      n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, 
      n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, 
      n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, 
      n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, 
      n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, 
      n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, 
      n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, 
      n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, 
      n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, 
      n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, 
      n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, 
      n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, 
      n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, 
      n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, 
      n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, 
      n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, 
      n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, 
      n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, 
      n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, 
      n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, 
      n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, 
      n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, 
      n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, 
      n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, 
      n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, 
      n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, 
      n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, 
      n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, 
      n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, 
      n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, 
      n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, 
      n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, 
      n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, 
      n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, 
      n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, 
      n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, 
      n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, 
      n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, 
      n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, 
      n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, 
      n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, 
      n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, 
      n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, 
      n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, 
      n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, 
      n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, 
      n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, 
      n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, 
      n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, 
      n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, 
      n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, 
      n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, 
      n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, 
      n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, 
      n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, 
      n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, 
      n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, 
      n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, 
      n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, 
      n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, 
      n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, 
      n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, 
      n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, 
      n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, 
      n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, 
      n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, 
      n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, 
      n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, 
      n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, 
      n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, 
      n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, 
      n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, 
      n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, 
      n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, 
      n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, 
      n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, 
      n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, 
      n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, 
      n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, 
      n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, 
      n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, 
      n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, 
      n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, 
      n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, 
      n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, 
      n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, 
      n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, 
      n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, 
      n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, 
      n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, 
      n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, 
      n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, 
      n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, 
      n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, 
      n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, 
      n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, 
      n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, 
      n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, 
      n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, 
      n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, 
      n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, 
      n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, 
      n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, 
      n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, 
      n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, 
      n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, 
      n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, 
      n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n_1004, 
      n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, 
      n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, 
      n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, 
      n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, 
      n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, 
      n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, 
      n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, 
      n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, 
      n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, 
      n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, 
      n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, 
      n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, 
      n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, 
      n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, 
      n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348 : std_logic;

begin
   
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n11230, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n1992, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n11230, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n1992, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n1992, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n1992, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n1992, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n11230, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n11230, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n1992, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n1992, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n1992, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n1992, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n11230, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n1992, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n11230, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n11230, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n1992, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n1992, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n11230, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n11230, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n1992, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n11230, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n11230, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n11230, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n1992, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n1992, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => n11229, GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => n11228, GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => n11227, GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => n9204, Q => n11226, QN => n7165);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => n9201, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => n9196, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => n9207, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => n9199, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3080);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => n9199, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => n9205, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => n9199, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => n9209, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3079);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => n9196, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => n9210, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => n9208, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => n9203, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3078);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => n9203, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => n9205, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => n9204, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => n9207, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => n9210, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => n9202, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => n9201, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => n9208, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3082);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => n9204, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => n9196, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => n9205, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => n9206, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => n9203, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => n9207, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => n9201, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => n9200, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => n9196, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => n9204, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3076);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => n9199, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => n9205, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => n9197, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => n9202, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => n9199, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => n9201, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => n9210, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => n9210, Q => n_1060, QN => n5126);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => n9205, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3095, CK => clk, RN => n9210, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => n9205, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => n9206, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => n9210, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => n9208, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => n9201, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => n9197, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => n9199, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => n9202, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => n9197, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => n9206, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => n9202, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n9203, Q => n_1106, QN => n5134);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => n9210, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => n9197, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => n9207, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => n9209, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => n9197, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => n9210, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => n9207, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => n9199, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => n9202, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1120);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => n9200, Q => n_1121, QN => n5133);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => n9204, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1122
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3094, CK => clk, RN => n9198, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1123
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => n9206, Q => boothmul_pipelined_i_sum_out_6_9_port
                           , QN => n_1124);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => n9201, Q => boothmul_pipelined_i_sum_out_6_8_port
                           , QN => n_1125);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => n9199, Q => boothmul_pipelined_i_sum_out_6_7_port
                           , QN => n_1126);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => n9198, Q => boothmul_pipelined_i_sum_out_6_6_port
                           , QN => n_1127);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => n9208, Q => boothmul_pipelined_i_sum_out_6_5_port
                           , QN => n_1128);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => n9206, Q => boothmul_pipelined_i_sum_out_6_4_port
                           , QN => n_1129);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => n9196, Q => boothmul_pipelined_i_sum_out_6_3_port
                           , QN => n_1130);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => n9200, Q => boothmul_pipelined_i_sum_out_6_2_port
                           , QN => n_1131);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => n9207, Q => boothmul_pipelined_i_sum_out_6_1_port
                           , QN => n_1132);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => n9209, Q => boothmul_pipelined_i_sum_out_6_0_port
                           , QN => n_1133);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => n5129
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => n9197, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => n5123
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1156);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1157);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1158);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1159);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1160);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1161);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1162);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1163);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => n9207, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1164);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => n9205, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1165);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => n9199, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1166);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1167);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => n9210, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => n9199, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => n9207, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => n9199, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1177);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => n9202, Q => n_1178, QN => n5132);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => n9207, Q => boothmul_pipelined_i_sum_out_5_9_port
                           , QN => n_1179);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3093, CK => clk, RN => n9206, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1180)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => n9204, Q => boothmul_pipelined_i_sum_out_5_7_port
                           , QN => n_1181);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => n9197, Q => boothmul_pipelined_i_sum_out_5_6_port
                           , QN => n_1182);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => n9207, Q => boothmul_pipelined_i_sum_out_5_5_port
                           , QN => n_1183);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => n9210, Q => boothmul_pipelined_i_sum_out_5_4_port
                           , QN => n_1184);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => n9203, Q => boothmul_pipelined_i_sum_out_5_3_port
                           , QN => n_1185);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => n9197, Q => boothmul_pipelined_i_sum_out_5_2_port
                           , QN => n_1186);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => n9206, Q => boothmul_pipelined_i_sum_out_5_1_port
                           , QN => n_1187);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => n9201, Q => boothmul_pipelined_i_sum_out_5_0_port
                           , QN => n_1188);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => n9197, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => n5128
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1189);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1190);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1191);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => n9197, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n5122);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => n9210, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => n9197, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => n9210, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => n9201, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => n9205, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => n9201, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => n9205, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1231);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1232
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => n9198, Q => n_1233, QN => n5131);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => n9196, Q => boothmul_pipelined_i_sum_out_4_7_port
                           , QN => n_1234);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3092, CK => clk, RN => n9207, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1235)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => n9209, Q => boothmul_pipelined_i_sum_out_4_5_port
                           , QN => n_1236);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => n9206, Q => boothmul_pipelined_i_sum_out_4_4_port
                           , QN => n_1237);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => n9199, Q => boothmul_pipelined_i_sum_out_4_3_port
                           , QN => n_1238);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => n9209, Q => boothmul_pipelined_i_sum_out_4_2_port
                           , QN => n_1239);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => n9196, Q => boothmul_pipelined_i_sum_out_4_1_port
                           , QN => n_1240);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => n9207, Q => boothmul_pipelined_i_sum_out_4_0_port
                           , QN => n_1241);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => n5127
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1242);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1243);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1244);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1245);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1246);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1249);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1250);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1251);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1252);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1253);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1254);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1255);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => n5121
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1256);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1257);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1258);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => n9198, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => n9197, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => n9201, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => n9201, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => n9202, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => n9209, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => n9205, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => n9205, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1282);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => n9205, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1283
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1284
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => n9201, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1285
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => n9205, Q => n_1286, QN => n5124);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => n9199, Q => boothmul_pipelined_i_sum_out_3_5_port
                           , QN => n_1287);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3091, CK => clk, RN => n9209, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1288)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => n9204, Q => boothmul_pipelined_i_sum_out_3_3_port
                           , QN => n_1289);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => n9200, Q => boothmul_pipelined_i_sum_out_3_2_port
                           , QN => n_1290);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => n9197, Q => boothmul_pipelined_i_sum_out_3_1_port
                           , QN => n_1291);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => n9208, Q => boothmul_pipelined_i_sum_out_3_0_port
                           , QN => n_1292);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => n7164
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1293);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1294);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1295);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1296);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1297);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1298);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => n9201, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => n9199, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => n9197, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => n9207, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => n9200, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => n9204, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => n9203, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => n9206, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => n9210, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => n9205, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => n9208, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => n9209, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => n9202, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => n9209, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => n9204, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => n9207, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => n9202, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => n9208, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => n9206, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => n9200, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => n9198, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => n9198, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1332
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => n9202, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1333
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => n9203, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1334
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => n9196, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1335
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => n9209, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1336
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => n9202, Q => n_1337, QN => n5130);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => n9205, Q => boothmul_pipelined_i_sum_out_2_3_port
                           , QN => n_1338);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3086, CK => clk, RN => n9207, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1339)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           n2022, CK => clk, RN => n9210, Q => 
                           boothmul_pipelined_i_sum_out_2_1_port, QN => n_1340)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => n9207, Q => boothmul_pipelined_i_sum_out_2_0_port
                           , QN => n_1341);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => n9196, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n3077);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n1992, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n2023, B => n2024, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n2021, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n2020, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n2018, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n2016, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n2014, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n2012, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n2010, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n2008, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n2006, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n2004, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n2002, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n2000, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1998, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1993, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => n2019, 
                           CI => n3083, CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => n2017, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => n2015, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => n2013, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => n2011, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => n2009, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => n2007, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => n2005, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => n2003, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => n2001, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => n1999, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => n1994, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1342, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3085,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1343, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3084,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n1991, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1344, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3090,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n1997, B => boothmul_pipelined_i_sum_B_in_4_24_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1345, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3089
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n1996, B => boothmul_pipelined_i_sum_B_in_5_26_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1346, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3088
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n1995, B => boothmul_pipelined_i_sum_B_in_6_28_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1347, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3087
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1348, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n11230, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n11230, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n11230, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n11230, Q => 
                           DATA2_I_27_port);
   U3 : CLKBUF_X1 port map( A => n9199, Z => n9196);
   U4 : CLKBUF_X1 port map( A => n9199, Z => n9197);
   U5 : CLKBUF_X1 port map( A => n9199, Z => n9198);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n9199);
   U7 : CLKBUF_X1 port map( A => n9203, Z => n9200);
   U8 : CLKBUF_X1 port map( A => n9196, Z => n9201);
   U9 : CLKBUF_X1 port map( A => n9197, Z => n9202);
   U10 : CLKBUF_X1 port map( A => n9197, Z => n9203);
   U11 : CLKBUF_X1 port map( A => n9197, Z => n9204);
   U12 : CLKBUF_X1 port map( A => n9197, Z => n9205);
   U13 : CLKBUF_X1 port map( A => n9198, Z => n9206);
   U14 : CLKBUF_X1 port map( A => n9198, Z => n9207);
   U15 : CLKBUF_X1 port map( A => n9198, Z => n9208);
   U16 : CLKBUF_X1 port map( A => n9198, Z => n9209);
   U17 : CLKBUF_X1 port map( A => n9198, Z => n9210);
   U18 : AOI211_X4 port map( C1 => n10927, C2 => n9468, A => n10926, B => 
                           n10925, ZN => n10373);
   U19 : NOR2_X2 port map( A1 => DATA2(4), A2 => DATA2(5), ZN => n10839);
   U20 : NOR2_X1 port map( A1 => n9211, A2 => FUNC(2), ZN => n10895);
   U21 : NOR2_X1 port map( A1 => FUNC(1), A2 => FUNC(0), ZN => n9410);
   U22 : INV_X1 port map( A => n9410, ZN => n9211);
   U23 : INV_X1 port map( A => n10895, ZN => n1992);
   U24 : CLKBUF_X1 port map( A => n1992, Z => n11230);
   U25 : CLKBUF_X1 port map( A => DATA1(3), Z => n11227);
   U26 : CLKBUF_X1 port map( A => DATA1(15), Z => n11229);
   U27 : CLKBUF_X1 port map( A => DATA1(11), Z => n11228);
   U28 : INV_X1 port map( A => data2_mul_1_port, ZN => n9212);
   U29 : NOR2_X1 port map( A1 => boothmul_pipelined_i_encoder_out_0_0_port, A2 
                           => n9212, ZN => n9226);
   U30 : CLKBUF_X1 port map( A => n9226, Z => n11202);
   U31 : NAND2_X1 port map( A1 => n9212, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n11205);
   U32 : INV_X1 port map( A => n11205, ZN => n9229);
   U33 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n10932);
   U34 : NOR2_X1 port map( A1 => n9212, A2 => n10932, ZN => n11203);
   U35 : CLKBUF_X1 port map( A => n11203, Z => n9225);
   U36 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, A2
                           => n11202, B1 => data1_mul_14_port, B2 => n9229, C1 
                           => boothmul_pipelined_i_muxes_in_0_103_port, C2 => 
                           n9225, ZN => n9213);
   U37 : INV_X1 port map( A => n9213, ZN => n1994);
   U38 : INV_X1 port map( A => data1_mul_0_port, ZN => n2024);
   U39 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, A2
                           => n11202, B1 => data1_mul_13_port, B2 => n9229, C1 
                           => boothmul_pipelined_i_muxes_in_0_104_port, C2 => 
                           n11203, ZN => n9214);
   U40 : INV_X1 port map( A => n9214, ZN => n1999);
   U41 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, A2
                           => n11202, B1 => data1_mul_11_port, B2 => n9229, C1 
                           => boothmul_pipelined_i_muxes_in_0_106_port, C2 => 
                           n11203, ZN => n9215);
   U42 : INV_X1 port map( A => n9215, ZN => n2003);
   U43 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, A2
                           => n11202, B1 => data1_mul_12_port, B2 => n9229, C1 
                           => boothmul_pipelined_i_muxes_in_0_105_port, C2 => 
                           n9225, ZN => n9216);
   U44 : INV_X1 port map( A => n9216, ZN => n2001);
   U45 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, A2
                           => n9226, B1 => data1_mul_9_port, B2 => n9229, C1 =>
                           boothmul_pipelined_i_muxes_in_0_108_port, C2 => 
                           n9225, ZN => n9217);
   U46 : INV_X1 port map( A => n9217, ZN => n2007);
   U47 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, A2
                           => n9226, B1 => data1_mul_10_port, B2 => n9229, C1 
                           => boothmul_pipelined_i_muxes_in_0_107_port, C2 => 
                           n9225, ZN => n9218);
   U48 : INV_X1 port map( A => n9218, ZN => n2005);
   U49 : AOI222_X1 port map( A1 => data1_mul_0_port, A2 => n11202, B1 => 
                           data1_mul_1_port, B2 => n9229, C1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C2 => 
                           n9225, ZN => n9219);
   U50 : INV_X1 port map( A => n9219, ZN => n2022);
   U51 : AOI222_X1 port map( A1 => n11202, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           data1_mul_3_port, B2 => n9229, C1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, C2 => 
                           n11203, ZN => n9220);
   U52 : INV_X1 port map( A => n9220, ZN => n2019);
   U53 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, A2
                           => n9226, B1 => data1_mul_4_port, B2 => n9229, C1 =>
                           boothmul_pipelined_i_muxes_in_0_113_port, C2 => 
                           n11203, ZN => n9221);
   U54 : INV_X1 port map( A => n9221, ZN => n2017);
   U55 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, A2
                           => n9226, B1 => data1_mul_5_port, B2 => n9229, C1 =>
                           boothmul_pipelined_i_muxes_in_0_112_port, C2 => 
                           n9225, ZN => n9222);
   U56 : INV_X1 port map( A => n9222, ZN => n2015);
   U57 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, A2
                           => n9226, B1 => data1_mul_6_port, B2 => n9229, C1 =>
                           boothmul_pipelined_i_muxes_in_0_111_port, C2 => 
                           n9225, ZN => n9223);
   U58 : INV_X1 port map( A => n9223, ZN => n2013);
   U59 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, A2
                           => n9226, B1 => data1_mul_7_port, B2 => n9229, C1 =>
                           boothmul_pipelined_i_muxes_in_0_110_port, C2 => 
                           n11203, ZN => n9224);
   U60 : INV_X1 port map( A => n9224, ZN => n2011);
   U61 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, A2
                           => n9226, B1 => data1_mul_8_port, B2 => n9229, C1 =>
                           boothmul_pipelined_i_muxes_in_0_109_port, C2 => 
                           n9225, ZN => n9227);
   U62 : INV_X1 port map( A => n9227, ZN => n2009);
   U63 : INV_X1 port map( A => data1_mul_14_port, ZN => n1998);
   U64 : INV_X1 port map( A => data1_mul_15_port, ZN => n1993);
   U65 : INV_X1 port map( A => data1_mul_13_port, ZN => n2000);
   U66 : INV_X1 port map( A => data1_mul_12_port, ZN => n2002);
   U67 : INV_X1 port map( A => data1_mul_11_port, ZN => n2004);
   U68 : INV_X1 port map( A => data1_mul_10_port, ZN => n2006);
   U69 : INV_X1 port map( A => data1_mul_9_port, ZN => n2008);
   U70 : INV_X1 port map( A => data1_mul_8_port, ZN => n2010);
   U71 : INV_X1 port map( A => data1_mul_7_port, ZN => n2012);
   U72 : INV_X1 port map( A => data1_mul_6_port, ZN => n2014);
   U73 : INV_X1 port map( A => data1_mul_1_port, ZN => n2023);
   U74 : INV_X1 port map( A => data1_mul_2_port, ZN => n2021);
   U75 : INV_X1 port map( A => data1_mul_3_port, ZN => n2020);
   U76 : INV_X1 port map( A => data1_mul_4_port, ZN => n2018);
   U77 : INV_X1 port map( A => data1_mul_5_port, ZN => n2016);
   U78 : XOR2_X1 port map( A => n1993, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => boothmul_pipelined_i_muxes_in_0_119_port);
   U79 : AOI22_X1 port map( A1 => n11203, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n11202, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n9228);
   U80 : OAI21_X1 port map( B1 => n11205, B2 => n1993, A => n9228, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U81 : AOI222_X1 port map( A1 => n9229, A2 => data1_mul_2_port, B1 => n11203,
                           B2 => boothmul_pipelined_i_muxes_in_0_115_port, C1 
                           => n11202, C2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n9231);
   U82 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n10973);
   U83 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n10973, ZN => n10933);
   U84 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n10933, ZN => n9230);
   U85 : NOR2_X1 port map( A1 => n9231, A2 => n9230, ZN => n3083);
   U86 : AOI21_X1 port map( B1 => n9231, B2 => n9230, A => n3083, ZN => n3086);
   U87 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n9232);
   U88 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n9232, ZN => n10975);
   U89 : NOR3_X1 port map( A1 => n5130, A2 => n10975, A3 => n2024, ZN => n3085)
                           ;
   U90 : OR2_X1 port map( A1 => n2024, A2 => n10975, ZN => n9233);
   U91 : AOI21_X1 port map( B1 => n5130, B2 => n9233, A => n3085, ZN => n3091);
   U92 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n9234);
   U93 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, A
                           => n9234, ZN => n11016);
   U94 : NOR3_X1 port map( A1 => n3077, A2 => n5124, A3 => n11016, ZN => n3084)
                           ;
   U95 : AOI221_X1 port map( B1 => n3077, B2 => n5124, C1 => n11016, C2 => 
                           n5124, A => n3084, ZN => n3092);
   U96 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n9235);
   U97 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, A
                           => n9235, ZN => n11052);
   U98 : NOR3_X1 port map( A1 => n5121, A2 => n5131, A3 => n11052, ZN => n3090)
                           ;
   U99 : AOI221_X1 port map( B1 => n5121, B2 => n5131, C1 => n11052, C2 => 
                           n5131, A => n3090, ZN => n3093);
   U100 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n9236);
   U101 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, A
                           => n9236, ZN => n11088);
   U102 : NOR3_X1 port map( A1 => n5122, A2 => n5132, A3 => n11088, ZN => n3089
                           );
   U103 : AOI221_X1 port map( B1 => n5122, B2 => n5132, C1 => n11088, C2 => 
                           n5132, A => n3089, ZN => n3094);
   U104 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n9237);
   U105 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           A => n9237, ZN => n11124);
   U106 : NOR3_X1 port map( A1 => n5123, A2 => n5133, A3 => n11124, ZN => n3088
                           );
   U107 : AOI221_X1 port map( B1 => n5123, B2 => n5133, C1 => n11124, C2 => 
                           n5133, A => n3088, ZN => n3095);
   U108 : INV_X1 port map( A => FUNC(3), ZN => n10894);
   U109 : NAND3_X1 port map( A1 => FUNC(2), A2 => n9410, A3 => n10894, ZN => 
                           n553);
   U110 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(4), ZN => n9378);
   U111 : INV_X1 port map( A => n9378, ZN => n9423);
   U112 : INV_X1 port map( A => DATA2(3), ZN => n10926);
   U113 : NOR2_X1 port map( A1 => n10926, A2 => n10839, ZN => n10797);
   U114 : NOR2_X1 port map( A1 => n9423, A2 => n10797, ZN => n10133);
   U115 : CLKBUF_X1 port map( A => n10133, Z => n10072);
   U116 : NAND2_X1 port map( A1 => DATA2(0), A2 => DATA2(1), ZN => n9339);
   U117 : INV_X1 port map( A => n9339, ZN => n9422);
   U118 : NAND2_X1 port map( A1 => n10926, A2 => n10839, ZN => n9248);
   U119 : NOR2_X1 port map( A1 => n9248, A2 => DATA2(2), ZN => n10109);
   U120 : NAND2_X1 port map( A1 => n9422, A2 => n10109, ZN => n10179);
   U121 : INV_X1 port map( A => n10179, ZN => n9697);
   U122 : CLKBUF_X1 port map( A => n9697, Z => n9715);
   U123 : CLKBUF_X1 port map( A => n10109, Z => n9800);
   U124 : INV_X1 port map( A => n9800, ZN => n9868);
   U125 : AOI22_X1 port map( A1 => DATA1(20), A2 => n9715, B1 => DATA1(21), B2 
                           => n9868, ZN => n9238);
   U126 : INV_X1 port map( A => DATA2(1), ZN => n10928);
   U127 : NOR2_X1 port map( A1 => n10928, A2 => DATA2(0), ZN => n9375);
   U128 : NAND2_X1 port map( A1 => n9800, A2 => n9375, ZN => n10162);
   U129 : INV_X1 port map( A => n10162, ZN => n10183);
   U130 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(19), ZN => n9685);
   U131 : NAND2_X1 port map( A1 => DATA2(0), A2 => n10928, ZN => n10036);
   U132 : INV_X1 port map( A => n9800, ZN => n9853);
   U133 : OR2_X1 port map( A1 => n10036, A2 => n9853, ZN => n10333);
   U134 : INV_X1 port map( A => n10333, ZN => n10803);
   U135 : NAND2_X1 port map( A1 => n10803, A2 => DATA1(18), ZN => n9655);
   U136 : NOR2_X1 port map( A1 => DATA2(0), A2 => DATA2(1), ZN => n9468);
   U137 : NAND2_X1 port map( A1 => n9468, A2 => n10109, ZN => n9837);
   U138 : INV_X1 port map( A => n9837, ZN => n10344);
   U139 : CLKBUF_X1 port map( A => n10344, Z => n10802);
   U140 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(17), ZN => n9672);
   U141 : NAND4_X1 port map( A1 => n9238, A2 => n9685, A3 => n9655, A4 => n9672
                           , ZN => n9247);
   U142 : INV_X1 port map( A => DATA2(2), ZN => n10927);
   U143 : NOR3_X1 port map( A1 => n10927, A2 => n10036, A3 => n9248, ZN => 
                           n10211);
   U144 : INV_X1 port map( A => n10211, ZN => n9943);
   U145 : INV_X1 port map( A => n9943, ZN => n10812);
   U146 : AOI22_X1 port map( A1 => DATA1(18), A2 => n10344, B1 => DATA1(22), B2
                           => n9868, ZN => n9240);
   U147 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(20), ZN => n9683);
   U148 : INV_X1 port map( A => DATA1(21), ZN => n10309);
   U149 : NOR2_X1 port map( A1 => n10179, A2 => n10309, ZN => n9708);
   U150 : INV_X1 port map( A => n9708, ZN => n9239);
   U151 : NAND2_X1 port map( A1 => n10803, A2 => DATA1(19), ZN => n9663);
   U152 : NAND4_X1 port map( A1 => n9240, A2 => n9683, A3 => n9239, A4 => n9663
                           , ZN => n9250);
   U153 : OAI21_X1 port map( B1 => n9248, B2 => DATA2(1), A => n9868, ZN => 
                           n9875);
   U154 : CLKBUF_X1 port map( A => n9875, Z => n9947);
   U155 : INV_X1 port map( A => n9947, ZN => n10114);
   U156 : AOI22_X1 port map( A1 => DATA1(16), A2 => n10802, B1 => DATA1(20), B2
                           => n9853, ZN => n9241);
   U157 : NAND2_X1 port map( A1 => n10803, A2 => DATA1(17), ZN => n9658);
   U158 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(19), ZN => n9680);
   U159 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(18), ZN => n9664);
   U160 : NAND4_X1 port map( A1 => n9241, A2 => n9658, A3 => n9680, A4 => n9664
                           , ZN => n9282);
   U161 : INV_X1 port map( A => DATA2(0), ZN => n10929);
   U162 : OAI21_X1 port map( B1 => n10929, B2 => n10927, A => n9875, ZN => 
                           n9945);
   U163 : CLKBUF_X1 port map( A => n9945, Z => n9897);
   U164 : INV_X1 port map( A => n9897, ZN => n10349);
   U165 : AOI222_X1 port map( A1 => n9247, A2 => n10812, B1 => n9250, B2 => 
                           n10114, C1 => n9282, C2 => n10349, ZN => n9242);
   U166 : INV_X1 port map( A => n9242, ZN => n9303);
   U167 : INV_X1 port map( A => n9248, ZN => n9243);
   U168 : AOI21_X1 port map( B1 => n10929, B2 => n9243, A => n9875, ZN => 
                           n10115);
   U169 : INV_X1 port map( A => n10115, ZN => n10056);
   U170 : INV_X1 port map( A => n10056, ZN => n10817);
   U171 : NAND2_X1 port map( A1 => n9243, A2 => n10817, ZN => n10818);
   U172 : INV_X1 port map( A => n10818, ZN => n10061);
   U173 : CLKBUF_X1 port map( A => n10061, Z => n9996);
   U174 : NAND4_X1 port map( A1 => n10927, A2 => DATA2(3), A3 => n10839, A4 => 
                           n9468, ZN => n10814);
   U175 : AOI22_X1 port map( A1 => DATA1(22), A2 => n9697, B1 => DATA1(23), B2 
                           => n9853, ZN => n9244);
   U176 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(21), ZN => n9699);
   U177 : NAND2_X1 port map( A1 => n10803, A2 => DATA1(20), ZN => n9684);
   U178 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(19), ZN => n9654);
   U179 : NAND4_X1 port map( A1 => n9244, A2 => n9699, A3 => n9684, A4 => n9654
                           , ZN => n9253);
   U180 : INV_X1 port map( A => n9875, ZN => n10810);
   U181 : INV_X1 port map( A => n9945, ZN => n10808);
   U182 : AOI222_X1 port map( A1 => n9250, A2 => n10211, B1 => n9253, B2 => 
                           n10810, C1 => n9247, C2 => n10808, ZN => n9294);
   U183 : INV_X1 port map( A => DATA1(16), ZN => n10675);
   U184 : NOR2_X1 port map( A1 => n10333, A2 => n10675, ZN => n9677);
   U185 : INV_X1 port map( A => DATA1(15), ZN => n10475);
   U186 : NAND2_X1 port map( A1 => n9697, A2 => DATA1(18), ZN => n9686);
   U187 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(17), ZN => n9656);
   U188 : OAI211_X1 port map( C1 => n10475, C2 => n9837, A => n9686, B => n9656
                           , ZN => n9245);
   U189 : AOI211_X1 port map( C1 => DATA1(19), C2 => n9868, A => n9677, B => 
                           n9245, ZN => n9246);
   U190 : INV_X1 port map( A => n9246, ZN => n9291);
   U191 : AOI222_X1 port map( A1 => n9282, A2 => n10211, B1 => n9247, B2 => 
                           n10810, C1 => n9291, C2 => n10808, ZN => n9300);
   U192 : OAI22_X1 port map( A1 => n10814, A2 => n9294, B1 => n10115, B2 => 
                           n9300, ZN => n9255);
   U193 : INV_X1 port map( A => n9468, ZN => n9626);
   U194 : OAI21_X1 port map( B1 => DATA2(2), B2 => DATA2(1), A => DATA2(3), ZN 
                           => n9490);
   U195 : NAND2_X1 port map( A1 => n9490, A2 => n10839, ZN => n10825);
   U196 : INV_X1 port map( A => n10825, ZN => n10352);
   U197 : NAND3_X1 port map( A1 => n9626, A2 => n9248, A3 => n10352, ZN => 
                           n10820);
   U198 : AOI22_X1 port map( A1 => DATA1(23), A2 => n9697, B1 => DATA1(24), B2 
                           => n9853, ZN => n9249);
   U199 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(22), ZN => n9711);
   U200 : INV_X1 port map( A => n10333, ZN => n9941);
   U201 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(21), ZN => n9679);
   U202 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(20), ZN => n9662);
   U203 : NAND4_X1 port map( A1 => n9249, A2 => n9711, A3 => n9679, A4 => n9662
                           , ZN => n9258);
   U204 : AOI222_X1 port map( A1 => n9253, A2 => n10211, B1 => n9258, B2 => 
                           n10810, C1 => n9250, C2 => n10808, ZN => n9283);
   U205 : INV_X1 port map( A => DATA1(22), ZN => n10768);
   U206 : NOR2_X1 port map( A1 => n10333, A2 => n10768, ZN => n9695);
   U207 : INV_X1 port map( A => DATA1(25), ZN => n10230);
   U208 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(23), ZN => n9706);
   U209 : NAND2_X1 port map( A1 => n9697, A2 => DATA1(24), ZN => n9734);
   U210 : OAI211_X1 port map( C1 => n9800, C2 => n10230, A => n9706, B => n9734
                           , ZN => n9251);
   U211 : AOI211_X1 port map( C1 => DATA1(21), C2 => n10802, A => n9695, B => 
                           n9251, ZN => n9252);
   U212 : INV_X1 port map( A => n9252, ZN => n9266);
   U213 : AOI222_X1 port map( A1 => n10114, A2 => n9266, B1 => n10808, B2 => 
                           n9253, C1 => n10812, C2 => n9258, ZN => n9271);
   U214 : OAI22_X1 port map( A1 => n10820, A2 => n9283, B1 => n10352, B2 => 
                           n9271, ZN => n9254);
   U215 : AOI211_X1 port map( C1 => n9303, C2 => n9996, A => n9255, B => n9254,
                           ZN => n9337);
   U216 : NAND2_X1 port map( A1 => DATA2(3), A2 => n9422, ZN => n9552);
   U217 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(2), ZN => n9286);
   U218 : NAND3_X1 port map( A1 => n10839, A2 => n9552, A3 => n9286, ZN => 
                           n10826);
   U219 : INV_X1 port map( A => n10839, ZN => n10071);
   U220 : OR3_X1 port map( A1 => DATA2(2), A2 => n9552, A3 => n10071, ZN => 
                           n10831);
   U221 : INV_X1 port map( A => n10831, ZN => n10554);
   U222 : INV_X1 port map( A => n10820, ZN => n10355);
   U223 : CLKBUF_X1 port map( A => n10355, Z => n9997);
   U224 : INV_X1 port map( A => n9271, ZN => n9279);
   U225 : AOI22_X1 port map( A1 => n9997, A2 => n9279, B1 => n10056, B2 => 
                           n9303, ZN => n9261);
   U226 : INV_X1 port map( A => n10814, ZN => n10058);
   U227 : CLKBUF_X1 port map( A => n10058, Z => n10012);
   U228 : INV_X1 port map( A => n9283, ZN => n9259);
   U229 : INV_X1 port map( A => DATA1(23), ZN => n10256);
   U230 : NOR2_X1 port map( A1 => n10333, A2 => n10256, ZN => n9709);
   U231 : INV_X1 port map( A => DATA1(26), ZN => n10778);
   U232 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(22), ZN => n9678);
   U233 : NAND2_X1 port map( A1 => n9697, A2 => DATA1(25), ZN => n9786);
   U234 : OAI211_X1 port map( C1 => n10109, C2 => n10778, A => n9678, B => 
                           n9786, ZN => n9256);
   U235 : AOI211_X1 port map( C1 => DATA1(24), C2 => n10183, A => n9709, B => 
                           n9256, ZN => n9257);
   U236 : INV_X1 port map( A => n9257, ZN => n9268);
   U237 : AOI222_X1 port map( A1 => n10114, A2 => n9268, B1 => n10808, B2 => 
                           n9258, C1 => n10812, C2 => n9266, ZN => n9351);
   U238 : INV_X1 port map( A => n9351, ZN => n9274);
   U239 : AOI22_X1 port map( A1 => n10012, A2 => n9259, B1 => n10825, B2 => 
                           n9274, ZN => n9260);
   U240 : OAI211_X1 port map( C1 => n9294, C2 => n10818, A => n9261, B => n9260
                           , ZN => n9333);
   U241 : OAI21_X1 port map( B1 => n10928, B2 => n9286, A => n10839, ZN => 
                           n10124);
   U242 : CLKBUF_X1 port map( A => n10124, Z => n9924);
   U243 : INV_X1 port map( A => n9924, ZN => n10834);
   U244 : INV_X1 port map( A => DATA1(27), ZN => n10193);
   U245 : NOR2_X1 port map( A1 => n10179, A2 => n10193, ZN => n9834);
   U246 : INV_X1 port map( A => DATA1(28), ZN => n10784);
   U247 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(24), ZN => n9710);
   U248 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(25), ZN => n9716);
   U249 : OAI211_X1 port map( C1 => n9800, C2 => n10784, A => n9710, B => n9716
                           , ZN => n9262);
   U250 : AOI211_X1 port map( C1 => DATA1(26), C2 => n10183, A => n9834, B => 
                           n9262, ZN => n9263);
   U251 : INV_X1 port map( A => n9263, ZN => n9350);
   U252 : AOI22_X1 port map( A1 => DATA1(24), A2 => n10803, B1 => DATA1(27), B2
                           => n9853, ZN => n9264);
   U253 : NAND2_X1 port map( A1 => n9697, A2 => DATA1(26), ZN => n9798);
   U254 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(25), ZN => n9735);
   U255 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(23), ZN => n9698);
   U256 : NAND4_X1 port map( A1 => n9264, A2 => n9798, A3 => n9735, A4 => n9698
                           , ZN => n9267);
   U257 : AOI222_X1 port map( A1 => n10114, A2 => n9350, B1 => n10808, B2 => 
                           n9268, C1 => n10812, C2 => n9267, ZN => n10292);
   U258 : OAI22_X1 port map( A1 => n9351, A2 => n10818, B1 => n10292, B2 => 
                           n10820, ZN => n9270);
   U259 : AOI22_X1 port map( A1 => DATA1(26), A2 => n10803, B1 => DATA1(29), B2
                           => n9853, ZN => n9265);
   U260 : NAND2_X1 port map( A1 => n9697, A2 => DATA1(28), ZN => n9937);
   U261 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(27), ZN => n9799);
   U262 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(25), ZN => n9704);
   U263 : NAND4_X1 port map( A1 => n9265, A2 => n9937, A3 => n9799, A4 => n9704
                           , ZN => n9363);
   U264 : AOI222_X1 port map( A1 => n9350, A2 => n10211, B1 => n9363, B2 => 
                           n10810, C1 => n9267, C2 => n10808, ZN => n10291);
   U265 : AOI222_X1 port map( A1 => n9268, A2 => n10812, B1 => n9267, B2 => 
                           n10810, C1 => n9266, C2 => n10808, ZN => n9364);
   U266 : OAI22_X1 port map( A1 => n10352, A2 => n10291, B1 => n9364, B2 => 
                           n10814, ZN => n9269);
   U267 : AOI211_X1 port map( C1 => n10056, C2 => n9279, A => n9270, B => n9269
                           , ZN => n9361);
   U268 : OAI22_X1 port map( A1 => n10352, A2 => n10292, B1 => n10115, B2 => 
                           n9283, ZN => n9273);
   U269 : OAI22_X1 port map( A1 => n10820, A2 => n9364, B1 => n10818, B2 => 
                           n9271, ZN => n9272);
   U270 : AOI211_X1 port map( C1 => n9274, C2 => n10012, A => n9273, B => n9272
                           , ZN => n9369);
   U271 : NOR3_X1 port map( A1 => n10929, A2 => n9286, A3 => n10124, ZN => 
                           n10414);
   U272 : INV_X1 port map( A => n10414, ZN => n10069);
   U273 : OAI22_X1 port map( A1 => n10834, A2 => n9361, B1 => n9369, B2 => 
                           n10069, ZN => n9275);
   U274 : AOI21_X1 port map( B1 => n10554, B2 => n9333, A => n9275, ZN => n9276
                           );
   U275 : OAI21_X1 port map( B1 => n9337, B2 => n10826, A => n9276, ZN => n9347
                           );
   U276 : CLKBUF_X1 port map( A => n10414, Z => n10838);
   U277 : OAI22_X1 port map( A1 => n10817, A2 => n9294, B1 => n9283, B2 => 
                           n10818, ZN => n9278);
   U278 : OAI22_X1 port map( A1 => n10352, A2 => n9364, B1 => n9351, B2 => 
                           n10820, ZN => n9277);
   U279 : AOI211_X1 port map( C1 => n10012, C2 => n9279, A => n9278, B => n9277
                           , ZN => n9368);
   U280 : INV_X1 port map( A => n9368, ZN => n9358);
   U281 : INV_X1 port map( A => n10826, ZN => n10576);
   U282 : OAI22_X1 port map( A1 => n9300, A2 => n10818, B1 => n9294, B2 => 
                           n10820, ZN => n9285);
   U283 : NOR2_X1 port map( A1 => n10333, A2 => n10475, ZN => n9670);
   U284 : INV_X1 port map( A => DATA1(14), ZN => n10486);
   U285 : NAND2_X1 port map( A1 => n9697, A2 => DATA1(17), ZN => n9665);
   U286 : NAND2_X1 port map( A1 => DATA1(18), A2 => n9853, ZN => n9681);
   U287 : OAI211_X1 port map( C1 => n9837, C2 => n10486, A => n9665, B => n9681
                           , ZN => n9280);
   U288 : AOI211_X1 port map( C1 => DATA1(16), C2 => n10183, A => n9670, B => 
                           n9280, ZN => n9281);
   U289 : INV_X1 port map( A => n9281, ZN => n9299);
   U290 : AOI222_X1 port map( A1 => n9291, A2 => n10812, B1 => n9282, B2 => 
                           n10810, C1 => n9299, C2 => n10808, ZN => n9313);
   U291 : OAI22_X1 port map( A1 => n10352, A2 => n9283, B1 => n10817, B2 => 
                           n9313, ZN => n9284);
   U292 : AOI211_X1 port map( C1 => n10058, C2 => n9303, A => n9285, B => n9284
                           , ZN => n9305);
   U293 : INV_X1 port map( A => n9305, ZN => n9332);
   U294 : AOI22_X1 port map( A1 => n10838, A2 => n9358, B1 => n10576, B2 => 
                           n9332, ZN => n9288);
   U295 : NOR3_X1 port map( A1 => n10071, A2 => n9626, A3 => n9286, ZN => 
                           n10065);
   U296 : INV_X1 port map( A => n10065, ZN => n10828);
   U297 : INV_X1 port map( A => n10828, ZN => n10525);
   U298 : INV_X1 port map( A => n9369, ZN => n10412);
   U299 : AOI22_X1 port map( A1 => n10525, A2 => n9333, B1 => n9924, B2 => 
                           n10412, ZN => n9287);
   U300 : OAI211_X1 port map( C1 => n9337, C2 => n10831, A => n9288, B => n9287
                           , ZN => n9348);
   U301 : OAI21_X1 port map( B1 => n10927, B2 => n9552, A => n10839, ZN => 
                           n10842);
   U302 : CLKBUF_X1 port map( A => n10842, Z => n9813);
   U303 : INV_X1 port map( A => n9813, ZN => n10488);
   U304 : NOR2_X1 port map( A1 => n10071, A2 => n10488, ZN => n10462);
   U305 : CLKBUF_X1 port map( A => n10462, Z => n9927);
   U306 : INV_X1 port map( A => n9333, ZN => n9355);
   U307 : OAI22_X1 port map( A1 => n10834, A2 => n9368, B1 => n9355, B2 => 
                           n10069, ZN => n9296);
   U308 : INV_X1 port map( A => n9300, ZN => n9316);
   U309 : INV_X1 port map( A => n9313, ZN => n9289);
   U310 : AOI22_X1 port map( A1 => n10058, A2 => n9316, B1 => n9996, B2 => 
                           n9289, ZN => n9293);
   U311 : AOI22_X1 port map( A1 => DATA1(16), A2 => n9697, B1 => DATA1(17), B2 
                           => n9853, ZN => n9290);
   U312 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(15), ZN => n9675);
   U313 : NAND2_X1 port map( A1 => DATA1(14), A2 => n9941, ZN => n9751);
   U314 : NAND2_X1 port map( A1 => DATA1(13), A2 => n10802, ZN => n9767);
   U315 : NAND4_X1 port map( A1 => n9290, A2 => n9675, A3 => n9751, A4 => n9767
                           , ZN => n9308);
   U316 : AOI222_X1 port map( A1 => n10114, A2 => n9291, B1 => n10349, B2 => 
                           n9308, C1 => n10812, C2 => n9299, ZN => n9323);
   U317 : INV_X1 port map( A => n9323, ZN => n9312);
   U318 : AOI22_X1 port map( A1 => n10355, A2 => n9303, B1 => n10056, B2 => 
                           n9312, ZN => n9292);
   U319 : OAI211_X1 port map( C1 => n10352, C2 => n9294, A => n9293, B => n9292
                           , ZN => n9334);
   U320 : INV_X1 port map( A => n9334, ZN => n9304);
   U321 : OAI22_X1 port map( A1 => n9304, A2 => n10826, B1 => n9305, B2 => 
                           n10831, ZN => n9295);
   U322 : NOR2_X1 port map( A1 => n9296, A2 => n9295, ZN => n9341);
   U323 : OAI21_X1 port map( B1 => n9337, B2 => n10828, A => n9341, ZN => n9340
                           );
   U324 : AOI222_X1 port map( A1 => n9347, A2 => n10071, B1 => n9348, B2 => 
                           n9927, C1 => n9340, C2 => n10488, ZN => n9360);
   U325 : NOR2_X1 port map( A1 => DATA2(2), A2 => n9626, ZN => n9297);
   U326 : AOI21_X1 port map( B1 => n9297, B2 => n10926, A => n10839, ZN => 
                           n10023);
   U327 : INV_X1 port map( A => n10023, ZN => n10848);
   U328 : AOI22_X1 port map( A1 => DATA1(15), A2 => n9697, B1 => DATA1(16), B2 
                           => n9853, ZN => n9298);
   U329 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(14), ZN => n9667);
   U330 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(13), ZN => n9760);
   U331 : NAND2_X1 port map( A1 => n10802, A2 => DATA1(12), ZN => n9823);
   U332 : NAND4_X1 port map( A1 => n9298, A2 => n9667, A3 => n9760, A4 => n9823
                           , ZN => n9309);
   U333 : AOI222_X1 port map( A1 => n10349, A2 => n9309, B1 => n10810, B2 => 
                           n9299, C1 => n10812, C2 => n9308, ZN => n9431);
   U334 : OAI22_X1 port map( A1 => n10814, A2 => n9313, B1 => n10817, B2 => 
                           n9431, ZN => n9302);
   U335 : OAI22_X1 port map( A1 => n10820, A2 => n9300, B1 => n10818, B2 => 
                           n9323, ZN => n9301);
   U336 : AOI211_X1 port map( C1 => n10825, C2 => n9303, A => n9302, B => n9301
                           , ZN => n9328);
   U337 : OAI22_X1 port map( A1 => n10834, A2 => n9305, B1 => n9304, B2 => 
                           n10069, ZN => n9318);
   U338 : INV_X1 port map( A => DATA1(12), ZN => n10744);
   U339 : NOR2_X1 port map( A1 => n10162, A2 => n10744, ZN => n9762);
   U340 : CLKBUF_X1 port map( A => DATA1(10), Z => n9763);
   U341 : NAND2_X1 port map( A1 => n10802, A2 => n9763, ZN => n9872);
   U342 : NAND2_X1 port map( A1 => DATA1(13), A2 => n9697, ZN => n9668);
   U343 : OAI211_X1 port map( C1 => n9800, C2 => n10486, A => n9872, B => n9668
                           , ZN => n9306);
   U344 : AOI211_X1 port map( C1 => n11228, C2 => n9941, A => n9762, B => n9306
                           , ZN => n9428);
   U345 : INV_X1 port map( A => n9428, ZN => n9320);
   U346 : AOI22_X1 port map( A1 => DATA1(11), A2 => n10344, B1 => DATA1(15), B2
                           => n9853, ZN => n9307);
   U347 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(12), ZN => n9766);
   U348 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(13), ZN => n9750);
   U349 : NAND2_X1 port map( A1 => DATA1(14), A2 => n9715, ZN => n9674);
   U350 : NAND4_X1 port map( A1 => n9307, A2 => n9766, A3 => n9750, A4 => n9674
                           , ZN => n9322);
   U351 : AOI222_X1 port map( A1 => n10114, A2 => n9309, B1 => n10808, B2 => 
                           n9320, C1 => n10812, C2 => n9322, ZN => n9499);
   U352 : AOI222_X1 port map( A1 => n9309, A2 => n10812, B1 => n9308, B2 => 
                           n10810, C1 => n9322, C2 => n10349, ZN => n9475);
   U353 : OAI22_X1 port map( A1 => n9499, A2 => n10817, B1 => n9475, B2 => 
                           n10818, ZN => n9311);
   U354 : OAI22_X1 port map( A1 => n10352, A2 => n9313, B1 => n9431, B2 => 
                           n10814, ZN => n9310);
   U355 : AOI211_X1 port map( C1 => n9997, C2 => n9312, A => n9311, B => n9310,
                           ZN => n9501);
   U356 : OAI22_X1 port map( A1 => n10814, A2 => n9323, B1 => n9475, B2 => 
                           n10115, ZN => n9315);
   U357 : OAI22_X1 port map( A1 => n10820, A2 => n9313, B1 => n10818, B2 => 
                           n9431, ZN => n9314);
   U358 : AOI211_X1 port map( C1 => n10825, C2 => n9316, A => n9315, B => n9314
                           , ZN => n9432);
   U359 : OAI22_X1 port map( A1 => n9501, A2 => n10826, B1 => n9432, B2 => 
                           n10831, ZN => n9317);
   U360 : NOR2_X1 port map( A1 => n9318, A2 => n9317, ZN => n9436);
   U361 : OAI21_X1 port map( B1 => n10828, B2 => n9328, A => n9436, ZN => n9338
                           );
   U362 : INV_X1 port map( A => n9499, ZN => n9472);
   U363 : INV_X1 port map( A => DATA1(11), ZN => n10555);
   U364 : NOR2_X1 port map( A1 => n10162, A2 => n10555, ZN => n9769);
   U365 : INV_X1 port map( A => DATA1(13), ZN => n10511);
   U366 : NAND2_X1 port map( A1 => n10344, A2 => DATA1(9), ZN => n9397);
   U367 : NAND2_X1 port map( A1 => DATA1(12), A2 => n9697, ZN => n9749);
   U368 : OAI211_X1 port map( C1 => n9800, C2 => n10511, A => n9397, B => n9749
                           , ZN => n9319);
   U369 : AOI211_X1 port map( C1 => DATA1(10), C2 => n9941, A => n9769, B => 
                           n9319, ZN => n9471);
   U370 : INV_X1 port map( A => n9471, ZN => n9321);
   U371 : AOI222_X1 port map( A1 => n10114, A2 => n9322, B1 => n10349, B2 => 
                           n9321, C1 => n10812, C2 => n9320, ZN => n9424);
   U372 : OAI22_X1 port map( A1 => n9424, A2 => n10817, B1 => n9475, B2 => 
                           n10814, ZN => n9325);
   U373 : OAI22_X1 port map( A1 => n10352, A2 => n9323, B1 => n9431, B2 => 
                           n10820, ZN => n9324);
   U374 : AOI211_X1 port map( C1 => n10061, C2 => n9472, A => n9325, B => n9324
                           , ZN => n9539);
   U375 : OAI22_X1 port map( A1 => n9539, A2 => n10826, B1 => n9432, B2 => 
                           n10828, ZN => n9327);
   U376 : OAI22_X1 port map( A1 => n9501, A2 => n10831, B1 => n9328, B2 => 
                           n10069, ZN => n9326);
   U377 : AOI211_X1 port map( C1 => n9924, C2 => n9334, A => n9327, B => n9326,
                           ZN => n9479);
   U378 : INV_X1 port map( A => n9479, ZN => n9331);
   U379 : INV_X1 port map( A => n9432, ZN => n9478);
   U380 : AOI22_X1 port map( A1 => n9478, A2 => n10576, B1 => n9334, B2 => 
                           n10525, ZN => n9330);
   U381 : INV_X1 port map( A => n9328, ZN => n9435);
   U382 : AOI22_X1 port map( A1 => n9435, A2 => n10554, B1 => n9332, B2 => 
                           n10838, ZN => n9329);
   U383 : OAI211_X1 port map( C1 => n10834, C2 => n9337, A => n9330, B => n9329
                           , ZN => n9343);
   U384 : AOI222_X1 port map( A1 => n9927, A2 => n9338, B1 => n10488, B2 => 
                           n9331, C1 => n9343, C2 => n10071, ZN => n9507);
   U385 : INV_X1 port map( A => n9507, ZN => n9543);
   U386 : NOR4_X1 port map( A1 => DATA2(2), A2 => DATA2(1), A3 => n10797, A4 =>
                           n10848, ZN => n10852);
   U387 : CLKBUF_X1 port map( A => n10852, Z => n10527);
   U388 : AOI22_X1 port map( A1 => n10525, A2 => n9332, B1 => n10576, B2 => 
                           n9435, ZN => n9336);
   U389 : AOI22_X1 port map( A1 => n10554, A2 => n9334, B1 => n10124, B2 => 
                           n9333, ZN => n9335);
   U390 : OAI211_X1 port map( C1 => n9337, C2 => n10069, A => n9336, B => n9335
                           , ZN => n9344);
   U391 : AOI222_X1 port map( A1 => n9344, A2 => n10071, B1 => n9343, B2 => 
                           n9927, C1 => n9338, C2 => n10488, ZN => n9508);
   U392 : INV_X1 port map( A => n9508, ZN => n9481);
   U393 : AOI22_X1 port map( A1 => n10848, A2 => n9543, B1 => n10527, B2 => 
                           n9481, ZN => n9346);
   U394 : INV_X1 port map( A => DATA2(4), ZN => n10925);
   U395 : INV_X1 port map( A => n10133, ZN => n10849);
   U396 : NOR3_X1 port map( A1 => n10925, A2 => n9339, A3 => n10849, ZN => 
                           n10531);
   U397 : CLKBUF_X1 port map( A => n10531, Z => n10130);
   U398 : AOI222_X1 port map( A1 => n9348, A2 => n10071, B1 => n9340, B2 => 
                           n10462, C1 => n9344, C2 => n10488, ZN => n9438);
   U399 : INV_X1 port map( A => n9438, ZN => n10528);
   U400 : NAND3_X1 port map( A1 => n9375, A2 => n10072, A3 => n10071, ZN => 
                           n10408);
   U401 : INV_X1 port map( A => n10408, ZN => n10846);
   U402 : INV_X1 port map( A => n9341, ZN => n9342);
   U403 : AOI222_X1 port map( A1 => n9927, A2 => n9344, B1 => n10488, B2 => 
                           n9343, C1 => n9342, C2 => n10071, ZN => n9437);
   U404 : INV_X1 port map( A => n9437, ZN => n9480);
   U405 : AOI22_X1 port map( A1 => n10130, A2 => n10528, B1 => n10846, B2 => 
                           n9480, ZN => n9345);
   U406 : OAI211_X1 port map( C1 => n10072, C2 => n9360, A => n9346, B => n9345
                           , ZN => n9548);
   U407 : INV_X1 port map( A => n10797, ZN => n10077);
   U408 : AOI21_X1 port map( B1 => n10077, B2 => n9468, A => n10072, ZN => 
                           n10322);
   U409 : INV_X1 port map( A => n10322, ZN => n10858);
   U410 : INV_X1 port map( A => n10527, ZN => n10431);
   U411 : INV_X1 port map( A => n9927, ZN => n10844);
   U412 : AOI21_X1 port map( B1 => n10525, B2 => n9358, A => n9347, ZN => n9372
                           );
   U413 : INV_X1 port map( A => n9348, ZN => n9359);
   U414 : INV_X1 port map( A => n10291, ZN => n9354);
   U415 : INV_X1 port map( A => DATA1(29), ZN => n10158);
   U416 : NOR2_X1 port map( A1 => n9837, A2 => n10778, ZN => n9713);
   U417 : NOR2_X1 port map( A1 => n10333, A2 => n10193, ZN => n9788);
   U418 : AOI211_X1 port map( C1 => DATA1(30), C2 => n9868, A => n9713, B => 
                           n9788, ZN => n9349);
   U419 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(28), ZN => n9835);
   U420 : OAI211_X1 port map( C1 => n10158, C2 => n10179, A => n9349, B => 
                           n9835, ZN => n10209);
   U421 : AOI222_X1 port map( A1 => n9363, A2 => n10812, B1 => n10209, B2 => 
                           n10810, C1 => n9350, C2 => n10349, ZN => n10294);
   U422 : OAI22_X1 port map( A1 => n10352, A2 => n10294, B1 => n10292, B2 => 
                           n10814, ZN => n9353);
   U423 : OAI22_X1 port map( A1 => n10115, A2 => n9351, B1 => n9364, B2 => 
                           n10818, ZN => n9352);
   U424 : AOI211_X1 port map( C1 => n10355, C2 => n9354, A => n9353, B => n9352
                           , ZN => n10390);
   U425 : OAI22_X1 port map( A1 => n10834, A2 => n10390, B1 => n9355, B2 => 
                           n10826, ZN => n9357);
   U426 : OAI22_X1 port map( A1 => n9369, A2 => n10828, B1 => n9361, B2 => 
                           n10069, ZN => n9356);
   U427 : AOI211_X1 port map( C1 => n10554, C2 => n9358, A => n9357, B => n9356
                           , ZN => n10447);
   U428 : OAI222_X1 port map( A1 => n10844, A2 => n9372, B1 => n9813, B2 => 
                           n9359, C1 => n10447, C2 => n10839, ZN => n10529);
   U429 : INV_X1 port map( A => n9360, ZN => n10526);
   U430 : AOI22_X1 port map( A1 => n10130, A2 => n10529, B1 => n10846, B2 => 
                           n10526, ZN => n9374);
   U431 : INV_X1 port map( A => n9361, ZN => n10411);
   U432 : INV_X1 port map( A => n10294, ZN => n9367);
   U433 : INV_X1 port map( A => DATA1(30), ZN => n10793);
   U434 : NOR2_X1 port map( A1 => n9837, A2 => n10193, ZN => n9737);
   U435 : NOR2_X1 port map( A1 => n10333, A2 => n10784, ZN => n9802);
   U436 : AOI211_X1 port map( C1 => DATA1(31), C2 => n9868, A => n9737, B => 
                           n9802, ZN => n9362);
   U437 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(29), ZN => n9938);
   U438 : OAI211_X1 port map( C1 => n10793, C2 => n10179, A => n9362, B => 
                           n9938, ZN => n10210);
   U439 : AOI222_X1 port map( A1 => n10209, A2 => n10812, B1 => n10210, B2 => 
                           n10810, C1 => n9363, C2 => n10349, ZN => n10293);
   U440 : OAI22_X1 port map( A1 => n10352, A2 => n10293, B1 => n10292, B2 => 
                           n10818, ZN => n9366);
   U441 : OAI22_X1 port map( A1 => n10817, A2 => n9364, B1 => n10291, B2 => 
                           n10814, ZN => n9365);
   U442 : AOI211_X1 port map( C1 => n9997, C2 => n9367, A => n9366, B => n9365,
                           ZN => n10391);
   U443 : OAI22_X1 port map( A1 => n10834, A2 => n10391, B1 => n9368, B2 => 
                           n10826, ZN => n9371);
   U444 : OAI22_X1 port map( A1 => n9369, A2 => n10831, B1 => n10390, B2 => 
                           n10069, ZN => n9370);
   U445 : AOI211_X1 port map( C1 => n10525, C2 => n10411, A => n9371, B => 
                           n9370, ZN => n10446);
   U446 : OAI222_X1 port map( A1 => n10844, A2 => n10447, B1 => n9813, B2 => 
                           n9372, C1 => n10446, C2 => n10839, ZN => n10530);
   U447 : AOI22_X1 port map( A1 => n10848, A2 => n9480, B1 => n10849, B2 => 
                           n10530, ZN => n9373);
   U448 : OAI211_X1 port map( C1 => n9438, C2 => n10431, A => n9374, B => n9373
                           , ZN => n10568);
   U449 : NAND3_X1 port map( A1 => n9423, A2 => n9375, A3 => n10077, ZN => 
                           n10863);
   U450 : INV_X1 port map( A => n10863, ZN => n10365);
   U451 : AOI22_X1 port map( A1 => n10527, A2 => n9480, B1 => n10849, B2 => 
                           n10529, ZN => n9376);
   U452 : OAI21_X1 port map( B1 => n9438, B2 => n10408, A => n9376, ZN => n9377
                           );
   U453 : AOI21_X1 port map( B1 => n10130, B2 => n10526, A => n9377, ZN => 
                           n9492);
   U454 : OAI21_X1 port map( B1 => n9508, B2 => n10023, A => n9492, ZN => 
                           n10567);
   U455 : NOR3_X1 port map( A1 => DATA2(3), A2 => n9378, A3 => n10036, ZN => 
                           n10799);
   U456 : CLKBUF_X1 port map( A => n10799, Z => n10569);
   U457 : AOI222_X1 port map( A1 => n9548, A2 => n10858, B1 => n10568, B2 => 
                           n10365, C1 => n10567, C2 => n10569, ZN => n9421);
   U458 : INV_X1 port map( A => FUNC(0), ZN => n10707);
   U459 : NAND2_X1 port map( A1 => FUNC(1), A2 => n10707, ZN => n9379);
   U460 : NOR2_X1 port map( A1 => DATA2(5), A2 => n9379, ZN => n10051);
   U461 : NAND2_X1 port map( A1 => DATA2(3), A2 => n9423, ZN => n10037);
   U462 : NOR2_X1 port map( A1 => n10037, A2 => n10928, ZN => n10879);
   U463 : NAND2_X1 port map( A1 => DATA2(0), A2 => n10879, ZN => n10053);
   U464 : NAND3_X1 port map( A1 => FUNC(2), A2 => n10051, A3 => n10053, ZN => 
                           n9387);
   U465 : NOR2_X1 port map( A1 => n10894, A2 => n9387, ZN => n10885);
   U466 : CLKBUF_X1 port map( A => n10885, Z => n10482);
   U467 : INV_X1 port map( A => n10482, ZN => n10591);
   U468 : NOR2_X1 port map( A1 => FUNC(2), A2 => n9379, ZN => n10556);
   U469 : INV_X1 port map( A => DATA2(9), ZN => n10918);
   U470 : NAND2_X1 port map( A1 => DATA1(9), A2 => n10918, ZN => n10736);
   U471 : NOR2_X1 port map( A1 => n10918, A2 => DATA1(9), ZN => n10664);
   U472 : INV_X1 port map( A => n10664, ZN => n10731);
   U473 : NAND2_X1 port map( A1 => n10736, A2 => n10731, ZN => n10618);
   U474 : CLKBUF_X1 port map( A => DATA1(8), Z => n10660);
   U475 : NOR2_X1 port map( A1 => n10660, A2 => DATA2_I_8_port, ZN => n9442);
   U476 : XOR2_X1 port map( A => DATA2_I_9_port, B => DATA1(9), Z => n9418);
   U477 : INV_X1 port map( A => n9418, ZN => n9641);
   U478 : NOR2_X1 port map( A1 => n9442, A2 => n9641, ZN => n10588);
   U479 : NAND2_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, ZN => n9385)
                           ;
   U480 : OAI21_X1 port map( B1 => DATA1(7), B2 => DATA2_I_7_port, A => n9385, 
                           ZN => n9488);
   U481 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n9460)
                           ;
   U482 : NAND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n9382)
                           ;
   U483 : INV_X1 port map( A => n9382, ZN => n9456);
   U484 : XOR2_X1 port map( A => DATA2_I_3_port, B => n11227, Z => n9631);
   U485 : NAND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n9453)
                           ;
   U486 : OAI21_X1 port map( B1 => DATA1(2), B2 => DATA2_I_2_port, A => n9453, 
                           ZN => n10151);
   U487 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n9451)
                           ;
   U488 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n10593
                           );
   U489 : INV_X1 port map( A => n10593, ZN => n10337);
   U490 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n10341)
                           ;
   U491 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n9451, 
                           ZN => n10340);
   U492 : NOR2_X1 port map( A1 => n10341, A2 => n10340, ZN => n10339);
   U493 : OAI21_X1 port map( B1 => n10337, B2 => cin, A => n10339, ZN => n9380)
                           ;
   U494 : OAI221_X1 port map( B1 => n10151, B2 => n9451, C1 => n10151, C2 => 
                           n9380, A => n9453, ZN => n9381);
   U495 : AND2_X1 port map( A1 => n11227, A2 => DATA2_I_3_port, ZN => n9454);
   U496 : AOI21_X1 port map( B1 => n9631, B2 => n9381, A => n9454, ZN => n9383)
                           ;
   U497 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n9455)
                           ;
   U498 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n9455, 
                           ZN => n9593);
   U499 : OAI21_X1 port map( B1 => DATA1(5), B2 => DATA2_I_5_port, A => n9382, 
                           ZN => n9555);
   U500 : AOI221_X1 port map( B1 => n9383, B2 => n9455, C1 => n9593, C2 => 
                           n9455, A => n9555, ZN => n9384);
   U501 : XOR2_X1 port map( A => DATA2_I_6_port, B => DATA1(6), Z => n9521);
   U502 : OAI21_X1 port map( B1 => n9456, B2 => n9384, A => n9521, ZN => n9386)
                           ;
   U503 : OAI221_X1 port map( B1 => n9488, B2 => n9460, C1 => n9488, C2 => 
                           n9386, A => n9385, ZN => n10515);
   U504 : NAND2_X1 port map( A1 => n10895, A2 => n10515, ZN => n10565);
   U505 : AOI211_X1 port map( C1 => n9442, C2 => n9641, A => n10588, B => 
                           n10565, ZN => n9416);
   U506 : NOR2_X1 port map( A1 => FUNC(3), A2 => n9387, ZN => n10577);
   U507 : CLKBUF_X1 port map( A => n10577, Z => n10438);
   U508 : INV_X1 port map( A => n10438, ZN => n10559);
   U509 : INV_X1 port map( A => DATA1(3), ZN => n9632);
   U510 : NOR2_X1 port map( A1 => n10333, A2 => n9632, ZN => n9390);
   U511 : INV_X1 port map( A => DATA1(0), ZN => n10645);
   U512 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(2), ZN => n10806);
   U513 : NAND2_X1 port map( A1 => n10344, A2 => DATA1(4), ZN => n9388);
   U514 : OAI211_X1 port map( C1 => n10109, C2 => n10645, A => n10806, B => 
                           n9388, ZN => n9389);
   U515 : AOI211_X1 port map( C1 => n9715, C2 => DATA1(1), A => n9390, B => 
                           n9389, ZN => n9561);
   U516 : INV_X1 port map( A => DATA1(4), ZN => n9562);
   U517 : NOR2_X1 port map( A1 => n10162, A2 => n9562, ZN => n10111);
   U518 : INV_X1 port map( A => DATA1(6), ZN => n10644);
   U519 : NOR2_X1 port map( A1 => n9837, A2 => n10644, ZN => n9391);
   U520 : AOI211_X1 port map( C1 => DATA1(2), C2 => n9868, A => n10111, B => 
                           n9391, ZN => n9392);
   U521 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(5), ZN => n9567);
   U522 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(3), ZN => n10805);
   U523 : AND3_X1 port map( A1 => n9392, A2 => n9567, A3 => n10805, ZN => n9400
                           );
   U524 : INV_X1 port map( A => DATA1(5), ZN => n9527);
   U525 : NOR2_X1 port map( A1 => n9837, A2 => n9527, ZN => n9394);
   U526 : INV_X1 port map( A => DATA1(2), ZN => n10715);
   U527 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(4), ZN => n9607);
   U528 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(3), ZN => n10347);
   U529 : OAI211_X1 port map( C1 => n10179, C2 => n10715, A => n9607, B => 
                           n10347, ZN => n9393);
   U530 : AOI211_X1 port map( C1 => DATA1(1), C2 => n9868, A => n9394, B => 
                           n9393, ZN => n9524);
   U531 : OAI222_X1 port map( A1 => n9947, A2 => n9561, B1 => n9897, B2 => 
                           n9400, C1 => n9943, C2 => n9524, ZN => n10059);
   U532 : INV_X1 port map( A => DATA1(7), ZN => n9462);
   U533 : NOR2_X1 port map( A1 => n9837, A2 => n9462, ZN => n9396);
   U534 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(6), ZN => n9531);
   U535 : NAND2_X1 port map( A1 => n10183, A2 => DATA1(5), ZN => n9605);
   U536 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(4), ZN => n10346);
   U537 : NAND3_X1 port map( A1 => n9531, A2 => n9605, A3 => n10346, ZN => 
                           n9395);
   U538 : AOI211_X1 port map( C1 => DATA1(3), C2 => n9868, A => n9396, B => 
                           n9395, ZN => n9401);
   U539 : NOR2_X1 port map( A1 => n10162, A2 => n9462, ZN => n9534);
   U540 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(8), ZN => n9469);
   U541 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(6), ZN => n9606);
   U542 : NAND2_X1 port map( A1 => DATA1(5), A2 => n9868, ZN => n10345);
   U543 : NAND4_X1 port map( A1 => n9397, A2 => n9469, A3 => n9606, A4 => 
                           n10345, ZN => n9398);
   U544 : NOR2_X1 port map( A1 => n9534, A2 => n9398, ZN => n9915);
   U545 : NOR2_X1 port map( A1 => n10162, A2 => n10644, ZN => n9569);
   U546 : NAND2_X1 port map( A1 => n10344, A2 => DATA1(8), ZN => n9426);
   U547 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(7), ZN => n9494);
   U548 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(5), ZN => n10107);
   U549 : NAND2_X1 port map( A1 => DATA1(4), A2 => n9853, ZN => n10804);
   U550 : NAND4_X1 port map( A1 => n9426, A2 => n9494, A3 => n10107, A4 => 
                           n10804, ZN => n9399);
   U551 : NOR2_X1 port map( A1 => n9569, A2 => n9399, ZN => n9917);
   U552 : OAI222_X1 port map( A1 => n9947, A2 => n9401, B1 => n9897, B2 => 
                           n9915, C1 => n9943, C2 => n9917, ZN => n10060);
   U553 : AOI22_X1 port map( A1 => n10355, A2 => n10059, B1 => n10056, B2 => 
                           n10060, ZN => n9414);
   U554 : OAI222_X1 port map( A1 => n9947, A2 => n9524, B1 => n9897, B2 => 
                           n9401, C1 => n9943, C2 => n9400, ZN => n10054);
   U555 : OAI222_X1 port map( A1 => n9401, A2 => n9943, B1 => n9400, B2 => 
                           n9947, C1 => n9917, C2 => n9897, ZN => n10057);
   U556 : AOI22_X1 port map( A1 => n10012, A2 => n10054, B1 => n9996, B2 => 
                           n10057, ZN => n9413);
   U557 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(8), A3 => DATA2(6), A4 
                           => DATA2(7), ZN => n9409);
   U558 : INV_X1 port map( A => DATA2(12), ZN => n10915);
   U559 : INV_X1 port map( A => DATA2(10), ZN => n10917);
   U560 : INV_X1 port map( A => DATA2(11), ZN => n10916);
   U561 : INV_X1 port map( A => DATA2(13), ZN => n10914);
   U562 : NAND4_X1 port map( A1 => n10915, A2 => n10917, A3 => n10916, A4 => 
                           n10914, ZN => n9402);
   U563 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n9837, A4 
                           => n9402, ZN => n9408);
   U564 : NOR4_X1 port map( A1 => DATA1(14), A2 => DATA1(12), A3 => n11228, A4 
                           => n9763, ZN => n9406);
   U565 : NOR4_X1 port map( A1 => DATA1(13), A2 => DATA1(9), A3 => DATA1(8), A4
                           => DATA1(7), ZN => n9405);
   U566 : NOR4_X1 port map( A1 => DATA1(15), A2 => DATA1(6), A3 => DATA1(5), A4
                           => DATA1(4), ZN => n9404);
   U567 : NOR4_X1 port map( A1 => n11227, A2 => DATA1(2), A3 => DATA1(1), A4 =>
                           DATA1(0), ZN => n9403);
   U568 : AND4_X1 port map( A1 => n9406, A2 => n9405, A3 => n9404, A4 => n9403,
                           ZN => n9407);
   U569 : AOI211_X1 port map( C1 => n9409, C2 => n9408, A => n9407, B => n553, 
                           ZN => n10214);
   U570 : CLKBUF_X1 port map( A => n10214, Z => n10583);
   U571 : INV_X1 port map( A => DATA1(9), ZN => n9532);
   U572 : NOR2_X1 port map( A1 => n9532, A2 => n10918, ZN => n9411);
   U573 : NAND3_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => n9410, ZN => 
                           n10601);
   U574 : NAND2_X1 port map( A1 => n10894, A2 => n10556, ZN => n10409);
   U575 : NAND2_X1 port map( A1 => n10601, A2 => n10409, ZN => n10578);
   U576 : AOI22_X1 port map( A1 => n10583, A2 => dataout_mul_9_port, B1 => 
                           n9411, B2 => n10578, ZN => n9412);
   U577 : OAI221_X1 port map( B1 => n10559, B2 => n9414, C1 => n10559, C2 => 
                           n9413, A => n9412, ZN => n9415);
   U578 : AOI211_X1 port map( C1 => n10556, C2 => n10618, A => n9416, B => 
                           n9415, ZN => n9420);
   U579 : AND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n9417);
   U580 : NOR2_X1 port map( A1 => n11230, A2 => n10515, ZN => n10548);
   U581 : NAND3_X1 port map( A1 => n10660, A2 => n9418, A3 => DATA2_I_8_port, 
                           ZN => n10574);
   U582 : OAI211_X1 port map( C1 => n9418, C2 => n9417, A => n10548, B => 
                           n10574, ZN => n9419);
   U583 : OAI211_X1 port map( C1 => n9421, C2 => n10591, A => n9420, B => n9419
                           , ZN => OUTALU(9));
   U584 : AOI22_X1 port map( A1 => n10569, A2 => n9548, B1 => n10365, B2 => 
                           n10567, ZN => n9450);
   U585 : NAND3_X1 port map( A1 => n10926, A2 => n9423, A3 => n9422, ZN => 
                           n10370);
   U586 : INV_X1 port map( A => n10370, ZN => n10860);
   U587 : INV_X1 port map( A => n9424, ZN => n9536);
   U588 : INV_X1 port map( A => n9475, ZN => n9425);
   U589 : AOI22_X1 port map( A1 => n9536, A2 => n10061, B1 => n9425, B2 => 
                           n9997, ZN => n9430);
   U590 : INV_X1 port map( A => n9763, ZN => n10628);
   U591 : NOR2_X1 port map( A1 => n10162, A2 => n10628, ZN => n9821);
   U592 : NAND2_X1 port map( A1 => n9715, A2 => n11228, ZN => n9759);
   U593 : OAI211_X1 port map( C1 => n10109, C2 => n10744, A => n9426, B => 
                           n9759, ZN => n9427);
   U594 : AOI211_X1 port map( C1 => DATA1(9), C2 => n10803, A => n9821, B => 
                           n9427, ZN => n9496);
   U595 : OAI222_X1 port map( A1 => n9947, A2 => n9428, B1 => n9897, B2 => 
                           n9496, C1 => n9943, C2 => n9471, ZN => n9571);
   U596 : AOI22_X1 port map( A1 => n9571, A2 => n10056, B1 => n9472, B2 => 
                           n10058, ZN => n9429);
   U597 : OAI211_X1 port map( C1 => n10352, C2 => n9431, A => n9430, B => n9429
                           , ZN => n9574);
   U598 : INV_X1 port map( A => n9574, ZN => n9500);
   U599 : OAI22_X1 port map( A1 => n9500, A2 => n10826, B1 => n9501, B2 => 
                           n10828, ZN => n9434);
   U600 : OAI22_X1 port map( A1 => n9539, A2 => n10831, B1 => n9432, B2 => 
                           n10069, ZN => n9433);
   U601 : AOI211_X1 port map( C1 => n9924, C2 => n9435, A => n9434, B => n9433,
                           ZN => n9505);
   U602 : OAI222_X1 port map( A1 => n10844, A2 => n9479, B1 => n9813, B2 => 
                           n9505, C1 => n9436, C2 => n10839, ZN => n9566);
   U603 : INV_X1 port map( A => n9566, ZN => n9506);
   U604 : CLKBUF_X1 port map( A => n10023, Z => n10448);
   U605 : OAI22_X1 port map( A1 => n9506, A2 => n10448, B1 => n9508, B2 => 
                           n10408, ZN => n9440);
   U606 : INV_X1 port map( A => n10130, ZN => n10855);
   U607 : OAI22_X1 port map( A1 => n10072, A2 => n9438, B1 => n9437, B2 => 
                           n10855, ZN => n9439);
   U608 : AOI211_X1 port map( C1 => n10527, C2 => n9543, A => n9440, B => n9439
                           , ZN => n9581);
   U609 : INV_X1 port map( A => n9581, ZN => n9441);
   U610 : AOI22_X1 port map( A1 => n10860, A2 => n10568, B1 => n10858, B2 => 
                           n9441, ZN => n9449);
   U611 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => n10660, A => n9442, ZN
                           => n9643);
   U612 : INV_X1 port map( A => n10565, ZN => n10586);
   U613 : INV_X1 port map( A => n9643, ZN => n9447);
   U614 : AOI222_X1 port map( A1 => n10057, A2 => n10056, B1 => n10054, B2 => 
                           n10061, C1 => n10059, C2 => n10012, ZN => n9445);
   U615 : CLKBUF_X1 port map( A => n10214, Z => n10602);
   U616 : INV_X1 port map( A => n10660, ZN => n10710);
   U617 : INV_X1 port map( A => DATA2(8), ZN => n10919);
   U618 : OAI22_X1 port map( A1 => n10710, A2 => DATA2(8), B1 => n10919, B2 => 
                           n10660, ZN => n10727);
   U619 : AOI22_X1 port map( A1 => dataout_mul_8_port, A2 => n10602, B1 => 
                           n10556, B2 => n10727, ZN => n9444);
   U620 : NAND3_X1 port map( A1 => DATA2(8), A2 => DATA1(8), A3 => n10578, ZN 
                           => n9443);
   U621 : OAI211_X1 port map( C1 => n9445, C2 => n10559, A => n9444, B => n9443
                           , ZN => n9446);
   U622 : AOI221_X1 port map( B1 => n10548, B2 => n9643, C1 => n10586, C2 => 
                           n9447, A => n9446, ZN => n9448);
   U623 : OAI221_X1 port map( B1 => n10591, B2 => n9450, C1 => n10591, C2 => 
                           n9449, A => n9448, ZN => OUTALU(8));
   U624 : NOR2_X1 port map( A1 => n1992, A2 => cin, ZN => n10105);
   U625 : INV_X1 port map( A => n10340, ZN => n10336);
   U626 : INV_X1 port map( A => n9451, ZN => n9452);
   U627 : AOI21_X1 port map( B1 => n10337, B2 => n10336, A => n9452, ZN => 
                           n10104);
   U628 : OAI21_X1 port map( B1 => n10104, B2 => n10151, A => n9453, ZN => 
                           n9599);
   U629 : AOI21_X1 port map( B1 => n9631, B2 => n9599, A => n9454, ZN => n9588)
                           ;
   U630 : OAI21_X1 port map( B1 => n9588, B2 => n9593, A => n9455, ZN => n9529)
                           ;
   U631 : INV_X1 port map( A => n9555, ZN => n9557);
   U632 : AOI21_X1 port map( B1 => n9529, B2 => n9557, A => n9456, ZN => n9459)
                           ;
   U633 : NAND2_X1 port map( A1 => n10895, A2 => cin, ZN => n10338);
   U634 : INV_X1 port map( A => n10338, ZN => n10599);
   U635 : NOR2_X1 port map( A1 => n9452, A2 => n10339, ZN => n10103);
   U636 : OAI21_X1 port map( B1 => n10103, B2 => n10151, A => n9453, ZN => 
                           n9598);
   U637 : AOI21_X1 port map( B1 => n9631, B2 => n9598, A => n9454, ZN => n9587)
                           ;
   U638 : OAI21_X1 port map( B1 => n9587, B2 => n9593, A => n9455, ZN => n9528)
                           ;
   U639 : AOI21_X1 port map( B1 => n9528, B2 => n9557, A => n9456, ZN => n9458)
                           ;
   U640 : AOI22_X1 port map( A1 => n10105, A2 => n9459, B1 => n10599, B2 => 
                           n9458, ZN => n9457);
   U641 : INV_X1 port map( A => n9457, ZN => n9520);
   U642 : INV_X1 port map( A => n9521, ZN => n9519);
   U643 : OAI211_X1 port map( C1 => n9520, C2 => n9519, A => n10895, B => n9460
                           , ZN => n9489);
   U644 : INV_X1 port map( A => n10105, ZN => n10596);
   U645 : OAI22_X1 port map( A1 => n9459, A2 => n10596, B1 => n9458, B2 => 
                           n10338, ZN => n9518);
   U646 : INV_X1 port map( A => n9518, ZN => n9461);
   U647 : OAI22_X1 port map( A1 => n9461, A2 => n9519, B1 => n1992, B2 => n9460
                           , ZN => n9467);
   U648 : AOI22_X1 port map( A1 => n10061, A2 => n10059, B1 => n10056, B2 => 
                           n10054, ZN => n9465);
   U649 : CLKBUF_X1 port map( A => n10556, Z => n10476);
   U650 : NOR2_X1 port map( A1 => n9462, A2 => DATA2(7), ZN => n10711);
   U651 : INV_X1 port map( A => DATA2(7), ZN => n10922);
   U652 : NOR2_X1 port map( A1 => n10922, A2 => DATA1(7), ZN => n10728);
   U653 : OR2_X1 port map( A1 => n10711, A2 => n10728, ZN => n10617);
   U654 : AOI22_X1 port map( A1 => dataout_mul_7_port, A2 => n10602, B1 => 
                           n10476, B2 => n10617, ZN => n9464);
   U655 : NAND3_X1 port map( A1 => DATA2(7), A2 => DATA1(7), A3 => n10578, ZN 
                           => n9463);
   U656 : OAI211_X1 port map( C1 => n9465, C2 => n10559, A => n9464, B => n9463
                           , ZN => n9466);
   U657 : AOI21_X1 port map( B1 => n9488, B2 => n9467, A => n9466, ZN => n9487)
                           ;
   U658 : INV_X1 port map( A => n10373, ZN => n10870);
   U659 : INV_X1 port map( A => n10569, ZN => n10304);
   U660 : NOR2_X1 port map( A1 => n10162, A2 => n9532, ZN => n9857);
   U661 : NAND2_X1 port map( A1 => n9715, A2 => n9763, ZN => n9765);
   U662 : OAI211_X1 port map( C1 => n9800, C2 => n10555, A => n9765, B => n9469
                           , ZN => n9470);
   U663 : AOI211_X1 port map( C1 => n10344, C2 => DATA1(7), A => n9857, B => 
                           n9470, ZN => n9535);
   U664 : OAI222_X1 port map( A1 => n9947, A2 => n9471, B1 => n9897, B2 => 
                           n9535, C1 => n9943, C2 => n9496, ZN => n9613);
   U665 : AOI22_X1 port map( A1 => n9996, A2 => n9571, B1 => n10056, B2 => 
                           n9613, ZN => n9474);
   U666 : AOI22_X1 port map( A1 => n10058, A2 => n9536, B1 => n9997, B2 => 
                           n9472, ZN => n9473);
   U667 : OAI211_X1 port map( C1 => n10352, C2 => n9475, A => n9474, B => n9473
                           , ZN => n9504);
   U668 : INV_X1 port map( A => n9504, ZN => n9602);
   U669 : OAI22_X1 port map( A1 => n9539, A2 => n10828, B1 => n9602, B2 => 
                           n10826, ZN => n9477);
   U670 : OAI22_X1 port map( A1 => n9501, A2 => n10069, B1 => n9500, B2 => 
                           n10831, ZN => n9476);
   U671 : AOI211_X1 port map( C1 => n9924, C2 => n9478, A => n9477, B => n9476,
                           ZN => n9542);
   U672 : OAI222_X1 port map( A1 => n10844, A2 => n9505, B1 => n9813, B2 => 
                           n9542, C1 => n9479, C2 => n10839, ZN => n9618);
   U673 : AOI22_X1 port map( A1 => n10531, A2 => n9481, B1 => n10849, B2 => 
                           n9480, ZN => n9482);
   U674 : OAI21_X1 port map( B1 => n9507, B2 => n10408, A => n9482, ZN => n9483
                           );
   U675 : AOI21_X1 port map( B1 => n10848, B2 => n9618, A => n9483, ZN => n9600
                           );
   U676 : OAI21_X1 port map( B1 => n10431, B2 => n9506, A => n9600, ZN => n9491
                           );
   U677 : AOI22_X1 port map( A1 => n10797, A2 => n10568, B1 => n10858, B2 => 
                           n9491, ZN => n9485);
   U678 : AOI22_X1 port map( A1 => n10860, A2 => n10567, B1 => n10365, B2 => 
                           n9548, ZN => n9484);
   U679 : OAI211_X1 port map( C1 => n9581, C2 => n10304, A => n9485, B => n9484
                           , ZN => n9550);
   U680 : NAND3_X1 port map( A1 => n10885, A2 => n10870, A3 => n9550, ZN => 
                           n9486);
   U681 : OAI211_X1 port map( C1 => n9489, C2 => n9488, A => n9487, B => n9486,
                           ZN => OUTALU(7));
   U682 : NOR2_X1 port map( A1 => n10925, A2 => n9490, ZN => n10866);
   U683 : INV_X1 port map( A => n10866, ZN => n10375);
   U684 : NAND2_X1 port map( A1 => n10375, A2 => n10373, ZN => n10376);
   U685 : INV_X1 port map( A => n10376, ZN => n10868);
   U686 : INV_X1 port map( A => n9491, ZN => n9582);
   U687 : OAI22_X1 port map( A1 => n9582, A2 => n10304, B1 => n9492, B2 => 
                           n10077, ZN => n9493);
   U688 : INV_X1 port map( A => n9493, ZN => n9512);
   U689 : AOI22_X1 port map( A1 => DATA1(6), A2 => n10344, B1 => DATA1(10), B2 
                           => n9853, ZN => n9495);
   U690 : NAND2_X1 port map( A1 => n10183, A2 => n10660, ZN => n9871);
   U691 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(9), ZN => n9822);
   U692 : AND4_X1 port map( A1 => n9495, A2 => n9494, A3 => n9871, A4 => n9822,
                           ZN => n9570);
   U693 : OAI222_X1 port map( A1 => n9535, A2 => n9943, B1 => n9496, B2 => 
                           n9947, C1 => n9570, C2 => n9897, ZN => n10118);
   U694 : AOI22_X1 port map( A1 => n9536, A2 => n10355, B1 => n10056, B2 => 
                           n10118, ZN => n9498);
   U695 : AOI22_X1 port map( A1 => n9571, A2 => n10058, B1 => n9613, B2 => 
                           n9996, ZN => n9497);
   U696 : OAI211_X1 port map( C1 => n10352, C2 => n9499, A => n9498, B => n9497
                           , ZN => n10123);
   U697 : INV_X1 port map( A => n10123, ZN => n9601);
   U698 : OAI22_X1 port map( A1 => n9500, A2 => n10828, B1 => n9601, B2 => 
                           n10826, ZN => n9503);
   U699 : OAI22_X1 port map( A1 => n10834, A2 => n9501, B1 => n9539, B2 => 
                           n10069, ZN => n9502);
   U700 : AOI211_X1 port map( C1 => n10554, C2 => n9504, A => n9503, B => n9502
                           , ZN => n9578);
   U701 : OAI222_X1 port map( A1 => n10842, A2 => n9578, B1 => n10844, B2 => 
                           n9542, C1 => n9505, C2 => n10839, ZN => n9619);
   U702 : INV_X1 port map( A => n9619, ZN => n10134);
   U703 : OAI22_X1 port map( A1 => n10134, A2 => n10448, B1 => n9506, B2 => 
                           n10408, ZN => n9510);
   U704 : OAI22_X1 port map( A1 => n10133, A2 => n9508, B1 => n9507, B2 => 
                           n10855, ZN => n9509);
   U705 : AOI211_X1 port map( C1 => n10852, C2 => n9618, A => n9510, B => n9509
                           , ZN => n9622);
   U706 : INV_X1 port map( A => n9622, ZN => n10139);
   U707 : AOI22_X1 port map( A1 => n10139, A2 => n10858, B1 => n9548, B2 => 
                           n10860, ZN => n9511);
   U708 : OAI211_X1 port map( C1 => n10863, C2 => n9581, A => n9512, B => n9511
                           , ZN => n9549);
   U709 : AOI22_X1 port map( A1 => n10868, A2 => n9550, B1 => n10870, B2 => 
                           n9549, ZN => n9523);
   U710 : NAND2_X1 port map( A1 => n10644, A2 => DATA2(6), ZN => n10725);
   U711 : OAI21_X1 port map( B1 => n10644, B2 => DATA2(6), A => n10725, ZN => 
                           n9513);
   U712 : INV_X1 port map( A => n9513, ZN => n10629);
   U713 : INV_X1 port map( A => n10556, ZN => n10594);
   U714 : OAI21_X1 port map( B1 => n10601, B2 => n10644, A => n10409, ZN => 
                           n9514);
   U715 : AOI22_X1 port map( A1 => DATA2(6), A2 => n9514, B1 => n10214, B2 => 
                           dataout_mul_6_port, ZN => n9516);
   U716 : NAND3_X1 port map( A1 => n10577, A2 => n10056, A3 => n10059, ZN => 
                           n9515);
   U717 : OAI211_X1 port map( C1 => n10629, C2 => n10594, A => n9516, B => 
                           n9515, ZN => n9517);
   U718 : AOI221_X1 port map( B1 => n9521, B2 => n9520, C1 => n9519, C2 => 
                           n9518, A => n9517, ZN => n9522);
   U719 : OAI21_X1 port map( B1 => n9523, B2 => n10591, A => n9522, ZN => 
                           OUTALU(6));
   U720 : OAI21_X1 port map( B1 => n10601, B2 => n9527, A => n10409, ZN => 
                           n9526);
   U721 : OAI22_X1 port map( A1 => n9524, A2 => n9897, B1 => n9561, B2 => n9943
                           , ZN => n9525);
   U722 : AOI22_X1 port map( A1 => DATA2(5), A2 => n9526, B1 => n10438, B2 => 
                           n9525, ZN => n9560);
   U723 : INV_X1 port map( A => DATA2(5), ZN => n10924);
   U724 : NAND2_X1 port map( A1 => DATA1(5), A2 => n10924, ZN => n10720);
   U725 : NAND2_X1 port map( A1 => DATA2(5), A2 => n9527, ZN => n10724);
   U726 : NAND2_X1 port map( A1 => n10720, A2 => n10724, ZN => n10613);
   U727 : AOI22_X1 port map( A1 => dataout_mul_5_port, A2 => n10602, B1 => 
                           n10476, B2 => n10613, ZN => n9559);
   U728 : OAI22_X1 port map( A1 => n10596, A2 => n9529, B1 => n10338, B2 => 
                           n9528, ZN => n9556);
   U729 : AOI22_X1 port map( A1 => n9529, A2 => n10105, B1 => n9528, B2 => 
                           n10599, ZN => n9530);
   U730 : INV_X1 port map( A => n9530, ZN => n9554);
   U731 : INV_X1 port map( A => n10118, ZN => n9610);
   U732 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(8), ZN => n9855);
   U733 : OAI211_X1 port map( C1 => n10109, C2 => n9532, A => n9855, B => n9531
                           , ZN => n9533);
   U734 : AOI211_X1 port map( C1 => n10344, C2 => DATA1(5), A => n9534, B => 
                           n9533, ZN => n9604);
   U735 : OAI222_X1 port map( A1 => n9875, A2 => n9535, B1 => n9945, B2 => 
                           n9604, C1 => n9943, C2 => n9570, ZN => n10119);
   U736 : AOI22_X1 port map( A1 => n10058, A2 => n9613, B1 => n10056, B2 => 
                           n10119, ZN => n9538);
   U737 : AOI22_X1 port map( A1 => n9997, A2 => n9571, B1 => n10825, B2 => 
                           n9536, ZN => n9537);
   U738 : OAI211_X1 port map( C1 => n9610, C2 => n10818, A => n9538, B => n9537
                           , ZN => n10122);
   U739 : INV_X1 port map( A => n10122, ZN => n10357);
   U740 : OAI22_X1 port map( A1 => n10826, A2 => n10357, B1 => n10828, B2 => 
                           n9602, ZN => n9541);
   U741 : OAI22_X1 port map( A1 => n10831, A2 => n9601, B1 => n9539, B2 => 
                           n10834, ZN => n9540);
   U742 : AOI211_X1 port map( C1 => n9574, C2 => n10838, A => n9541, B => n9540
                           , ZN => n9617);
   U743 : OAI222_X1 port map( A1 => n9542, A2 => n10839, B1 => n9578, B2 => 
                           n10844, C1 => n9617, C2 => n9813, ZN => n10361);
   U744 : AOI22_X1 port map( A1 => n10848, A2 => n10361, B1 => n10846, B2 => 
                           n9618, ZN => n9545);
   U745 : AOI22_X1 port map( A1 => n10531, A2 => n9566, B1 => n10849, B2 => 
                           n9543, ZN => n9544);
   U746 : OAI211_X1 port map( C1 => n10134, C2 => n10431, A => n9545, B => 
                           n9544, ZN => n10366);
   U747 : INV_X1 port map( A => n10366, ZN => n10135);
   U748 : CLKBUF_X1 port map( A => n10322, Z => n10284);
   U749 : OAI22_X1 port map( A1 => n10135, A2 => n10284, B1 => n9622, B2 => 
                           n10304, ZN => n9547);
   U750 : OAI22_X1 port map( A1 => n9582, A2 => n10863, B1 => n9581, B2 => 
                           n10370, ZN => n9546);
   U751 : AOI211_X1 port map( C1 => n10797, C2 => n9548, A => n9547, B => n9546
                           , ZN => n9625);
   U752 : INV_X1 port map( A => n9549, ZN => n9585);
   U753 : INV_X1 port map( A => n9550, ZN => n9551);
   U754 : OAI222_X1 port map( A1 => n9625, A2 => n10373, B1 => n9585, B2 => 
                           n10376, C1 => n9551, C2 => n10375, ZN => n10141);
   U755 : INV_X1 port map( A => n10141, ZN => n10381);
   U756 : OAI21_X1 port map( B1 => n10925, B2 => n9552, A => n10037, ZN => 
                           n10882);
   U757 : NOR3_X1 port map( A1 => n10381, A2 => n10591, A3 => n10882, ZN => 
                           n9553);
   U758 : AOI221_X1 port map( B1 => n9557, B2 => n9556, C1 => n9555, C2 => 
                           n9554, A => n9553, ZN => n9558);
   U759 : NAND3_X1 port map( A1 => n9560, A2 => n9559, A3 => n9558, ZN => 
                           OUTALU(5));
   U760 : AOI22_X1 port map( A1 => n10105, A2 => n9588, B1 => n10599, B2 => 
                           n9587, ZN => n9594);
   U761 : NOR3_X1 port map( A1 => n9561, A2 => n10559, A3 => n9897, ZN => n9565
                           );
   U762 : NAND2_X1 port map( A1 => n9562, A2 => DATA2(4), ZN => n10652);
   U763 : NAND2_X1 port map( A1 => n10925, A2 => DATA1(4), ZN => n10721);
   U764 : NAND3_X1 port map( A1 => DATA1(4), A2 => DATA2(4), A3 => n10578, ZN 
                           => n9563);
   U765 : OAI221_X1 port map( B1 => n10594, B2 => n10652, C1 => n10594, C2 => 
                           n10721, A => n9563, ZN => n9564);
   U766 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n10583, A => 
                           n9565, B => n9564, ZN => n9592);
   U767 : AOI22_X1 port map( A1 => n10130, A2 => n9618, B1 => n10849, B2 => 
                           n9566, ZN => n9580);
   U768 : INV_X1 port map( A => n10119, ZN => n10351);
   U769 : NAND2_X1 port map( A1 => n9715, A2 => DATA1(7), ZN => n9870);
   U770 : OAI211_X1 port map( C1 => n9800, C2 => n10710, A => n9567, B => n9870
                           , ZN => n9568);
   U771 : AOI211_X1 port map( C1 => n10344, C2 => DATA1(4), A => n9569, B => 
                           n9568, ZN => n9603);
   U772 : OAI222_X1 port map( A1 => n9875, A2 => n9570, B1 => n9897, B2 => 
                           n9603, C1 => n9943, C2 => n9604, ZN => n10824);
   U773 : AOI22_X1 port map( A1 => n10012, A2 => n10118, B1 => n10056, B2 => 
                           n10824, ZN => n9573);
   U774 : AOI22_X1 port map( A1 => n10355, A2 => n9613, B1 => n10825, B2 => 
                           n9571, ZN => n9572);
   U775 : OAI211_X1 port map( C1 => n10351, C2 => n10818, A => n9573, B => 
                           n9572, ZN => n10830);
   U776 : AOI22_X1 port map( A1 => n10525, A2 => n10123, B1 => n10576, B2 => 
                           n10830, ZN => n9576);
   U777 : AOI22_X1 port map( A1 => n10554, A2 => n10122, B1 => n10124, B2 => 
                           n9574, ZN => n9575);
   U778 : OAI211_X1 port map( C1 => n9602, C2 => n10069, A => n9576, B => n9575
                           , ZN => n9577);
   U779 : INV_X1 port map( A => n9577, ZN => n10129);
   U780 : OAI222_X1 port map( A1 => n9578, A2 => n10839, B1 => n9617, B2 => 
                           n10844, C1 => n10129, C2 => n10842, ZN => n10850);
   U781 : AOI22_X1 port map( A1 => n10848, A2 => n10850, B1 => n10846, B2 => 
                           n9619, ZN => n9579);
   U782 : NAND2_X1 port map( A1 => n9580, A2 => n9579, ZN => n10796);
   U783 : AOI21_X1 port map( B1 => n10527, B2 => n10361, A => n10796, ZN => 
                           n10371);
   U784 : OAI22_X1 port map( A1 => n10371, A2 => n10284, B1 => n9581, B2 => 
                           n10077, ZN => n9584);
   U785 : OAI22_X1 port map( A1 => n10135, A2 => n10304, B1 => n9582, B2 => 
                           n10370, ZN => n9583);
   U786 : AOI211_X1 port map( C1 => n10365, C2 => n10139, A => n9584, B => 
                           n9583, ZN => n10140);
   U787 : OAI222_X1 port map( A1 => n10376, A2 => n9625, B1 => n10375, B2 => 
                           n9585, C1 => n10140, C2 => n10373, ZN => n10878);
   U788 : INV_X1 port map( A => n10882, ZN => n10377);
   U789 : NAND2_X1 port map( A1 => n10037, A2 => n10882, ZN => n10043);
   U790 : INV_X1 port map( A => n10043, ZN => n10875);
   U791 : AOI22_X1 port map( A1 => n10878, A2 => n10377, B1 => n10141, B2 => 
                           n10875, ZN => n9586);
   U792 : INV_X1 port map( A => n9586, ZN => n9590);
   U793 : OAI22_X1 port map( A1 => n9588, A2 => n10596, B1 => n9587, B2 => 
                           n10338, ZN => n9589);
   U794 : AOI22_X1 port map( A1 => n10482, A2 => n9590, B1 => n9593, B2 => 
                           n9589, ZN => n9591);
   U795 : OAI211_X1 port map( C1 => n9594, C2 => n9593, A => n9592, B => n9591,
                           ZN => OUTALU(4));
   U796 : INV_X1 port map( A => DATA1(1), ZN => n10335);
   U797 : AOI22_X1 port map( A1 => n10803, A2 => DATA1(2), B1 => n9697, B2 => 
                           DATA1(0), ZN => n9596);
   U798 : NAND2_X1 port map( A1 => n10802, A2 => n11227, ZN => n9595);
   U799 : OAI211_X1 port map( C1 => n10162, C2 => n10335, A => n9596, B => 
                           n9595, ZN => n9597);
   U800 : AOI22_X1 port map( A1 => n10583, A2 => dataout_mul_3_port, B1 => 
                           n10577, B2 => n9597, ZN => n9636);
   U801 : OAI22_X1 port map( A1 => n10596, A2 => n9599, B1 => n10338, B2 => 
                           n9598, ZN => n9630);
   U802 : AOI22_X1 port map( A1 => n10105, A2 => n9599, B1 => n10599, B2 => 
                           n9598, ZN => n9628);
   U803 : OAI22_X1 port map( A1 => n10371, A2 => n10304, B1 => n9600, B2 => 
                           n10077, ZN => n9624);
   U804 : INV_X1 port map( A => n10850, ZN => n10364);
   U805 : OAI22_X1 port map( A1 => n9602, A2 => n10834, B1 => n9601, B2 => 
                           n10069, ZN => n9615);
   U806 : INV_X1 port map( A => n9603, ZN => n10113);
   U807 : INV_X1 port map( A => n9604, ZN => n9609);
   U808 : AOI22_X1 port map( A1 => DATA1(3), A2 => n10344, B1 => DATA1(7), B2 
                           => n9853, ZN => n9608);
   U809 : NAND4_X1 port map( A1 => n9608, A2 => n9607, A3 => n9606, A4 => n9605
                           , ZN => n10350);
   U810 : AOI222_X1 port map( A1 => n10113, A2 => n10812, B1 => n9609, B2 => 
                           n10810, C1 => n10350, C2 => n10349, ZN => n10821);
   U811 : OAI22_X1 port map( A1 => n10115, A2 => n10821, B1 => n9610, B2 => 
                           n10820, ZN => n9612);
   U812 : INV_X1 port map( A => n10824, ZN => n10116);
   U813 : OAI22_X1 port map( A1 => n10351, A2 => n10814, B1 => n10116, B2 => 
                           n10818, ZN => n9611);
   U814 : AOI211_X1 port map( C1 => n10825, C2 => n9613, A => n9612, B => n9611
                           , ZN => n10801);
   U815 : OAI22_X1 port map( A1 => n10357, A2 => n10828, B1 => n10801, B2 => 
                           n10826, ZN => n9614);
   U816 : NOR2_X1 port map( A1 => n9615, A2 => n9614, ZN => n10360);
   U817 : INV_X1 port map( A => n10360, ZN => n9616);
   U818 : AOI21_X1 port map( B1 => n10830, B2 => n10554, A => n9616, ZN => 
                           n10128);
   U819 : OAI222_X1 port map( A1 => n9617, A2 => n10839, B1 => n10129, B2 => 
                           n10844, C1 => n10128, C2 => n10842, ZN => n10800);
   U820 : AOI22_X1 port map( A1 => n10848, A2 => n10800, B1 => n10846, B2 => 
                           n10361, ZN => n9621);
   U821 : AOI22_X1 port map( A1 => n10531, A2 => n9619, B1 => n10849, B2 => 
                           n9618, ZN => n9620);
   U822 : OAI211_X1 port map( C1 => n10364, C2 => n10431, A => n9621, B => 
                           n9620, ZN => n10859);
   U823 : INV_X1 port map( A => n10859, ZN => n10136);
   U824 : OAI22_X1 port map( A1 => n10136, A2 => n10284, B1 => n9622, B2 => 
                           n10370, ZN => n9623);
   U825 : AOI211_X1 port map( C1 => n10365, C2 => n10366, A => n9624, B => 
                           n9623, ZN => n10374);
   U826 : OAI222_X1 port map( A1 => n10376, A2 => n10140, B1 => n10375, B2 => 
                           n9625, C1 => n10374, C2 => n10373, ZN => n10876);
   U827 : NOR2_X1 port map( A1 => n10037, A2 => n9626, ZN => n10873);
   U828 : AOI222_X1 port map( A1 => n10876, A2 => n10377, B1 => n10141, B2 => 
                           n10873, C1 => n10878, C2 => n10875, ZN => n9627);
   U829 : OAI22_X1 port map( A1 => n9631, A2 => n9628, B1 => n9627, B2 => 
                           n10591, ZN => n9629);
   U830 : AOI21_X1 port map( B1 => n9631, B2 => n9630, A => n9629, ZN => n9635)
                           ;
   U831 : NAND3_X1 port map( A1 => n11227, A2 => DATA2(3), A3 => n10578, ZN => 
                           n9634);
   U832 : NOR2_X1 port map( A1 => DATA2(3), A2 => n9632, ZN => n10716);
   U833 : NOR2_X1 port map( A1 => n11227, A2 => n10926, ZN => n10649);
   U834 : OAI21_X1 port map( B1 => n10716, B2 => n10649, A => n10556, ZN => 
                           n9633);
   U835 : NAND4_X1 port map( A1 => n9636, A2 => n9635, A3 => n9634, A4 => n9633
                           , ZN => OUTALU(3));
   U836 : INV_X1 port map( A => DATA1(31), ZN => n10180);
   U837 : NOR2_X1 port map( A1 => n9837, A2 => n10180, ZN => n9940);
   U838 : AOI22_X1 port map( A1 => n10482, A2 => n9940, B1 => n10214, B2 => 
                           dataout_mul_31_port, ZN => n10089);
   U839 : NOR2_X1 port map( A1 => n10180, A2 => DATA2(31), ZN => n10703);
   U840 : INV_X1 port map( A => n10703, ZN => n10795);
   U841 : INV_X1 port map( A => DATA2(31), ZN => n10896);
   U842 : NOR2_X1 port map( A1 => n10896, A2 => DATA1(31), ZN => n10706);
   U843 : INV_X1 port map( A => n10706, ZN => n10791);
   U844 : NAND2_X1 port map( A1 => n10795, A2 => n10791, ZN => n10605);
   U845 : AOI211_X1 port map( C1 => n10409, C2 => n10601, A => n10180, B => 
                           n10896, ZN => n9653);
   U846 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n9637);
   U847 : OAI21_X1 port map( B1 => DATA1(30), B2 => DATA2_I_30_port, A => n9637
                           , ZN => n10091);
   U848 : NAND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => 
                           n10092);
   U849 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n10170);
   U850 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n10177);
   U851 : INV_X1 port map( A => n10177, ZN => n10196);
   U852 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n9638);
   U853 : INV_X1 port map( A => n9638, ZN => n10215);
   U854 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n10246);
   U855 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => n9638
                           , ZN => n10236);
   U856 : NOR2_X1 port map( A1 => n10246, A2 => n10236, ZN => n10229);
   U857 : NOR2_X1 port map( A1 => n10215, A2 => n10229, ZN => n10219);
   U858 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n9649);
   U859 : OAI21_X1 port map( B1 => DATA1(26), B2 => DATA2_I_26_port, A => n9649
                           , ZN => n10221);
   U860 : OAI21_X1 port map( B1 => n10219, B2 => n10221, A => n9649, ZN => 
                           n10198);
   U861 : NOR2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n10195);
   U862 : OAI21_X1 port map( B1 => DATA1(28), B2 => DATA2_I_28_port, A => 
                           n10170, ZN => n10189);
   U863 : NOR2_X1 port map( A1 => n10195, A2 => n10189, ZN => n9650);
   U864 : OAI21_X1 port map( B1 => n10196, B2 => n10198, A => n9650, ZN => 
                           n10175);
   U865 : OAI21_X1 port map( B1 => DATA1(29), B2 => DATA2_I_29_port, A => 
                           n10092, ZN => n10171);
   U866 : AOI21_X1 port map( B1 => n10170, B2 => n10175, A => n10171, ZN => 
                           n10046);
   U867 : XOR2_X1 port map( A => DATA2_I_23_port, B => DATA1(23), Z => n10278);
   U868 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n10273);
   U869 : OAI21_X1 port map( B1 => DATA1(22), B2 => DATA2_I_22_port, A => 
                           n10273, ZN => n10287);
   U870 : XOR2_X1 port map( A => DATA2_I_21_port, B => DATA1(21), Z => n10317);
   U871 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n9639);
   U872 : INV_X1 port map( A => n9639, ZN => n10264);
   U873 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n10428);
   U874 : INV_X1 port map( A => n10428, ZN => n10445);
   U875 : XOR2_X1 port map( A => DATA2_I_17_port, B => DATA1(17), Z => n10443);
   U876 : AOI22_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, B1 => 
                           n10445, B2 => n10443, ZN => n10406);
   U877 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n10262);
   U878 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => 
                           n10262, ZN => n10424);
   U879 : OAI21_X1 port map( B1 => n10406, B2 => n10424, A => n10262, ZN => 
                           n10387);
   U880 : OAI22_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, B1 => 
                           n10264, B2 => n10387, ZN => n10319);
   U881 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n10265);
   U882 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n10265, ZN => n10330);
   U883 : OAI21_X1 port map( B1 => n10319, B2 => n10330, A => n10265, ZN => 
                           n10302);
   U884 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, B1 => 
                           n10317, B2 => n10302, ZN => n10276);
   U885 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n10444);
   U886 : INV_X1 port map( A => n10443, ZN => n10441);
   U887 : NOR2_X1 port map( A1 => n10444, A2 => n10441, ZN => n10260);
   U888 : INV_X1 port map( A => n10317, ZN => n10315);
   U889 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => n9639
                           , ZN => n10401);
   U890 : NOR4_X1 port map( A1 => n10424, A2 => n10330, A3 => n10315, A4 => 
                           n10401, ZN => n9646);
   U891 : NAND2_X1 port map( A1 => n11229, A2 => DATA2_I_15_port, ZN => n9644);
   U892 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => n9644
                           , ZN => n10473);
   U893 : XOR2_X1 port map( A => DATA2_I_14_port, B => DATA1(14), Z => n10499);
   U894 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n10495);
   U895 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => 
                           n10495, ZN => n10521);
   U896 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n10522);
   U897 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => 
                           n10522, ZN => n10542);
   U898 : NOR2_X1 port map( A1 => n10521, A2 => n10542, ZN => n10472);
   U899 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n10470);
   U900 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n10465
                           );
   U901 : NAND2_X1 port map( A1 => n9763, A2 => DATA2_I_10_port, ZN => n10467);
   U902 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n10467, ZN => n10466);
   U903 : AOI21_X1 port map( B1 => n10465, B2 => n10574, A => n10466, ZN => 
                           n10573);
   U904 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => n9763, A => n10573, 
                           ZN => n10552);
   U905 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n10468);
   U906 : OAI21_X1 port map( B1 => n10470, B2 => n10552, A => n10468, ZN => 
                           n10541);
   U907 : NOR2_X1 port map( A1 => n10522, A2 => n10521, ZN => n10471);
   U908 : AOI21_X1 port map( B1 => n10472, B2 => n10541, A => n10471, ZN => 
                           n10497);
   U909 : NAND2_X1 port map( A1 => n10497, A2 => n10495, ZN => n10492);
   U910 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n10499, B2 => n10492, ZN => n10464);
   U911 : INV_X1 port map( A => n10499, ZN => n9640);
   U912 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n10468, ZN => n10551);
   U913 : NOR4_X1 port map( A1 => n10466, A2 => n9641, A3 => n9640, A4 => 
                           n10551, ZN => n9642);
   U914 : NAND4_X1 port map( A1 => n10472, A2 => n9643, A3 => n9642, A4 => 
                           n10515, ZN => n9645);
   U915 : OAI221_X1 port map( B1 => n10473, B2 => n10464, C1 => n10473, C2 => 
                           n9645, A => n9644, ZN => n10268);
   U916 : NAND3_X1 port map( A1 => n10260, A2 => n9646, A3 => n10268, ZN => 
                           n9647);
   U917 : OAI221_X1 port map( B1 => n10287, B2 => n10276, C1 => n10287, C2 => 
                           n9647, A => n10273, ZN => n9648);
   U918 : AOI22_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, B1 => 
                           n10278, B2 => n9648, ZN => n9651);
   U919 : NAND2_X1 port map( A1 => n10895, A2 => n9651, ZN => n10228);
   U920 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n10253);
   U921 : NOR2_X1 port map( A1 => n10253, A2 => n10236, ZN => n10216);
   U922 : NOR2_X1 port map( A1 => n10215, A2 => n10216, ZN => n10218);
   U923 : OAI21_X1 port map( B1 => n10218, B2 => n10221, A => n9649, ZN => 
                           n10197);
   U924 : OAI21_X1 port map( B1 => n10196, B2 => n10197, A => n9650, ZN => 
                           n10174);
   U925 : AOI21_X1 port map( B1 => n10170, B2 => n10174, A => n10171, ZN => 
                           n10045);
   U926 : NOR2_X1 port map( A1 => n11230, A2 => n9651, ZN => n10252);
   U927 : INV_X1 port map( A => n10252, ZN => n10217);
   U928 : OAI22_X1 port map( A1 => n10046, A2 => n10228, B1 => n10045, B2 => 
                           n10217, ZN => n10154);
   U929 : AOI22_X1 port map( A1 => n10895, A2 => n10091, B1 => n10092, B2 => 
                           n10154, ZN => n10090);
   U930 : XOR2_X1 port map( A => n10180, B => DATA2_I_31_port, Z => n10049);
   U931 : AOI211_X1 port map( C1 => DATA1(30), C2 => DATA2_I_30_port, A => 
                           n10090, B => n10049, ZN => n9652);
   U932 : AOI211_X1 port map( C1 => n10556, C2 => n10605, A => n9653, B => 
                           n9652, ZN => n10088);
   U933 : AOI22_X1 port map( A1 => DATA1(16), A2 => n9697, B1 => n11229, B2 => 
                           n9853, ZN => n9657);
   U934 : NAND4_X1 port map( A1 => n9657, A2 => n9656, A3 => n9655, A4 => n9654
                           , ZN => n9692);
   U935 : AOI22_X1 port map( A1 => n10183, A2 => DATA1(16), B1 => n10802, B2 =>
                           DATA1(18), ZN => n9661);
   U936 : NAND2_X1 port map( A1 => n9715, A2 => n11229, ZN => n9660);
   U937 : NAND2_X1 port map( A1 => DATA1(14), A2 => n9868, ZN => n9659);
   U938 : NAND4_X1 port map( A1 => n9661, A2 => n9660, A3 => n9659, A4 => n9658
                           , ZN => n9671);
   U939 : AND3_X1 port map( A1 => n9664, A2 => n9663, A3 => n9662, ZN => n9666)
                           ;
   U940 : OAI211_X1 port map( C1 => n9800, C2 => n10675, A => n9666, B => n9665
                           , ZN => n9691);
   U941 : AOI222_X1 port map( A1 => n9692, A2 => n10812, B1 => n9671, B2 => 
                           n10810, C1 => n9691, C2 => n10349, ZN => n9778);
   U942 : OAI211_X1 port map( C1 => n10109, C2 => n10744, A => n9668, B => 
                           n9667, ZN => n9669);
   U943 : AOI211_X1 port map( C1 => DATA1(16), C2 => n10344, A => n9670, B => 
                           n9669, ZN => n9764);
   U944 : INV_X1 port map( A => n9671, ZN => n9689);
   U945 : NAND2_X1 port map( A1 => DATA1(13), A2 => n9853, ZN => n9673);
   U946 : NAND4_X1 port map( A1 => n9675, A2 => n9674, A3 => n9673, A4 => n9672
                           , ZN => n9676);
   U947 : NOR2_X1 port map( A1 => n9677, A2 => n9676, ZN => n9753);
   U948 : OAI222_X1 port map( A1 => n9947, A2 => n9764, B1 => n9945, B2 => 
                           n9689, C1 => n9943, C2 => n9753, ZN => n9826);
   U949 : AND4_X1 port map( A1 => n9681, A2 => n9680, A3 => n9679, A4 => n9678,
                           ZN => n9682);
   U950 : NAND2_X1 port map( A1 => n9683, A2 => n9682, ZN => n9719);
   U951 : NAND2_X1 port map( A1 => DATA1(17), A2 => n9853, ZN => n9687);
   U952 : AND4_X1 port map( A1 => n9687, A2 => n9686, A3 => n9685, A4 => n9684,
                           ZN => n9688);
   U953 : OAI21_X1 port map( B1 => n9837, B2 => n10309, A => n9688, ZN => n9701
                           );
   U954 : AOI222_X1 port map( A1 => n10114, A2 => n9691, B1 => n10808, B2 => 
                           n9719, C1 => n10812, C2 => n9701, ZN => n9723);
   U955 : INV_X1 port map( A => n9723, ZN => n9730);
   U956 : AOI22_X1 port map( A1 => n10825, A2 => n9826, B1 => n10056, B2 => 
                           n9730, ZN => n9694);
   U957 : INV_X1 port map( A => n9692, ZN => n9690);
   U958 : OAI222_X1 port map( A1 => n9947, A2 => n9753, B1 => n9897, B2 => 
                           n9690, C1 => n9943, C2 => n9689, ZN => n9775);
   U959 : AOI222_X1 port map( A1 => n10114, A2 => n9692, B1 => n10808, B2 => 
                           n9701, C1 => n10812, C2 => n9691, ZN => n9727);
   U960 : INV_X1 port map( A => n9727, ZN => n9754);
   U961 : AOI22_X1 port map( A1 => n9997, A2 => n9775, B1 => n10061, B2 => 
                           n9754, ZN => n9693);
   U962 : OAI211_X1 port map( C1 => n9778, C2 => n10814, A => n9694, B => n9693
                           , ZN => n9819);
   U963 : INV_X1 port map( A => DATA1(19), ZN => n10392);
   U964 : NOR2_X1 port map( A1 => n9800, A2 => n10392, ZN => n9696);
   U965 : AOI211_X1 port map( C1 => n9697, C2 => DATA1(20), A => n9696, B => 
                           n9695, ZN => n9700);
   U966 : NAND3_X1 port map( A1 => n9700, A2 => n9699, A3 => n9698, ZN => n9720
                           );
   U967 : AOI222_X1 port map( A1 => n9719, A2 => n10812, B1 => n9701, B2 => 
                           n10114, C1 => n9720, C2 => n10349, ZN => n9726);
   U968 : OAI22_X1 port map( A1 => n10115, A2 => n9726, B1 => n9727, B2 => 
                           n10814, ZN => n9703);
   U969 : INV_X1 port map( A => n9775, ZN => n9773);
   U970 : OAI22_X1 port map( A1 => n10352, A2 => n9773, B1 => n9778, B2 => 
                           n10820, ZN => n9702);
   U971 : AOI211_X1 port map( C1 => n9996, C2 => n9730, A => n9703, B => n9702,
                           ZN => n9783);
   U972 : AOI22_X1 port map( A1 => DATA1(22), A2 => n9715, B1 => DATA1(21), B2 
                           => n9853, ZN => n9707);
   U973 : NAND2_X1 port map( A1 => n9941, A2 => DATA1(24), ZN => n9705);
   U974 : NAND4_X1 port map( A1 => n9707, A2 => n9706, A3 => n9705, A4 => n9704
                           , ZN => n9733);
   U975 : AOI211_X1 port map( C1 => DATA1(20), C2 => n9868, A => n9709, B => 
                           n9708, ZN => n9712);
   U976 : NAND3_X1 port map( A1 => n9712, A2 => n9711, A3 => n9710, ZN => n9718
                           );
   U977 : INV_X1 port map( A => DATA1(24), ZN => n10694);
   U978 : NOR2_X1 port map( A1 => n10109, A2 => n10768, ZN => n9714);
   U979 : AOI211_X1 port map( C1 => n9715, C2 => DATA1(23), A => n9714, B => 
                           n9713, ZN => n9717);
   U980 : OAI211_X1 port map( C1 => n10694, C2 => n10162, A => n9717, B => 
                           n9716, ZN => n9738);
   U981 : AOI222_X1 port map( A1 => n9733, A2 => n10812, B1 => n9718, B2 => 
                           n10114, C1 => n9738, C2 => n10349, ZN => n9740);
   U982 : AOI222_X1 port map( A1 => n9718, A2 => n10812, B1 => n9720, B2 => 
                           n10114, C1 => n9733, C2 => n10349, ZN => n9806);
   U983 : OAI22_X1 port map( A1 => n10817, A2 => n9740, B1 => n9806, B2 => 
                           n10818, ZN => n9722);
   U984 : AOI222_X1 port map( A1 => n9720, A2 => n10812, B1 => n9719, B2 => 
                           n10114, C1 => n9718, C2 => n10349, ZN => n9793);
   U985 : OAI22_X1 port map( A1 => n9726, A2 => n10820, B1 => n9793, B2 => 
                           n10814, ZN => n9721);
   U986 : AOI211_X1 port map( C1 => n10825, C2 => n9730, A => n9722, B => n9721
                           , ZN => n9745);
   U987 : OAI22_X1 port map( A1 => n9783, A2 => n10069, B1 => n9745, B2 => 
                           n10826, ZN => n9732);
   U988 : INV_X1 port map( A => n9726, ZN => n9741);
   U989 : OAI22_X1 port map( A1 => n10817, A2 => n9793, B1 => n9723, B2 => 
                           n10814, ZN => n9725);
   U990 : OAI22_X1 port map( A1 => n10352, A2 => n9778, B1 => n9727, B2 => 
                           n10820, ZN => n9724);
   U991 : AOI211_X1 port map( C1 => n10061, C2 => n9741, A => n9725, B => n9724
                           , ZN => n9797);
   U992 : OAI22_X1 port map( A1 => n10817, A2 => n9806, B1 => n9726, B2 => 
                           n10814, ZN => n9729);
   U993 : OAI22_X1 port map( A1 => n10352, A2 => n9727, B1 => n9793, B2 => 
                           n10818, ZN => n9728);
   U994 : AOI211_X1 port map( C1 => n9997, C2 => n9730, A => n9729, B => n9728,
                           ZN => n9809);
   U995 : OAI22_X1 port map( A1 => n9797, A2 => n10828, B1 => n9809, B2 => 
                           n10831, ZN => n9731);
   U996 : AOI211_X1 port map( C1 => n9924, C2 => n9819, A => n9732, B => n9731,
                           ZN => n9816);
   U997 : INV_X1 port map( A => n9809, ZN => n9794);
   U998 : INV_X1 port map( A => n9797, ZN => n9744);
   U999 : INV_X1 port map( A => n9806, ZN => n9790);
   U1000 : INV_X1 port map( A => n9733, ZN => n9739);
   U1001 : OAI211_X1 port map( C1 => n9800, C2 => n10256, A => n9735, B => 
                           n9734, ZN => n9736);
   U1002 : AOI211_X1 port map( C1 => DATA1(26), C2 => n9941, A => n9737, B => 
                           n9736, ZN => n9803);
   U1003 : INV_X1 port map( A => n9738, ZN => n9789);
   U1004 : OAI222_X1 port map( A1 => n9875, A2 => n9739, B1 => n9945, B2 => 
                           n9803, C1 => n9943, C2 => n9789, ZN => n9950);
   U1005 : AOI22_X1 port map( A1 => n10058, A2 => n9790, B1 => n10056, B2 => 
                           n9950, ZN => n9743);
   U1006 : INV_X1 port map( A => n9740, ZN => n9840);
   U1007 : AOI22_X1 port map( A1 => n10061, A2 => n9840, B1 => n10825, B2 => 
                           n9741, ZN => n9742);
   U1008 : OAI211_X1 port map( C1 => n9793, C2 => n10820, A => n9743, B => 
                           n9742, ZN => n9957);
   U1009 : AOI22_X1 port map( A1 => n10838, A2 => n9744, B1 => n10576, B2 => 
                           n9957, ZN => n9747);
   U1010 : INV_X1 port map( A => n9745, ZN => n9844);
   U1011 : NAND2_X1 port map( A1 => n10554, A2 => n9844, ZN => n9746);
   U1012 : OAI211_X1 port map( C1 => n10834, C2 => n9783, A => n9747, B => 
                           n9746, ZN => n9810);
   U1013 : AOI21_X1 port map( B1 => n10525, B2 => n9794, A => n9810, ZN => 
                           n9815);
   U1014 : NAND2_X1 port map( A1 => n11228, A2 => n9868, ZN => n9748);
   U1015 : NAND4_X1 port map( A1 => n9751, A2 => n9750, A3 => n9749, A4 => 
                           n9748, ZN => n9752);
   U1016 : AOI21_X1 port map( B1 => n10344, B2 => n11229, A => n9752, ZN => 
                           n9770);
   U1017 : OAI222_X1 port map( A1 => n9947, A2 => n9770, B1 => n9897, B2 => 
                           n9753, C1 => n9943, C2 => n9764, ZN => n9859);
   U1018 : AOI22_X1 port map( A1 => n10825, A2 => n9859, B1 => n10056, B2 => 
                           n9754, ZN => n9756);
   U1019 : AOI22_X1 port map( A1 => n9997, A2 => n9826, B1 => n10012, B2 => 
                           n9775, ZN => n9755);
   U1020 : OAI211_X1 port map( C1 => n9778, C2 => n10818, A => n9756, B => 
                           n9755, ZN => n9864);
   U1021 : INV_X1 port map( A => n9819, ZN => n9781);
   U1022 : OAI22_X1 port map( A1 => n9781, A2 => n10069, B1 => n9809, B2 => 
                           n10826, ZN => n9758);
   U1023 : OAI22_X1 port map( A1 => n9797, A2 => n10831, B1 => n9783, B2 => 
                           n10828, ZN => n9757);
   U1024 : AOI211_X1 port map( C1 => n9924, C2 => n9864, A => n9758, B => n9757
                           , ZN => n9811);
   U1025 : OAI222_X1 port map( A1 => n10844, A2 => n9816, B1 => n9813, B2 => 
                           n9815, C1 => n9811, C2 => n10839, ZN => n9887);
   U1026 : OAI211_X1 port map( C1 => n10486, C2 => n9837, A => n9760, B => 
                           n9759, ZN => n9761);
   U1027 : AOI211_X1 port map( C1 => n9763, C2 => n9868, A => n9762, B => n9761
                           , ZN => n9825);
   U1028 : OAI222_X1 port map( A1 => n9947, A2 => n9825, B1 => n9945, B2 => 
                           n9764, C1 => n9943, C2 => n9770, ZN => n9860);
   U1029 : NAND3_X1 port map( A1 => n9767, A2 => n9766, A3 => n9765, ZN => 
                           n9768);
   U1030 : AOI211_X1 port map( C1 => DATA1(9), C2 => n9868, A => n9769, B => 
                           n9768, ZN => n9858);
   U1031 : OAI222_X1 port map( A1 => n9947, A2 => n9858, B1 => n9897, B2 => 
                           n9770, C1 => n9943, C2 => n9825, ZN => n9896);
   U1032 : AOI22_X1 port map( A1 => n10355, A2 => n9860, B1 => n10825, B2 => 
                           n9896, ZN => n9772);
   U1033 : AOI22_X1 port map( A1 => n10012, A2 => n9859, B1 => n9996, B2 => 
                           n9826, ZN => n9771);
   U1034 : OAI211_X1 port map( C1 => n10115, C2 => n9773, A => n9772, B => 
                           n9771, ZN => n9879);
   U1035 : INV_X1 port map( A => n9879, ZN => n9905);
   U1036 : OAI22_X1 port map( A1 => n10826, A2 => n9783, B1 => n10834, B2 => 
                           n9905, ZN => n9774);
   U1037 : INV_X1 port map( A => n9774, ZN => n9780);
   U1038 : AOI22_X1 port map( A1 => n10355, A2 => n9859, B1 => n10012, B2 => 
                           n9826, ZN => n9777);
   U1039 : AOI22_X1 port map( A1 => n9996, A2 => n9775, B1 => n10825, B2 => 
                           n9860, ZN => n9776);
   U1040 : OAI211_X1 port map( C1 => n10817, C2 => n9778, A => n9777, B => 
                           n9776, ZN => n9880);
   U1041 : AOI22_X1 port map( A1 => n10414, A2 => n9880, B1 => n10525, B2 => 
                           n9864, ZN => n9779);
   U1042 : OAI211_X1 port map( C1 => n9781, C2 => n10831, A => n9780, B => 
                           n9779, ZN => n9867);
   U1043 : AOI22_X1 port map( A1 => n10414, A2 => n9864, B1 => n10124, B2 => 
                           n9880, ZN => n9782);
   U1044 : OAI21_X1 port map( B1 => n9783, B2 => n10831, A => n9782, ZN => 
                           n9784);
   U1045 : AOI21_X1 port map( B1 => n10525, B2 => n9819, A => n9784, ZN => 
                           n9812);
   U1046 : OAI21_X1 port map( B1 => n9797, B2 => n10826, A => n9812, ZN => 
                           n9831);
   U1047 : INV_X1 port map( A => n9811, ZN => n9785);
   U1048 : AOI222_X1 port map( A1 => n9867, A2 => n10071, B1 => n9831, B2 => 
                           n10462, C1 => n9785, C2 => n10488, ZN => n9907);
   U1049 : NAND2_X1 port map( A1 => n10344, A2 => DATA1(28), ZN => n10178);
   U1050 : OAI211_X1 port map( C1 => n9800, C2 => n10694, A => n10178, B => 
                           n9786, ZN => n9787);
   U1051 : AOI211_X1 port map( C1 => DATA1(26), C2 => n10183, A => n9788, B => 
                           n9787, ZN => n9839);
   U1052 : OAI222_X1 port map( A1 => n9947, A2 => n9789, B1 => n9945, B2 => 
                           n9839, C1 => n9943, C2 => n9803, ZN => n9936);
   U1053 : AOI22_X1 port map( A1 => n10058, A2 => n9840, B1 => n10056, B2 => 
                           n9936, ZN => n9792);
   U1054 : AOI22_X1 port map( A1 => n9997, A2 => n9790, B1 => n9996, B2 => 
                           n9950, ZN => n9791);
   U1055 : OAI211_X1 port map( C1 => n10352, C2 => n9793, A => n9792, B => 
                           n9791, ZN => n9935);
   U1056 : AOI22_X1 port map( A1 => n10525, A2 => n9844, B1 => n10576, B2 => 
                           n9935, ZN => n9796);
   U1057 : AOI22_X1 port map( A1 => n10554, A2 => n9957, B1 => n10838, B2 => 
                           n9794, ZN => n9795);
   U1058 : OAI211_X1 port map( C1 => n10834, C2 => n9797, A => n9796, B => 
                           n9795, ZN => n9848);
   U1059 : OAI211_X1 port map( C1 => n9800, C2 => n10230, A => n9799, B => 
                           n9798, ZN => n9801);
   U1060 : AOI211_X1 port map( C1 => DATA1(29), C2 => n10802, A => n9802, B => 
                           n9801, ZN => n9946);
   U1061 : OAI222_X1 port map( A1 => n9947, A2 => n9803, B1 => n9945, B2 => 
                           n9946, C1 => n9943, C2 => n9839, ZN => n9949);
   U1062 : AOI22_X1 port map( A1 => n10355, A2 => n9840, B1 => n10056, B2 => 
                           n9949, ZN => n9805);
   U1063 : AOI22_X1 port map( A1 => n10058, A2 => n9950, B1 => n10061, B2 => 
                           n9936, ZN => n9804);
   U1064 : OAI211_X1 port map( C1 => n10352, C2 => n9806, A => n9805, B => 
                           n9804, ZN => n9956);
   U1065 : AOI22_X1 port map( A1 => n10065, A2 => n9957, B1 => n10576, B2 => 
                           n9956, ZN => n9808);
   U1066 : AOI22_X1 port map( A1 => n10554, A2 => n9935, B1 => n10838, B2 => 
                           n9844, ZN => n9807);
   U1067 : OAI211_X1 port map( C1 => n10834, C2 => n9809, A => n9808, B => 
                           n9807, ZN => n9964);
   U1068 : AOI222_X1 port map( A1 => n9810, A2 => n10071, B1 => n9848, B2 => 
                           n10462, C1 => n9964, C2 => n10488, ZN => n9966);
   U1069 : OAI22_X1 port map( A1 => n10133, A2 => n9907, B1 => n9966, B2 => 
                           n10023, ZN => n9818);
   U1070 : OAI222_X1 port map( A1 => n9812, A2 => n10839, B1 => n9811, B2 => 
                           n10844, C1 => n9816, C2 => n9813, ZN => n9884);
   U1071 : INV_X1 port map( A => n9884, ZN => n9889);
   U1072 : INV_X1 port map( A => n9848, ZN => n9814);
   U1073 : OAI222_X1 port map( A1 => n9816, A2 => n10839, B1 => n9815, B2 => 
                           n10844, C1 => n9814, C2 => n9813, ZN => n9850);
   U1074 : INV_X1 port map( A => n9850, ZN => n9967);
   U1075 : OAI22_X1 port map( A1 => n9889, A2 => n10855, B1 => n9967, B2 => 
                           n10431, ZN => n9817);
   U1076 : AOI211_X1 port map( C1 => n10846, C2 => n9887, A => n9818, B => 
                           n9817, ZN => n9972);
   U1077 : INV_X1 port map( A => n9907, ZN => n9892);
   U1078 : AOI22_X1 port map( A1 => n10848, A2 => n9850, B1 => n10130, B2 => 
                           n9892, ZN => n9833);
   U1079 : AOI22_X1 port map( A1 => n9819, A2 => n10576, B1 => n9864, B2 => 
                           n10554, ZN => n9830);
   U1080 : INV_X1 port map( A => n9860, ZN => n9878);
   U1081 : NOR2_X1 port map( A1 => n10109, A2 => n10710, ZN => n9820);
   U1082 : AOI211_X1 port map( C1 => DATA1(11), C2 => n10803, A => n9821, B => 
                           n9820, ZN => n9824);
   U1083 : AND3_X1 port map( A1 => n9824, A2 => n9823, A3 => n9822, ZN => n9874
                           );
   U1084 : OAI222_X1 port map( A1 => n9858, A2 => n9943, B1 => n9874, B2 => 
                           n9875, C1 => n9825, C2 => n9897, ZN => n9918);
   U1085 : AOI22_X1 port map( A1 => n10825, A2 => n9918, B1 => n10056, B2 => 
                           n9826, ZN => n9828);
   U1086 : AOI22_X1 port map( A1 => n9859, A2 => n10061, B1 => n9896, B2 => 
                           n9997, ZN => n9827);
   U1087 : OAI211_X1 port map( C1 => n10814, C2 => n9878, A => n9828, B => 
                           n9827, ZN => n9902);
   U1088 : AOI22_X1 port map( A1 => n9924, A2 => n9902, B1 => n9880, B2 => 
                           n10525, ZN => n9829);
   U1089 : OAI211_X1 port map( C1 => n10069, C2 => n9905, A => n9830, B => 
                           n9829, ZN => n9883);
   U1090 : AOI222_X1 port map( A1 => n9927, A2 => n9867, B1 => n10488, B2 => 
                           n9831, C1 => n9883, C2 => n10071, ZN => n9888);
   U1091 : INV_X1 port map( A => n9888, ZN => n9930);
   U1092 : AOI22_X1 port map( A1 => n10527, A2 => n9887, B1 => n10849, B2 => 
                           n9930, ZN => n9832);
   U1093 : OAI211_X1 port map( C1 => n9889, C2 => n10408, A => n9833, B => 
                           n9832, ZN => n9913);
   U1094 : INV_X1 port map( A => n9956, ZN => n9847);
   U1095 : INV_X1 port map( A => n9949, ZN => n9843);
   U1096 : NOR2_X1 port map( A1 => n10333, A2 => n10158, ZN => n10182);
   U1097 : AOI211_X1 port map( C1 => DATA1(26), C2 => n9868, A => n10182, B => 
                           n9834, ZN => n9836);
   U1098 : OAI211_X1 port map( C1 => n9837, C2 => n10793, A => n9836, B => 
                           n9835, ZN => n9838);
   U1099 : INV_X1 port map( A => n9838, ZN => n9942);
   U1100 : OAI222_X1 port map( A1 => n9946, A2 => n9943, B1 => n9839, B2 => 
                           n9875, C1 => n9942, C2 => n9897, ZN => n9951);
   U1101 : AOI22_X1 port map( A1 => n10056, A2 => n9951, B1 => n9936, B2 => 
                           n10012, ZN => n9842);
   U1102 : AOI22_X1 port map( A1 => n10825, A2 => n9840, B1 => n9950, B2 => 
                           n10355, ZN => n9841);
   U1103 : OAI211_X1 port map( C1 => n10818, C2 => n9843, A => n9842, B => 
                           n9841, ZN => n9958);
   U1104 : AOI22_X1 port map( A1 => n9935, A2 => n10065, B1 => n9958, B2 => 
                           n10576, ZN => n9846);
   U1105 : AOI22_X1 port map( A1 => n9924, A2 => n9844, B1 => n9957, B2 => 
                           n10838, ZN => n9845);
   U1106 : OAI211_X1 port map( C1 => n10831, C2 => n9847, A => n9846, B => 
                           n9845, ZN => n9963);
   U1107 : AOI222_X1 port map( A1 => n9927, A2 => n9964, B1 => n10488, B2 => 
                           n9963, C1 => n9848, C2 => n10071, ZN => n9849);
   U1108 : INV_X1 port map( A => n9849, ZN => n9971);
   U1109 : AOI22_X1 port map( A1 => n10848, A2 => n9971, B1 => n10846, B2 => 
                           n9850, ZN => n9852);
   U1110 : AOI22_X1 port map( A1 => n10531, A2 => n9887, B1 => n10849, B2 => 
                           n9884, ZN => n9851);
   U1111 : OAI211_X1 port map( C1 => n9966, C2 => n10431, A => n9852, B => 
                           n9851, ZN => n9978);
   U1112 : AOI22_X1 port map( A1 => n10365, A2 => n9913, B1 => n10858, B2 => 
                           n9978, ZN => n9894);
   U1113 : INV_X1 port map( A => n9918, ZN => n9863);
   U1114 : NAND2_X1 port map( A1 => DATA1(7), A2 => n9853, ZN => n9854);
   U1115 : OAI211_X1 port map( C1 => n10628, C2 => n10333, A => n9855, B => 
                           n9854, ZN => n9856);
   U1116 : AOI211_X1 port map( C1 => n11228, C2 => n10344, A => n9857, B => 
                           n9856, ZN => n9898);
   U1117 : OAI222_X1 port map( A1 => n9947, A2 => n9898, B1 => n9897, B2 => 
                           n9858, C1 => n9943, C2 => n9874, ZN => n9914);
   U1118 : AOI22_X1 port map( A1 => n10058, A2 => n9896, B1 => n10825, B2 => 
                           n9914, ZN => n9862);
   U1119 : AOI22_X1 port map( A1 => n9996, A2 => n9860, B1 => n10056, B2 => 
                           n9859, ZN => n9861);
   U1120 : OAI211_X1 port map( C1 => n9863, C2 => n10820, A => n9862, B => 
                           n9861, ZN => n9984);
   U1121 : AOI22_X1 port map( A1 => n10576, A2 => n9864, B1 => n10124, B2 => 
                           n9984, ZN => n9866);
   U1122 : AOI22_X1 port map( A1 => n10554, A2 => n9880, B1 => n10838, B2 => 
                           n9902, ZN => n9865);
   U1123 : OAI211_X1 port map( C1 => n9905, C2 => n10828, A => n9866, B => 
                           n9865, ZN => n9906);
   U1124 : AOI222_X1 port map( A1 => n9906, A2 => n10071, B1 => n9883, B2 => 
                           n10462, C1 => n9867, C2 => n10488, ZN => n9991);
   U1125 : INV_X1 port map( A => n9902, ZN => n9989);
   U1126 : NAND2_X1 port map( A1 => DATA1(6), A2 => n9868, ZN => n9869);
   U1127 : NAND4_X1 port map( A1 => n9872, A2 => n9871, A3 => n9870, A4 => 
                           n9869, ZN => n9873);
   U1128 : AOI21_X1 port map( B1 => n9941, B2 => DATA1(9), A => n9873, ZN => 
                           n9916);
   U1129 : OAI222_X1 port map( A1 => n9898, A2 => n9943, B1 => n9916, B2 => 
                           n9875, C1 => n9874, C2 => n9897, ZN => n9995);
   U1130 : AOI22_X1 port map( A1 => n10825, A2 => n9995, B1 => n9914, B2 => 
                           n9997, ZN => n9877);
   U1131 : AOI22_X1 port map( A1 => n9896, A2 => n9996, B1 => n9918, B2 => 
                           n10012, ZN => n9876);
   U1132 : OAI211_X1 port map( C1 => n10817, C2 => n9878, A => n9877, B => 
                           n9876, ZN => n10020);
   U1133 : AOI22_X1 port map( A1 => n9924, A2 => n10020, B1 => n9879, B2 => 
                           n10554, ZN => n9882);
   U1134 : AOI22_X1 port map( A1 => n9880, A2 => n10576, B1 => n9984, B2 => 
                           n10838, ZN => n9881);
   U1135 : OAI211_X1 port map( C1 => n10828, C2 => n9989, A => n9882, B => 
                           n9881, ZN => n9926);
   U1136 : AOI222_X1 port map( A1 => n9927, A2 => n9906, B1 => n10488, B2 => 
                           n9883, C1 => n9926, C2 => n10071, ZN => n10009);
   U1137 : INV_X1 port map( A => n10009, ZN => n9994);
   U1138 : AOI22_X1 port map( A1 => n10848, A2 => n9884, B1 => n10849, B2 => 
                           n9994, ZN => n9886);
   U1139 : AOI22_X1 port map( A1 => n10527, A2 => n9892, B1 => n10846, B2 => 
                           n9930, ZN => n9885);
   U1140 : OAI211_X1 port map( C1 => n9991, C2 => n10855, A => n9886, B => 
                           n9885, ZN => n9933);
   U1141 : INV_X1 port map( A => n9887, ZN => n9968);
   U1142 : OAI22_X1 port map( A1 => n10023, A2 => n9968, B1 => n10855, B2 => 
                           n9888, ZN => n9891);
   U1143 : OAI22_X1 port map( A1 => n10431, A2 => n9889, B1 => n10133, B2 => 
                           n9991, ZN => n9890);
   U1144 : AOI211_X1 port map( C1 => n9892, C2 => n10846, A => n9891, B => 
                           n9890, ZN => n9975);
   U1145 : INV_X1 port map( A => n9975, ZN => n10034);
   U1146 : AOI22_X1 port map( A1 => n10797, A2 => n9933, B1 => n10860, B2 => 
                           n10034, ZN => n9893);
   U1147 : OAI211_X1 port map( C1 => n9972, C2 => n10304, A => n9894, B => 
                           n9893, ZN => n9895);
   U1148 : INV_X1 port map( A => n9895, ZN => n9980);
   U1149 : INV_X1 port map( A => n9896, ZN => n9901);
   U1150 : OAI222_X1 port map( A1 => n9916, A2 => n9943, B1 => n9915, B2 => 
                           n9947, C1 => n9898, C2 => n9897, ZN => n10011);
   U1151 : AOI22_X1 port map( A1 => n10825, A2 => n10011, B1 => n9914, B2 => 
                           n10058, ZN => n9900);
   U1152 : AOI22_X1 port map( A1 => n9918, A2 => n10061, B1 => n9995, B2 => 
                           n10355, ZN => n9899);
   U1153 : OAI211_X1 port map( C1 => n10817, C2 => n9901, A => n9900, B => 
                           n9899, ZN => n10010);
   U1154 : AOI22_X1 port map( A1 => n9924, A2 => n10010, B1 => n9984, B2 => 
                           n10525, ZN => n9904);
   U1155 : AOI22_X1 port map( A1 => n9902, A2 => n10554, B1 => n10020, B2 => 
                           n10838, ZN => n9903);
   U1156 : OAI211_X1 port map( C1 => n10826, C2 => n9905, A => n9904, B => 
                           n9903, ZN => n9990);
   U1157 : AOI222_X1 port map( A1 => n9927, A2 => n9926, B1 => n10488, B2 => 
                           n9906, C1 => n9990, C2 => n10071, ZN => n10024);
   U1158 : OAI22_X1 port map( A1 => n10023, A2 => n9907, B1 => n10072, B2 => 
                           n10024, ZN => n9908);
   U1159 : INV_X1 port map( A => n9908, ZN => n9910);
   U1160 : AOI22_X1 port map( A1 => n10527, A2 => n9930, B1 => n10531, B2 => 
                           n9994, ZN => n9909);
   U1161 : OAI211_X1 port map( C1 => n9991, C2 => n10408, A => n9910, B => 
                           n9909, ZN => n10007);
   U1162 : INV_X1 port map( A => n10007, ZN => n10030);
   U1163 : OAI22_X1 port map( A1 => n10077, A2 => n10030, B1 => n10284, B2 => 
                           n9972, ZN => n9912);
   U1164 : INV_X1 port map( A => n9933, ZN => n10031);
   U1165 : OAI22_X1 port map( A1 => n10370, A2 => n10031, B1 => n10863, B2 => 
                           n9975, ZN => n9911);
   U1166 : AOI211_X1 port map( C1 => n9913, C2 => n10799, A => n9912, B => 
                           n9911, ZN => n10038);
   U1167 : INV_X1 port map( A => n9913, ZN => n9974);
   U1168 : OAI22_X1 port map( A1 => n10370, A2 => n10030, B1 => n10322, B2 => 
                           n9974, ZN => n9932);
   U1169 : OAI22_X1 port map( A1 => n10855, A2 => n10024, B1 => n10408, B2 => 
                           n10009, ZN => n9929);
   U1170 : INV_X1 port map( A => n9914, ZN => n9983);
   U1171 : OAI222_X1 port map( A1 => n9947, A2 => n9917, B1 => n9945, B2 => 
                           n9916, C1 => n9943, C2 => n9915, ZN => n10055);
   U1172 : AOI22_X1 port map( A1 => n10058, A2 => n9995, B1 => n10825, B2 => 
                           n10055, ZN => n9920);
   U1173 : AOI22_X1 port map( A1 => n10355, A2 => n10011, B1 => n10056, B2 => 
                           n9918, ZN => n9919);
   U1174 : OAI211_X1 port map( C1 => n9983, C2 => n10818, A => n9920, B => 
                           n9919, ZN => n10066);
   U1175 : INV_X1 port map( A => n10020, ZN => n9922);
   U1176 : AOI22_X1 port map( A1 => n10554, A2 => n9984, B1 => n10838, B2 => 
                           n10010, ZN => n9921);
   U1177 : OAI21_X1 port map( B1 => n9922, B2 => n10828, A => n9921, ZN => 
                           n9923);
   U1178 : AOI21_X1 port map( B1 => n9924, B2 => n10066, A => n9923, ZN => 
                           n9988);
   U1179 : INV_X1 port map( A => n9988, ZN => n9925);
   U1180 : AOI222_X1 port map( A1 => n9927, A2 => n9990, B1 => n10488, B2 => 
                           n9926, C1 => n9925, C2 => n10071, ZN => n10073);
   U1181 : OAI22_X1 port map( A1 => n10431, A2 => n9991, B1 => n10072, B2 => 
                           n10073, ZN => n9928);
   U1182 : AOI211_X1 port map( C1 => n9930, C2 => n10848, A => n9929, B => 
                           n9928, ZN => n10078);
   U1183 : OAI22_X1 port map( A1 => n10304, A2 => n9975, B1 => n10077, B2 => 
                           n10078, ZN => n9931);
   U1184 : AOI211_X1 port map( C1 => n9933, C2 => n10365, A => n9932, B => 
                           n9931, ZN => n10040);
   U1185 : OAI222_X1 port map( A1 => n9980, A2 => n10373, B1 => n10038, B2 => 
                           n10376, C1 => n10040, C2 => n10375, ZN => n9934);
   U1186 : INV_X1 port map( A => n9934, ZN => n10085);
   U1187 : INV_X1 port map( A => n9935, ZN => n9961);
   U1188 : INV_X1 port map( A => n9936, ZN => n9954);
   U1189 : OAI211_X1 port map( C1 => n10109, C2 => n10193, A => n9938, B => 
                           n9937, ZN => n9939);
   U1190 : AOI211_X1 port map( C1 => DATA1(30), C2 => n9941, A => n9940, B => 
                           n9939, ZN => n9944);
   U1191 : OAI222_X1 port map( A1 => n9947, A2 => n9946, B1 => n9945, B2 => 
                           n9944, C1 => n9943, C2 => n9942, ZN => n9948);
   U1192 : AOI22_X1 port map( A1 => n10058, A2 => n9949, B1 => n10056, B2 => 
                           n9948, ZN => n9953);
   U1193 : AOI22_X1 port map( A1 => n9996, A2 => n9951, B1 => n10825, B2 => 
                           n9950, ZN => n9952);
   U1194 : OAI211_X1 port map( C1 => n9954, C2 => n10820, A => n9953, B => 
                           n9952, ZN => n9955);
   U1195 : AOI22_X1 port map( A1 => n10065, A2 => n9956, B1 => n10576, B2 => 
                           n9955, ZN => n9960);
   U1196 : AOI22_X1 port map( A1 => n10554, A2 => n9958, B1 => n10124, B2 => 
                           n9957, ZN => n9959);
   U1197 : OAI211_X1 port map( C1 => n9961, C2 => n10069, A => n9960, B => 
                           n9959, ZN => n9962);
   U1198 : AOI222_X1 port map( A1 => n9964, A2 => n10071, B1 => n9963, B2 => 
                           n10462, C1 => n9962, C2 => n10488, ZN => n9965);
   U1199 : OAI22_X1 port map( A1 => n9966, A2 => n10408, B1 => n9965, B2 => 
                           n10448, ZN => n9970);
   U1200 : OAI22_X1 port map( A1 => n10133, A2 => n9968, B1 => n9967, B2 => 
                           n10855, ZN => n9969);
   U1201 : AOI211_X1 port map( C1 => n10527, C2 => n9971, A => n9970, B => 
                           n9969, ZN => n9973);
   U1202 : OAI22_X1 port map( A1 => n10284, A2 => n9973, B1 => n9972, B2 => 
                           n10863, ZN => n9977);
   U1203 : OAI22_X1 port map( A1 => n9975, A2 => n10077, B1 => n9974, B2 => 
                           n10370, ZN => n9976);
   U1204 : AOI211_X1 port map( C1 => n10799, C2 => n9978, A => n9977, B => 
                           n9976, ZN => n9979);
   U1205 : OAI222_X1 port map( A1 => n10376, A2 => n9980, B1 => n10375, B2 => 
                           n10038, C1 => n9979, C2 => n10373, ZN => n10035);
   U1206 : INV_X1 port map( A => n10066, ZN => n9987);
   U1207 : AOI22_X1 port map( A1 => n9997, A2 => n10055, B1 => n10012, B2 => 
                           n10011, ZN => n9982);
   U1208 : AOI22_X1 port map( A1 => n10061, A2 => n9995, B1 => n10825, B2 => 
                           n10060, ZN => n9981);
   U1209 : OAI211_X1 port map( C1 => n10115, C2 => n9983, A => n9982, B => 
                           n9981, ZN => n10507);
   U1210 : AOI22_X1 port map( A1 => n10065, A2 => n10010, B1 => n10124, B2 => 
                           n10507, ZN => n9986);
   U1211 : AOI22_X1 port map( A1 => n10554, A2 => n10020, B1 => n10576, B2 => 
                           n9984, ZN => n9985);
   U1212 : OAI211_X1 port map( C1 => n9987, C2 => n10069, A => n9986, B => 
                           n9985, ZN => n10022);
   U1213 : OAI21_X1 port map( B1 => n9989, B2 => n10826, A => n9988, ZN => 
                           n10002);
   U1214 : AOI222_X1 port map( A1 => n10022, A2 => n10071, B1 => n10002, B2 => 
                           n10462, C1 => n9990, C2 => n10488, ZN => n10389);
   U1215 : OAI22_X1 port map( A1 => n10133, A2 => n10389, B1 => n10073, B2 => 
                           n10855, ZN => n9993);
   U1216 : OAI22_X1 port map( A1 => n9991, A2 => n10023, B1 => n10024, B2 => 
                           n10408, ZN => n9992);
   U1217 : AOI211_X1 port map( C1 => n10852, C2 => n9994, A => n9993, B => 
                           n9992, ZN => n10259);
   U1218 : OAI22_X1 port map( A1 => n10073, A2 => n10408, B1 => n10024, B2 => 
                           n10431, ZN => n10004);
   U1219 : INV_X1 port map( A => n10057, ZN => n10015);
   U1220 : AOI22_X1 port map( A1 => n10012, A2 => n10055, B1 => n10056, B2 => 
                           n9995, ZN => n9999);
   U1221 : AOI22_X1 port map( A1 => n9997, A2 => n10060, B1 => n9996, B2 => 
                           n10011, ZN => n9998);
   U1222 : OAI211_X1 port map( C1 => n10352, C2 => n10015, A => n9999, B => 
                           n9998, ZN => n10524);
   U1223 : AOI22_X1 port map( A1 => n10554, A2 => n10010, B1 => n10124, B2 => 
                           n10524, ZN => n10001);
   U1224 : AOI22_X1 port map( A1 => n10414, A2 => n10507, B1 => n10525, B2 => 
                           n10066, ZN => n10000);
   U1225 : NAND2_X1 port map( A1 => n10001, A2 => n10000, ZN => n10019);
   U1226 : AOI222_X1 port map( A1 => n10019, A2 => n10071, B1 => n10022, B2 => 
                           n10462, C1 => n10002, C2 => n10488, ZN => n10407);
   U1227 : OAI22_X1 port map( A1 => n10072, A2 => n10407, B1 => n10389, B2 => 
                           n10855, ZN => n10003);
   U1228 : NOR2_X1 port map( A1 => n10004, A2 => n10003, ZN => n10008);
   U1229 : OAI22_X1 port map( A1 => n10259, A2 => n10370, B1 => n10008, B2 => 
                           n10077, ZN => n10006);
   U1230 : OAI22_X1 port map( A1 => n10322, A2 => n10031, B1 => n10078, B2 => 
                           n10863, ZN => n10005);
   U1231 : AOI211_X1 port map( C1 => n10799, C2 => n10007, A => n10006, B => 
                           n10005, ZN => n10082);
   U1232 : INV_X1 port map( A => n10259, ZN => n10029);
   U1233 : OAI21_X1 port map( B1 => n10023, B2 => n10009, A => n10008, ZN => 
                           n10081);
   U1234 : INV_X1 port map( A => n10081, ZN => n10285);
   U1235 : INV_X1 port map( A => n10407, ZN => n10076);
   U1236 : INV_X1 port map( A => n10010, ZN => n10018);
   U1237 : AOI22_X1 port map( A1 => n10012, A2 => n10060, B1 => n10056, B2 => 
                           n10011, ZN => n10014);
   U1238 : AOI22_X1 port map( A1 => n10061, A2 => n10055, B1 => n10825, B2 => 
                           n10054, ZN => n10013);
   U1239 : OAI211_X1 port map( C1 => n10015, C2 => n10820, A => n10014, B => 
                           n10013, ZN => n10553);
   U1240 : AOI22_X1 port map( A1 => n10065, A2 => n10507, B1 => n10124, B2 => 
                           n10553, ZN => n10017);
   U1241 : AOI22_X1 port map( A1 => n10554, A2 => n10066, B1 => n10838, B2 => 
                           n10524, ZN => n10016);
   U1242 : OAI211_X1 port map( C1 => n10018, C2 => n10826, A => n10017, B => 
                           n10016, ZN => n10463);
   U1243 : AOI21_X1 port map( B1 => n10020, B2 => n10576, A => n10019, ZN => 
                           n10021);
   U1244 : INV_X1 port map( A => n10021, ZN => n10070);
   U1245 : AOI222_X1 port map( A1 => n10463, A2 => n10071, B1 => n10070, B2 => 
                           n10462, C1 => n10022, C2 => n10488, ZN => n10432);
   U1246 : OAI22_X1 port map( A1 => n10133, A2 => n10432, B1 => n10389, B2 => 
                           n10408, ZN => n10026);
   U1247 : OAI22_X1 port map( A1 => n10073, A2 => n10431, B1 => n10024, B2 => 
                           n10023, ZN => n10025);
   U1248 : AOI211_X1 port map( C1 => n10130, C2 => n10076, A => n10026, B => 
                           n10025, ZN => n10305);
   U1249 : OAI22_X1 port map( A1 => n10285, A2 => n10370, B1 => n10305, B2 => 
                           n10077, ZN => n10028);
   U1250 : OAI22_X1 port map( A1 => n10284, A2 => n10030, B1 => n10078, B2 => 
                           n10304, ZN => n10027);
   U1251 : AOI211_X1 port map( C1 => n10365, C2 => n10029, A => n10028, B => 
                           n10027, ZN => n10235);
   U1252 : OAI22_X1 port map( A1 => n10078, A2 => n10370, B1 => n10259, B2 => 
                           n10077, ZN => n10033);
   U1253 : OAI22_X1 port map( A1 => n10031, A2 => n10304, B1 => n10030, B2 => 
                           n10863, ZN => n10032);
   U1254 : AOI211_X1 port map( C1 => n10858, C2 => n10034, A => n10033, B => 
                           n10032, ZN => n10039);
   U1255 : OAI222_X1 port map( A1 => n10376, A2 => n10082, B1 => n10375, B2 => 
                           n10235, C1 => n10039, C2 => n10373, ZN => n10199);
   U1256 : AOI22_X1 port map( A1 => n10377, A2 => n10035, B1 => n10879, B2 => 
                           n10199, ZN => n10042);
   U1257 : NOR2_X1 port map( A1 => n10037, A2 => n10036, ZN => n10877);
   U1258 : OAI222_X1 port map( A1 => n10376, A2 => n10039, B1 => n10375, B2 => 
                           n10082, C1 => n10040, C2 => n10373, ZN => n10173);
   U1259 : OAI222_X1 port map( A1 => n10376, A2 => n10040, B1 => n10375, B2 => 
                           n10039, C1 => n10038, C2 => n10373, ZN => n10155);
   U1260 : AOI22_X1 port map( A1 => n10877, A2 => n10173, B1 => n10873, B2 => 
                           n10155, ZN => n10041);
   U1261 : OAI211_X1 port map( C1 => n10085, C2 => n10043, A => n10042, B => 
                           n10041, ZN => n10050);
   U1262 : INV_X1 port map( A => n10092, ZN => n10044);
   U1263 : INV_X1 port map( A => n10091, ZN => n10101);
   U1264 : AOI22_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, B1 => 
                           n10044, B2 => n10101, ZN => n10047);
   U1265 : INV_X1 port map( A => n10228, ZN => n10247);
   U1266 : AOI22_X1 port map( A1 => n10247, A2 => n10046, B1 => n10252, B2 => 
                           n10045, ZN => n10100);
   U1267 : OAI22_X1 port map( A1 => n10047, A2 => n11230, B1 => n10100, B2 => 
                           n10091, ZN => n10048);
   U1268 : AOI22_X1 port map( A1 => n10438, A2 => n10050, B1 => n10049, B2 => 
                           n10048, ZN => n10087);
   U1269 : INV_X1 port map( A => n10051, ZN => n10052);
   U1270 : NOR2_X1 port map( A1 => n10053, A2 => n10052, ZN => n10889);
   U1271 : AOI22_X1 port map( A1 => n10873, A2 => n10173, B1 => n10875, B2 => 
                           n10155, ZN => n10084);
   U1272 : INV_X1 port map( A => n10553, ZN => n10509);
   U1273 : INV_X1 port map( A => n10054, ZN => n10064);
   U1274 : AOI22_X1 port map( A1 => n10058, A2 => n10057, B1 => n10056, B2 => 
                           n10055, ZN => n10063);
   U1275 : AOI22_X1 port map( A1 => n10061, A2 => n10060, B1 => n10825, B2 => 
                           n10059, ZN => n10062);
   U1276 : OAI211_X1 port map( C1 => n10064, C2 => n10820, A => n10063, B => 
                           n10062, ZN => n10575);
   U1277 : AOI22_X1 port map( A1 => n10065, A2 => n10524, B1 => n10124, B2 => 
                           n10575, ZN => n10068);
   U1278 : AOI22_X1 port map( A1 => n10554, A2 => n10507, B1 => n10576, B2 => 
                           n10066, ZN => n10067);
   U1279 : OAI211_X1 port map( C1 => n10509, C2 => n10069, A => n10068, B => 
                           n10067, ZN => n10487);
   U1280 : AOI222_X1 port map( A1 => n10487, A2 => n10071, B1 => n10463, B2 => 
                           n10462, C1 => n10070, C2 => n10488, ZN => n10449);
   U1281 : OAI22_X1 port map( A1 => n10072, A2 => n10449, B1 => n10432, B2 => 
                           n10855, ZN => n10075);
   U1282 : OAI22_X1 port map( A1 => n10073, A2 => n10448, B1 => n10389, B2 => 
                           n10431, ZN => n10074);
   U1283 : AOI211_X1 port map( C1 => n10846, C2 => n10076, A => n10075, B => 
                           n10074, ZN => n10321);
   U1284 : OAI22_X1 port map( A1 => n10305, A2 => n10370, B1 => n10321, B2 => 
                           n10077, ZN => n10080);
   U1285 : OAI22_X1 port map( A1 => n10284, A2 => n10078, B1 => n10259, B2 => 
                           n10304, ZN => n10079);
   U1286 : AOI211_X1 port map( C1 => n10365, C2 => n10081, A => n10080, B => 
                           n10079, ZN => n10243);
   U1287 : OAI222_X1 port map( A1 => n10376, A2 => n10235, B1 => n10375, B2 => 
                           n10243, C1 => n10082, C2 => n10373, ZN => n10223);
   U1288 : AOI22_X1 port map( A1 => n10877, A2 => n10199, B1 => n10879, B2 => 
                           n10223, ZN => n10083);
   U1289 : OAI211_X1 port map( C1 => n10085, C2 => n10882, A => n10084, B => 
                           n10083, ZN => n10098);
   U1290 : NAND4_X1 port map( A1 => FUNC(2), A2 => n10889, A3 => n10894, A4 => 
                           n10098, ZN => n10086);
   U1291 : NAND4_X1 port map( A1 => n10089, A2 => n10088, A3 => n10087, A4 => 
                           n10086, ZN => OUTALU(31));
   U1292 : AOI21_X1 port map( B1 => n10092, B2 => n10091, A => n10090, ZN => 
                           n10097);
   U1293 : AOI22_X1 port map( A1 => n10802, A2 => n10482, B1 => DATA2(30), B2 
                           => n10578, ZN => n10095);
   U1294 : INV_X1 port map( A => DATA2(30), ZN => n10897);
   U1295 : OAI22_X1 port map( A1 => n10793, A2 => DATA2(30), B1 => n10897, B2 
                           => DATA1(30), ZN => n10701);
   U1296 : AOI22_X1 port map( A1 => dataout_mul_30_port, A2 => n10602, B1 => 
                           n10476, B2 => n10701, ZN => n10094);
   U1297 : NAND3_X1 port map( A1 => n10803, A2 => n10885, A3 => DATA1(31), ZN 
                           => n10093);
   U1298 : OAI211_X1 port map( C1 => n10095, C2 => n10793, A => n10094, B => 
                           n10093, ZN => n10096);
   U1299 : AOI211_X1 port map( C1 => n10438, C2 => n10098, A => n10097, B => 
                           n10096, ZN => n10099);
   U1300 : OAI21_X1 port map( B1 => n10101, B2 => n10100, A => n10099, ZN => 
                           OUTALU(30));
   U1301 : INV_X1 port map( A => n10151, ZN => n10153);
   U1302 : OAI22_X1 port map( A1 => n10596, A2 => n10104, B1 => n10338, B2 => 
                           n10103, ZN => n10102);
   U1303 : INV_X1 port map( A => n10102, ZN => n10152);
   U1304 : AOI22_X1 port map( A1 => n10105, A2 => n10104, B1 => n10599, B2 => 
                           n10103, ZN => n10150);
   U1305 : NAND2_X1 port map( A1 => n10344, A2 => DATA1(2), ZN => n10108);
   U1306 : NAND2_X1 port map( A1 => n10803, A2 => DATA1(1), ZN => n10106);
   U1307 : OAI211_X1 port map( C1 => n10162, C2 => n10645, A => n10108, B => 
                           n10106, ZN => n10148);
   U1308 : AOI22_X1 port map( A1 => n10873, A2 => n10878, B1 => n10875, B2 => 
                           n10876, ZN => n10143);
   U1309 : OAI211_X1 port map( C1 => n10109, C2 => n10644, A => n10108, B => 
                           n10107, ZN => n10110);
   U1310 : AOI211_X1 port map( C1 => DATA1(3), C2 => n10803, A => n10111, B => 
                           n10110, ZN => n10112);
   U1311 : INV_X1 port map( A => n10112, ZN => n10811);
   U1312 : AOI222_X1 port map( A1 => n10114, A2 => n10113, B1 => n10808, B2 => 
                           n10811, C1 => n10812, C2 => n10350, ZN => n10815);
   U1313 : OAI22_X1 port map( A1 => n10814, A2 => n10116, B1 => n10115, B2 => 
                           n10815, ZN => n10117);
   U1314 : INV_X1 port map( A => n10117, ZN => n10121);
   U1315 : AOI22_X1 port map( A1 => n10355, A2 => n10119, B1 => n10825, B2 => 
                           n10118, ZN => n10120);
   U1316 : OAI211_X1 port map( C1 => n10821, C2 => n10818, A => n10121, B => 
                           n10120, ZN => n10356);
   U1317 : AOI22_X1 port map( A1 => n10414, A2 => n10122, B1 => n10576, B2 => 
                           n10356, ZN => n10126);
   U1318 : AOI22_X1 port map( A1 => n10525, A2 => n10830, B1 => n10124, B2 => 
                           n10123, ZN => n10125);
   U1319 : OAI211_X1 port map( C1 => n10801, C2 => n10831, A => n10126, B => 
                           n10125, ZN => n10127);
   U1320 : INV_X1 port map( A => n10127, ZN => n10840);
   U1321 : OAI222_X1 port map( A1 => n10129, A2 => n10839, B1 => n10128, B2 => 
                           n10844, C1 => n10840, C2 => n10842, ZN => n10845);
   U1322 : AOI22_X1 port map( A1 => n10850, A2 => n10846, B1 => n10845, B2 => 
                           n10848, ZN => n10132);
   U1323 : AOI22_X1 port map( A1 => n10361, A2 => n10130, B1 => n10800, B2 => 
                           n10527, ZN => n10131);
   U1324 : OAI211_X1 port map( C1 => n10134, C2 => n10133, A => n10132, B => 
                           n10131, ZN => n10367);
   U1325 : INV_X1 port map( A => n10367, ZN => n10864);
   U1326 : OAI22_X1 port map( A1 => n10863, A2 => n10371, B1 => n10322, B2 => 
                           n10864, ZN => n10138);
   U1327 : OAI22_X1 port map( A1 => n10304, A2 => n10136, B1 => n10370, B2 => 
                           n10135, ZN => n10137);
   U1328 : AOI211_X1 port map( C1 => n10139, C2 => n10797, A => n10138, B => 
                           n10137, ZN => n10865);
   U1329 : OAI222_X1 port map( A1 => n10376, A2 => n10374, B1 => n10375, B2 => 
                           n10140, C1 => n10373, C2 => n10865, ZN => n10872);
   U1330 : AOI22_X1 port map( A1 => n10377, A2 => n10872, B1 => n10877, B2 => 
                           n10141, ZN => n10142);
   U1331 : AOI21_X1 port map( B1 => n10143, B2 => n10142, A => n10591, ZN => 
                           n10147);
   U1332 : AOI22_X1 port map( A1 => DATA2(2), A2 => n10715, B1 => DATA1(2), B2 
                           => n10927, ZN => n10719);
   U1333 : NOR2_X1 port map( A1 => n10927, A2 => n10715, ZN => n10144);
   U1334 : AOI22_X1 port map( A1 => n10583, A2 => dataout_mul_2_port, B1 => 
                           n10144, B2 => n10578, ZN => n10145);
   U1335 : OAI21_X1 port map( B1 => n10719, B2 => n10594, A => n10145, ZN => 
                           n10146);
   U1336 : AOI211_X1 port map( C1 => n10438, C2 => n10148, A => n10147, B => 
                           n10146, ZN => n10149);
   U1337 : OAI221_X1 port map( B1 => n10153, B2 => n10152, C1 => n10151, C2 => 
                           n10150, A => n10149, ZN => OUTALU(2));
   U1338 : INV_X1 port map( A => n10154, ZN => n10172);
   U1339 : OAI22_X1 port map( A1 => n10228, A2 => n10175, B1 => n10217, B2 => 
                           n10174, ZN => n10168);
   U1340 : AOI22_X1 port map( A1 => n10377, A2 => n10155, B1 => n10875, B2 => 
                           n10173, ZN => n10157);
   U1341 : AOI22_X1 port map( A1 => n10877, A2 => n10223, B1 => n10873, B2 => 
                           n10199, ZN => n10156);
   U1342 : AOI21_X1 port map( B1 => n10157, B2 => n10156, A => n10559, ZN => 
                           n10167);
   U1343 : NOR2_X1 port map( A1 => DATA2(29), A2 => n10158, ZN => n10790);
   U1344 : NAND2_X1 port map( A1 => n10158, A2 => DATA2(29), ZN => n10787);
   U1345 : INV_X1 port map( A => n10787, ZN => n10159);
   U1346 : NOR2_X1 port map( A1 => n10790, A2 => n10159, ZN => n10609);
   U1347 : NAND2_X1 port map( A1 => n10344, A2 => DATA1(29), ZN => n10161);
   U1348 : NAND2_X1 port map( A1 => n10803, A2 => DATA1(30), ZN => n10160);
   U1349 : OAI211_X1 port map( C1 => n10180, C2 => n10162, A => n10161, B => 
                           n10160, ZN => n10163);
   U1350 : AOI22_X1 port map( A1 => n10482, A2 => n10163, B1 => n10214, B2 => 
                           dataout_mul_29_port, ZN => n10165);
   U1351 : NAND3_X1 port map( A1 => DATA2(29), A2 => DATA1(29), A3 => n10578, 
                           ZN => n10164);
   U1352 : OAI211_X1 port map( C1 => n10609, C2 => n10594, A => n10165, B => 
                           n10164, ZN => n10166);
   U1353 : AOI211_X1 port map( C1 => n10171, C2 => n10168, A => n10167, B => 
                           n10166, ZN => n10169);
   U1354 : OAI221_X1 port map( B1 => n10172, B2 => n10171, C1 => n10172, C2 => 
                           n10170, A => n10169, ZN => OUTALU(29));
   U1355 : AOI222_X1 port map( A1 => n10173, A2 => n10377, B1 => n10223, B2 => 
                           n10873, C1 => n10199, C2 => n10875, ZN => n10192);
   U1356 : AOI22_X1 port map( A1 => n10247, A2 => n10198, B1 => n10252, B2 => 
                           n10197, ZN => n10201);
   U1357 : NOR2_X1 port map( A1 => n10195, A2 => n10201, ZN => n10190);
   U1358 : AOI22_X1 port map( A1 => n10247, A2 => n10175, B1 => n10252, B2 => 
                           n10174, ZN => n10176);
   U1359 : AOI21_X1 port map( B1 => n10177, B2 => n10189, A => n10176, ZN => 
                           n10188);
   U1360 : OAI21_X1 port map( B1 => n10180, B2 => n10179, A => n10178, ZN => 
                           n10181);
   U1361 : AOI211_X1 port map( C1 => DATA1(30), C2 => n10183, A => n10182, B =>
                           n10181, ZN => n10186);
   U1362 : INV_X1 port map( A => DATA2(28), ZN => n10899);
   U1363 : OAI22_X1 port map( A1 => n10784, A2 => DATA2(28), B1 => n10899, B2 
                           => DATA1(28), ZN => n10698);
   U1364 : AOI22_X1 port map( A1 => dataout_mul_28_port, A2 => n10602, B1 => 
                           n10476, B2 => n10698, ZN => n10185);
   U1365 : NAND3_X1 port map( A1 => DATA2(28), A2 => DATA1(28), A3 => n10578, 
                           ZN => n10184);
   U1366 : OAI211_X1 port map( C1 => n10186, C2 => n10591, A => n10185, B => 
                           n10184, ZN => n10187);
   U1367 : AOI211_X1 port map( C1 => n10190, C2 => n10189, A => n10188, B => 
                           n10187, ZN => n10191);
   U1368 : OAI21_X1 port map( B1 => n10192, B2 => n10559, A => n10191, ZN => 
                           OUTALU(28));
   U1369 : NOR2_X1 port map( A1 => n10193, A2 => DATA2(27), ZN => n10779);
   U1370 : INV_X1 port map( A => n10779, ZN => n10194);
   U1371 : NAND2_X1 port map( A1 => DATA2(27), A2 => n10193, ZN => n10783);
   U1372 : NAND2_X1 port map( A1 => n10194, A2 => n10783, ZN => n10612);
   U1373 : AOI22_X1 port map( A1 => dataout_mul_27_port, A2 => n10602, B1 => 
                           n10476, B2 => n10612, ZN => n10208);
   U1374 : NOR2_X1 port map( A1 => n10196, A2 => n10195, ZN => n10204);
   U1375 : OAI22_X1 port map( A1 => n10228, A2 => n10198, B1 => n10217, B2 => 
                           n10197, ZN => n10203);
   U1376 : AOI22_X1 port map( A1 => n10377, A2 => n10199, B1 => n10875, B2 => 
                           n10223, ZN => n10200);
   U1377 : OAI22_X1 port map( A1 => n10201, A2 => n10204, B1 => n10200, B2 => 
                           n10559, ZN => n10202);
   U1378 : AOI21_X1 port map( B1 => n10204, B2 => n10203, A => n10202, ZN => 
                           n10207);
   U1379 : NAND3_X1 port map( A1 => DATA2(27), A2 => DATA1(27), A3 => n10578, 
                           ZN => n10206);
   U1380 : NAND3_X1 port map( A1 => n10482, A2 => n10349, A3 => n10210, ZN => 
                           n10205);
   U1381 : NAND4_X1 port map( A1 => n10208, A2 => n10207, A3 => n10206, A4 => 
                           n10205, ZN => OUTALU(27));
   U1382 : NOR2_X1 port map( A1 => DATA2(26), A2 => n10778, ZN => n10780);
   U1383 : AOI21_X1 port map( B1 => DATA2(26), B2 => n10778, A => n10780, ZN =>
                           n10631);
   U1384 : AOI22_X1 port map( A1 => n10211, A2 => n10210, B1 => n10808, B2 => 
                           n10209, ZN => n10212);
   U1385 : OAI22_X1 port map( A1 => n10631, A2 => n10594, B1 => n10212, B2 => 
                           n10591, ZN => n10213);
   U1386 : AOI21_X1 port map( B1 => n10214, B2 => dataout_mul_26_port, A => 
                           n10213, ZN => n10227);
   U1387 : NOR2_X1 port map( A1 => n10215, A2 => n10221, ZN => n10222);
   U1388 : OAI22_X1 port map( A1 => n10229, A2 => n10228, B1 => n10216, B2 => 
                           n10217, ZN => n10237);
   U1389 : OAI22_X1 port map( A1 => n10219, A2 => n10228, B1 => n10218, B2 => 
                           n10217, ZN => n10220);
   U1390 : AOI22_X1 port map( A1 => n10222, A2 => n10237, B1 => n10221, B2 => 
                           n10220, ZN => n10226);
   U1391 : NAND3_X1 port map( A1 => n10577, A2 => n10377, A3 => n10223, ZN => 
                           n10225);
   U1392 : NAND3_X1 port map( A1 => DATA2(26), A2 => DATA1(26), A3 => n10578, 
                           ZN => n10224);
   U1393 : NAND4_X1 port map( A1 => n10227, A2 => n10226, A3 => n10225, A4 => 
                           n10224, ZN => OUTALU(26));
   U1394 : OR2_X1 port map( A1 => n10229, A2 => n10228, ZN => n10242);
   U1395 : NOR3_X1 port map( A1 => n10817, A2 => n10293, A3 => n10591, ZN => 
                           n10234);
   U1396 : NOR2_X1 port map( A1 => n10230, A2 => DATA2(25), ZN => n10773);
   U1397 : INV_X1 port map( A => DATA2(25), ZN => n10902);
   U1398 : NOR2_X1 port map( A1 => n10902, A2 => DATA1(25), ZN => n10777);
   U1399 : NOR2_X1 port map( A1 => n10773, A2 => n10777, ZN => n10611);
   U1400 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n10578, 
                           ZN => n10232);
   U1401 : INV_X1 port map( A => n10253, ZN => n10245);
   U1402 : NAND3_X1 port map( A1 => n10252, A2 => n10236, A3 => n10245, ZN => 
                           n10231);
   U1403 : OAI211_X1 port map( C1 => n10611, C2 => n10594, A => n10232, B => 
                           n10231, ZN => n10233);
   U1404 : AOI211_X1 port map( C1 => dataout_mul_25_port, C2 => n10583, A => 
                           n10234, B => n10233, ZN => n10241);
   U1405 : OAI22_X1 port map( A1 => n10373, A2 => n10235, B1 => n10243, B2 => 
                           n10376, ZN => n10239);
   U1406 : INV_X1 port map( A => n10236, ZN => n10238);
   U1407 : AOI22_X1 port map( A1 => n10438, A2 => n10239, B1 => n10238, B2 => 
                           n10237, ZN => n10240);
   U1408 : OAI211_X1 port map( C1 => n10246, C2 => n10242, A => n10241, B => 
                           n10240, ZN => OUTALU(25));
   U1409 : INV_X1 port map( A => n10601, ZN => n10451);
   U1410 : AOI22_X1 port map( A1 => DATA2(24), A2 => n10451, B1 => 
                           DATA2_I_24_port, B2 => n10252, ZN => n10255);
   U1411 : NOR3_X1 port map( A1 => n10373, A2 => n10243, A3 => n10559, ZN => 
                           n10251);
   U1412 : INV_X1 port map( A => DATA2(24), ZN => n10903);
   U1413 : OAI22_X1 port map( A1 => n10694, A2 => DATA2(24), B1 => n10903, B2 
                           => DATA1(24), ZN => n10690);
   U1414 : INV_X1 port map( A => n10690, ZN => n10770);
   U1415 : OAI22_X1 port map( A1 => n10817, A2 => n10294, B1 => n10293, B2 => 
                           n10818, ZN => n10244);
   U1416 : AOI22_X1 port map( A1 => n10482, A2 => n10244, B1 => n10583, B2 => 
                           dataout_mul_24_port, ZN => n10249);
   U1417 : NAND3_X1 port map( A1 => n10247, A2 => n10246, A3 => n10245, ZN => 
                           n10248);
   U1418 : OAI211_X1 port map( C1 => n10770, C2 => n10594, A => n10249, B => 
                           n10248, ZN => n10250);
   U1419 : AOI211_X1 port map( C1 => n10253, C2 => n10252, A => n10251, B => 
                           n10250, ZN => n10254);
   U1420 : OAI221_X1 port map( B1 => n10694, B2 => n10255, C1 => n10694, C2 => 
                           n10409, A => n10254, ZN => OUTALU(24));
   U1421 : INV_X1 port map( A => DATA2(23), ZN => n10904);
   U1422 : NOR2_X1 port map( A1 => n10256, A2 => n10904, ZN => n10257);
   U1423 : NOR2_X1 port map( A1 => n10256, A2 => DATA2(23), ZN => n10691);
   U1424 : INV_X1 port map( A => n10691, ZN => n10767);
   U1425 : NAND2_X1 port map( A1 => DATA2(23), A2 => n10256, ZN => n10769);
   U1426 : NAND2_X1 port map( A1 => n10767, A2 => n10769, ZN => n10614);
   U1427 : AOI22_X1 port map( A1 => n10257, A2 => n10578, B1 => n10476, B2 => 
                           n10614, ZN => n10283);
   U1428 : OAI222_X1 port map( A1 => n10818, A2 => n10294, B1 => n10814, B2 => 
                           n10293, C1 => n10291, C2 => n10817, ZN => n10258);
   U1429 : AOI22_X1 port map( A1 => n10885, A2 => n10258, B1 => n10583, B2 => 
                           dataout_mul_23_port, ZN => n10282);
   U1430 : OAI22_X1 port map( A1 => n10322, A2 => n10259, B1 => n10285, B2 => 
                           n10304, ZN => n10272);
   U1431 : OAI22_X1 port map( A1 => n10305, A2 => n10863, B1 => n10321, B2 => 
                           n10370, ZN => n10271);
   U1432 : NAND2_X1 port map( A1 => n10268, A2 => n10895, ZN => n10460);
   U1433 : INV_X1 port map( A => n10460, ZN => n10430);
   U1434 : AND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n10261);
   U1435 : NOR2_X1 port map( A1 => n10261, A2 => n10260, ZN => n10405);
   U1436 : OAI21_X1 port map( B1 => n10424, B2 => n10405, A => n10262, ZN => 
                           n10386);
   U1437 : OR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n10263);
   U1438 : OAI21_X1 port map( B1 => n10386, B2 => n10264, A => n10263, ZN => 
                           n10320);
   U1439 : OAI21_X1 port map( B1 => n10330, B2 => n10320, A => n10265, ZN => 
                           n10301);
   U1440 : INV_X1 port map( A => n10301, ZN => n10267);
   U1441 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n10266);
   U1442 : OAI21_X1 port map( B1 => n10267, B2 => n10315, A => n10266, ZN => 
                           n10274);
   U1443 : NOR2_X1 port map( A1 => n1992, A2 => n10268, ZN => n10429);
   U1444 : INV_X1 port map( A => n10276, ZN => n10269);
   U1445 : AOI22_X1 port map( A1 => n10430, A2 => n10274, B1 => n10429, B2 => 
                           n10269, ZN => n10288);
   U1446 : NOR3_X1 port map( A1 => n10278, A2 => n10288, A3 => n10287, ZN => 
                           n10270);
   U1447 : AOI221_X1 port map( B1 => n10272, B2 => n10577, C1 => n10271, C2 => 
                           n10438, A => n10270, ZN => n10281);
   U1448 : INV_X1 port map( A => n10273, ZN => n10279);
   U1449 : NOR2_X1 port map( A1 => n10460, A2 => n10274, ZN => n10275);
   U1450 : AOI211_X1 port map( C1 => n10276, C2 => n10429, A => n10275, B => 
                           n10287, ZN => n10286);
   U1451 : OAI21_X1 port map( B1 => n10279, B2 => n10286, A => n10278, ZN => 
                           n10277);
   U1452 : OAI211_X1 port map( C1 => n10279, C2 => n10278, A => n10895, B => 
                           n10277, ZN => n10280);
   U1453 : NAND4_X1 port map( A1 => n10283, A2 => n10282, A3 => n10281, A4 => 
                           n10280, ZN => OUTALU(23));
   U1454 : INV_X1 port map( A => DATA2(22), ZN => n10905);
   U1455 : OAI22_X1 port map( A1 => n10768, A2 => DATA2(22), B1 => n10905, B2 
                           => DATA1(22), ZN => n10763);
   U1456 : AOI22_X1 port map( A1 => dataout_mul_22_port, A2 => n10602, B1 => 
                           n10476, B2 => n10763, ZN => n10300);
   U1457 : OAI222_X1 port map( A1 => n10863, A2 => n10321, B1 => n10304, B2 => 
                           n10305, C1 => n10285, C2 => n10284, ZN => n10290);
   U1458 : AOI21_X1 port map( B1 => n10288, B2 => n10287, A => n10286, ZN => 
                           n10289);
   U1459 : AOI21_X1 port map( B1 => n10438, B2 => n10290, A => n10289, ZN => 
                           n10299);
   U1460 : OAI22_X1 port map( A1 => n10817, A2 => n10292, B1 => n10291, B2 => 
                           n10818, ZN => n10296);
   U1461 : OAI22_X1 port map( A1 => n10294, A2 => n10814, B1 => n10293, B2 => 
                           n10820, ZN => n10295);
   U1462 : OAI21_X1 port map( B1 => n10296, B2 => n10295, A => n10885, ZN => 
                           n10298);
   U1463 : NAND3_X1 port map( A1 => DATA2(22), A2 => DATA1(22), A3 => n10578, 
                           ZN => n10297);
   U1464 : NAND4_X1 port map( A1 => n10300, A2 => n10299, A3 => n10298, A4 => 
                           n10297, ZN => OUTALU(22));
   U1465 : AOI22_X1 port map( A1 => n10430, A2 => n10301, B1 => n10429, B2 => 
                           n10302, ZN => n10316);
   U1466 : INV_X1 port map( A => n10429, ZN => n10458);
   U1467 : OAI22_X1 port map( A1 => n10302, A2 => n10458, B1 => n10460, B2 => 
                           n10301, ZN => n10303);
   U1468 : INV_X1 port map( A => n10303, ZN => n10314);
   U1469 : OAI22_X1 port map( A1 => n10322, A2 => n10305, B1 => n10321, B2 => 
                           n10304, ZN => n10312);
   U1470 : INV_X1 port map( A => n10409, ZN => n10450);
   U1471 : AOI21_X1 port map( B1 => n10451, B2 => DATA2(21), A => n10450, ZN =>
                           n10310);
   U1472 : NOR3_X1 port map( A1 => n10391, A2 => n10591, A3 => n10826, ZN => 
                           n10306);
   U1473 : AOI21_X1 port map( B1 => dataout_mul_21_port, B2 => n10583, A => 
                           n10306, ZN => n10308);
   U1474 : NOR2_X1 port map( A1 => DATA2(21), A2 => n10309, ZN => n10686);
   U1475 : INV_X1 port map( A => DATA2(21), ZN => n10906);
   U1476 : NOR2_X1 port map( A1 => n10906, A2 => DATA1(21), ZN => n10764);
   U1477 : OAI21_X1 port map( B1 => n10686, B2 => n10764, A => n10556, ZN => 
                           n10307);
   U1478 : OAI211_X1 port map( C1 => n10310, C2 => n10309, A => n10308, B => 
                           n10307, ZN => n10311);
   U1479 : AOI21_X1 port map( B1 => n10577, B2 => n10312, A => n10311, ZN => 
                           n10313);
   U1480 : OAI221_X1 port map( B1 => n10317, B2 => n10316, C1 => n10315, C2 => 
                           n10314, A => n10313, ZN => OUTALU(21));
   U1481 : INV_X1 port map( A => n10330, ZN => n10332);
   U1482 : OAI22_X1 port map( A1 => n10319, A2 => n10458, B1 => n10460, B2 => 
                           n10320, ZN => n10318);
   U1483 : INV_X1 port map( A => n10318, ZN => n10331);
   U1484 : AOI22_X1 port map( A1 => n10430, A2 => n10320, B1 => n10429, B2 => 
                           n10319, ZN => n10329);
   U1485 : INV_X1 port map( A => DATA2(20), ZN => n10907);
   U1486 : OAI21_X1 port map( B1 => n10601, B2 => n10907, A => n10409, ZN => 
                           n10327);
   U1487 : NOR3_X1 port map( A1 => n10322, A2 => n10321, A3 => n10559, ZN => 
                           n10326);
   U1488 : NOR2_X1 port map( A1 => n10907, A2 => DATA1(20), ZN => n10616);
   U1489 : INV_X1 port map( A => n10616, ZN => n10759);
   U1490 : NAND2_X1 port map( A1 => n10907, A2 => DATA1(20), ZN => n10682);
   U1491 : OAI22_X1 port map( A1 => n10390, A2 => n10826, B1 => n10391, B2 => 
                           n10831, ZN => n10323);
   U1492 : AOI22_X1 port map( A1 => n10885, A2 => n10323, B1 => n10602, B2 => 
                           dataout_mul_20_port, ZN => n10324);
   U1493 : OAI221_X1 port map( B1 => n10594, B2 => n10759, C1 => n10594, C2 => 
                           n10682, A => n10324, ZN => n10325);
   U1494 : AOI211_X1 port map( C1 => DATA1(20), C2 => n10327, A => n10326, B =>
                           n10325, ZN => n10328);
   U1495 : OAI221_X1 port map( B1 => n10332, B2 => n10331, C1 => n10330, C2 => 
                           n10329, A => n10328, ZN => OUTALU(20));
   U1496 : NOR2_X1 port map( A1 => n10333, A2 => n10645, ZN => n10334);
   U1497 : AOI22_X1 port map( A1 => n10583, A2 => dataout_mul_1_port, B1 => 
                           n10577, B2 => n10334, ZN => n10385);
   U1498 : NOR2_X1 port map( A1 => n10335, A2 => DATA2(1), ZN => n10648);
   U1499 : INV_X1 port map( A => n10648, ZN => n10712);
   U1500 : NOR2_X1 port map( A1 => n10928, A2 => DATA1(1), ZN => n10714);
   U1501 : INV_X1 port map( A => n10714, ZN => n10646);
   U1502 : NAND2_X1 port map( A1 => n10712, A2 => n10646, ZN => n10643);
   U1503 : AOI221_X1 port map( B1 => n10337, B2 => n10336, C1 => n10593, C2 => 
                           n10340, A => n10596, ZN => n10343);
   U1504 : AOI211_X1 port map( C1 => n10341, C2 => n10340, A => n10339, B => 
                           n10338, ZN => n10342);
   U1505 : AOI211_X1 port map( C1 => n10556, C2 => n10643, A => n10343, B => 
                           n10342, ZN => n10384);
   U1506 : AOI21_X1 port map( B1 => n10577, B2 => n10344, A => n10450, ZN => 
                           n10600);
   U1507 : OAI21_X1 port map( B1 => n10928, B2 => n10601, A => n10600, ZN => 
                           n10382);
   U1508 : INV_X1 port map( A => n10879, ZN => n10380);
   U1509 : AOI22_X1 port map( A1 => n10803, A2 => DATA1(2), B1 => n10802, B2 =>
                           DATA1(1), ZN => n10348);
   U1510 : NAND4_X1 port map( A1 => n10348, A2 => n10347, A3 => n10346, A4 => 
                           n10345, ZN => n10813);
   U1511 : AOI222_X1 port map( A1 => n10811, A2 => n10812, B1 => n10350, B2 => 
                           n10810, C1 => n10813, C2 => n10349, ZN => n10819);
   U1512 : OAI22_X1 port map( A1 => n10817, A2 => n10819, B1 => n10821, B2 => 
                           n10814, ZN => n10354);
   U1513 : OAI22_X1 port map( A1 => n10352, A2 => n10351, B1 => n10815, B2 => 
                           n10818, ZN => n10353);
   U1514 : AOI211_X1 port map( C1 => n10355, C2 => n10824, A => n10354, B => 
                           n10353, ZN => n10832);
   U1515 : OAI22_X1 port map( A1 => n10801, A2 => n10828, B1 => n10832, B2 => 
                           n10826, ZN => n10359);
   U1516 : INV_X1 port map( A => n10356, ZN => n10829);
   U1517 : OAI22_X1 port map( A1 => n10834, A2 => n10357, B1 => n10829, B2 => 
                           n10831, ZN => n10358);
   U1518 : AOI211_X1 port map( C1 => n10838, C2 => n10830, A => n10359, B => 
                           n10358, ZN => n10843);
   U1519 : OAI222_X1 port map( A1 => n10844, A2 => n10840, B1 => n10842, B2 => 
                           n10843, C1 => n10360, C2 => n10839, ZN => n10851);
   U1520 : AOI22_X1 port map( A1 => n10848, A2 => n10851, B1 => n10846, B2 => 
                           n10800, ZN => n10363);
   U1521 : AOI22_X1 port map( A1 => n10852, A2 => n10845, B1 => n10849, B2 => 
                           n10361, ZN => n10362);
   U1522 : OAI211_X1 port map( C1 => n10364, C2 => n10855, A => n10363, B => 
                           n10362, ZN => n10798);
   U1523 : AOI22_X1 port map( A1 => n10365, A2 => n10859, B1 => n10858, B2 => 
                           n10798, ZN => n10369);
   U1524 : AOI22_X1 port map( A1 => n10569, A2 => n10367, B1 => n10797, B2 => 
                           n10366, ZN => n10368);
   U1525 : OAI211_X1 port map( C1 => n10371, C2 => n10370, A => n10369, B => 
                           n10368, ZN => n10869);
   U1526 : INV_X1 port map( A => n10869, ZN => n10372);
   U1527 : OAI222_X1 port map( A1 => n10376, A2 => n10865, B1 => n10375, B2 => 
                           n10374, C1 => n10373, C2 => n10372, ZN => n10874);
   U1528 : AOI22_X1 port map( A1 => n10377, A2 => n10874, B1 => n10877, B2 => 
                           n10878, ZN => n10379);
   U1529 : AOI22_X1 port map( A1 => n10875, A2 => n10872, B1 => n10873, B2 => 
                           n10876, ZN => n10378);
   U1530 : OAI211_X1 port map( C1 => n10381, C2 => n10380, A => n10379, B => 
                           n10378, ZN => n10888);
   U1531 : AOI22_X1 port map( A1 => DATA1(1), A2 => n10382, B1 => n10482, B2 =>
                           n10888, ZN => n10383);
   U1532 : NAND3_X1 port map( A1 => n10385, A2 => n10384, A3 => n10383, ZN => 
                           OUTALU(1));
   U1533 : INV_X1 port map( A => n10401, ZN => n10403);
   U1534 : AOI22_X1 port map( A1 => n10430, A2 => n10386, B1 => n10429, B2 => 
                           n10387, ZN => n10402);
   U1535 : OAI22_X1 port map( A1 => n10387, A2 => n10458, B1 => n10460, B2 => 
                           n10386, ZN => n10388);
   U1536 : INV_X1 port map( A => n10388, ZN => n10400);
   U1537 : OAI22_X1 port map( A1 => n10389, A2 => n10448, B1 => n10407, B2 => 
                           n10431, ZN => n10398);
   U1538 : OAI22_X1 port map( A1 => n10432, A2 => n10408, B1 => n10449, B2 => 
                           n10855, ZN => n10397);
   U1539 : INV_X1 port map( A => n10390, ZN => n10410);
   U1540 : INV_X1 port map( A => n10391, ZN => n10413);
   U1541 : AOI222_X1 port map( A1 => n10410, A2 => n10554, B1 => n10413, B2 => 
                           n10525, C1 => n10411, C2 => n10576, ZN => n10395);
   U1542 : NOR2_X1 port map( A1 => n10392, A2 => DATA2(19), ZN => n10762);
   U1543 : INV_X1 port map( A => n10762, ZN => n10683);
   U1544 : NAND2_X1 port map( A1 => DATA2(19), A2 => n10392, ZN => n10760);
   U1545 : NAND2_X1 port map( A1 => n10683, A2 => n10760, ZN => n10642);
   U1546 : AOI22_X1 port map( A1 => dataout_mul_19_port, A2 => n10602, B1 => 
                           n10476, B2 => n10642, ZN => n10394);
   U1547 : NAND3_X1 port map( A1 => DATA2(19), A2 => DATA1(19), A3 => n10578, 
                           ZN => n10393);
   U1548 : OAI211_X1 port map( C1 => n10395, C2 => n10591, A => n10394, B => 
                           n10393, ZN => n10396);
   U1549 : AOI221_X1 port map( B1 => n10398, B2 => n10577, C1 => n10397, C2 => 
                           n10438, A => n10396, ZN => n10399);
   U1550 : OAI221_X1 port map( B1 => n10403, B2 => n10402, C1 => n10401, C2 => 
                           n10400, A => n10399, ZN => OUTALU(19));
   U1551 : INV_X1 port map( A => n10424, ZN => n10426);
   U1552 : OAI22_X1 port map( A1 => n10460, A2 => n10405, B1 => n10458, B2 => 
                           n10406, ZN => n10404);
   U1553 : INV_X1 port map( A => n10404, ZN => n10425);
   U1554 : AOI22_X1 port map( A1 => n10406, A2 => n10429, B1 => n10430, B2 => 
                           n10405, ZN => n10423);
   U1555 : OAI222_X1 port map( A1 => n10431, A2 => n10432, B1 => n10408, B2 => 
                           n10449, C1 => n10448, C2 => n10407, ZN => n10421);
   U1556 : INV_X1 port map( A => DATA1(18), ZN => n10415);
   U1557 : INV_X1 port map( A => DATA2(18), ZN => n10909);
   U1558 : AOI211_X1 port map( C1 => n10409, C2 => n10601, A => n10415, B => 
                           n10909, ZN => n10420);
   U1559 : AOI22_X1 port map( A1 => n10554, A2 => n10411, B1 => n10525, B2 => 
                           n10410, ZN => n10418);
   U1560 : AOI22_X1 port map( A1 => n10414, A2 => n10413, B1 => n10576, B2 => 
                           n10412, ZN => n10417);
   U1561 : NOR2_X1 port map( A1 => n10909, A2 => DATA1(18), ZN => n10758);
   U1562 : INV_X1 port map( A => n10758, ZN => n10681);
   U1563 : NOR2_X1 port map( A1 => n10415, A2 => DATA2(18), ZN => n10679);
   U1564 : INV_X1 port map( A => n10679, ZN => n10756);
   U1565 : NAND2_X1 port map( A1 => n10681, A2 => n10756, ZN => n10607);
   U1566 : AOI22_X1 port map( A1 => dataout_mul_18_port, A2 => n10602, B1 => 
                           n10476, B2 => n10607, ZN => n10416);
   U1567 : OAI221_X1 port map( B1 => n10591, B2 => n10418, C1 => n10591, C2 => 
                           n10417, A => n10416, ZN => n10419);
   U1568 : AOI211_X1 port map( C1 => n10438, C2 => n10421, A => n10420, B => 
                           n10419, ZN => n10422);
   U1569 : OAI221_X1 port map( B1 => n10426, B2 => n10425, C1 => n10424, C2 => 
                           n10423, A => n10422, ZN => OUTALU(18));
   U1570 : OAI22_X1 port map( A1 => n10428, A2 => n10458, B1 => n10460, B2 => 
                           n10444, ZN => n10427);
   U1571 : INV_X1 port map( A => n10427, ZN => n10442);
   U1572 : AOI22_X1 port map( A1 => n10430, A2 => n10444, B1 => n10429, B2 => 
                           n10428, ZN => n10440);
   U1573 : OAI22_X1 port map( A1 => n10432, A2 => n10448, B1 => n10449, B2 => 
                           n10431, ZN => n10437);
   U1574 : NOR3_X1 port map( A1 => n10446, A2 => n10591, A3 => n10842, ZN => 
                           n10436);
   U1575 : NAND3_X1 port map( A1 => n10578, A2 => DATA2(17), A3 => DATA1(17), 
                           ZN => n10434);
   U1576 : INV_X1 port map( A => DATA2(17), ZN => n10910);
   U1577 : NAND2_X1 port map( A1 => DATA1(17), A2 => n10910, ZN => n10678);
   U1578 : OR2_X1 port map( A1 => n10910, A2 => DATA1(17), ZN => n10754);
   U1579 : NAND2_X1 port map( A1 => n10678, A2 => n10754, ZN => n10606);
   U1580 : AOI22_X1 port map( A1 => dataout_mul_17_port, A2 => n10602, B1 => 
                           n10476, B2 => n10606, ZN => n10433);
   U1581 : NAND2_X1 port map( A1 => n10434, A2 => n10433, ZN => n10435);
   U1582 : AOI211_X1 port map( C1 => n10438, C2 => n10437, A => n10436, B => 
                           n10435, ZN => n10439);
   U1583 : OAI221_X1 port map( B1 => n10443, B2 => n10442, C1 => n10441, C2 => 
                           n10440, A => n10439, ZN => OUTALU(17));
   U1584 : NOR2_X1 port map( A1 => n10445, A2 => n10444, ZN => n10461);
   U1585 : INV_X1 port map( A => n10461, ZN => n10459);
   U1586 : OAI22_X1 port map( A1 => n10447, A2 => n10842, B1 => n10446, B2 => 
                           n10844, ZN => n10456);
   U1587 : NOR3_X1 port map( A1 => n10449, A2 => n10559, A3 => n10448, ZN => 
                           n10455);
   U1588 : AOI21_X1 port map( B1 => n10451, B2 => DATA2(16), A => n10450, ZN =>
                           n10453);
   U1589 : NOR2_X1 port map( A1 => DATA2(16), A2 => n10675, ZN => n10755);
   U1590 : AOI21_X1 port map( B1 => DATA2(16), B2 => n10675, A => n10755, ZN =>
                           n10622);
   U1591 : INV_X1 port map( A => n10622, ZN => n10749);
   U1592 : AOI22_X1 port map( A1 => dataout_mul_16_port, A2 => n10602, B1 => 
                           n10476, B2 => n10749, ZN => n10452);
   U1593 : OAI21_X1 port map( B1 => n10453, B2 => n10675, A => n10452, ZN => 
                           n10454);
   U1594 : AOI211_X1 port map( C1 => n10885, C2 => n10456, A => n10455, B => 
                           n10454, ZN => n10457);
   U1595 : OAI221_X1 port map( B1 => n10461, B2 => n10460, C1 => n10459, C2 => 
                           n10458, A => n10457, ZN => OUTALU(16));
   U1596 : AOI22_X1 port map( A1 => n10488, A2 => n10463, B1 => n10462, B2 => 
                           n10487, ZN => n10485);
   U1597 : XOR2_X1 port map( A => n10464, B => n10473, Z => n10481);
   U1598 : INV_X1 port map( A => n10465, ZN => n10570);
   U1599 : INV_X1 port map( A => n10466, ZN => n10571);
   U1600 : OAI21_X1 port map( B1 => n10570, B2 => n10588, A => n10571, ZN => 
                           n10585);
   U1601 : NAND2_X1 port map( A1 => n10467, A2 => n10585, ZN => n10547);
   U1602 : INV_X1 port map( A => n10547, ZN => n10469);
   U1603 : OAI21_X1 port map( B1 => n10470, B2 => n10469, A => n10468, ZN => 
                           n10535);
   U1604 : AOI21_X1 port map( B1 => n10472, B2 => n10535, A => n10471, ZN => 
                           n10496);
   U1605 : NAND2_X1 port map( A1 => n10496, A2 => n10495, ZN => n10493);
   U1606 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n10499, B2 => n10493, ZN => n10474);
   U1607 : XNOR2_X1 port map( A => n10474, B => n10473, ZN => n10479);
   U1608 : NOR2_X1 port map( A1 => n10475, A2 => DATA2(15), ZN => n10745);
   U1609 : INV_X1 port map( A => DATA2(15), ZN => n10912);
   U1610 : NOR2_X1 port map( A1 => n10912, A2 => n11229, ZN => n10750);
   U1611 : OR2_X1 port map( A1 => n10745, A2 => n10750, ZN => n10604);
   U1612 : AOI22_X1 port map( A1 => dataout_mul_15_port, A2 => n10602, B1 => 
                           n10476, B2 => n10604, ZN => n10478);
   U1613 : NAND3_X1 port map( A1 => DATA2(15), A2 => n11229, A3 => n10578, ZN 
                           => n10477);
   U1614 : OAI211_X1 port map( C1 => n10479, C2 => n10565, A => n10478, B => 
                           n10477, ZN => n10480);
   U1615 : AOI21_X1 port map( B1 => n10548, B2 => n10481, A => n10480, ZN => 
                           n10484);
   U1616 : NAND3_X1 port map( A1 => n10482, A2 => n10848, A3 => n10530, ZN => 
                           n10483);
   U1617 : OAI211_X1 port map( C1 => n10485, C2 => n10559, A => n10484, B => 
                           n10483, ZN => OUTALU(15));
   U1618 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           ZN => n11159);
   U1619 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           A => n11159, ZN => n11160);
   U1620 : NOR3_X1 port map( A1 => n5126, A2 => n5134, A3 => n11160, ZN => 
                           n3087);
   U1621 : AOI22_X1 port map( A1 => n10848, A2 => n10529, B1 => n10527, B2 => 
                           n10530, ZN => n10506);
   U1622 : AOI221_X1 port map( B1 => n5134, B2 => n5126, C1 => n11160, C2 => 
                           n5126, A => n3087, ZN => n10504);
   U1623 : NAND3_X1 port map( A1 => DATA2(14), A2 => DATA1(14), A3 => n10578, 
                           ZN => n10491);
   U1624 : NAND2_X1 port map( A1 => n10486, A2 => DATA2(14), ZN => n10672);
   U1625 : INV_X1 port map( A => n10672, ZN => n10620);
   U1626 : NOR2_X1 port map( A1 => n10486, A2 => DATA2(14), ZN => n10746);
   U1627 : OAI21_X1 port map( B1 => n10620, B2 => n10746, A => n10556, ZN => 
                           n10490);
   U1628 : NAND3_X1 port map( A1 => n10577, A2 => n10488, A3 => n10487, ZN => 
                           n10489);
   U1629 : NAND3_X1 port map( A1 => n10491, A2 => n10490, A3 => n10489, ZN => 
                           n10503);
   U1630 : AOI22_X1 port map( A1 => n10586, A2 => n10493, B1 => n10548, B2 => 
                           n10492, ZN => n10494);
   U1631 : INV_X1 port map( A => n10494, ZN => n10501);
   U1632 : INV_X1 port map( A => n10495, ZN => n10498);
   U1633 : AOI22_X1 port map( A1 => n10497, A2 => n10548, B1 => n10586, B2 => 
                           n10496, ZN => n10523);
   U1634 : NOR2_X1 port map( A1 => n10498, A2 => n10523, ZN => n10500);
   U1635 : MUX2_X1 port map( A => n10501, B => n10500, S => n10499, Z => n10502
                           );
   U1636 : AOI211_X1 port map( C1 => n10583, C2 => n10504, A => n10503, B => 
                           n10502, ZN => n10505);
   U1637 : OAI21_X1 port map( B1 => n10506, B2 => n10591, A => n10505, ZN => 
                           OUTALU(14));
   U1638 : AOI22_X1 port map( A1 => n10554, A2 => n10524, B1 => n10576, B2 => 
                           n10507, ZN => n10508);
   U1639 : OAI21_X1 port map( B1 => n10509, B2 => n10828, A => n10508, ZN => 
                           n10510);
   U1640 : AOI21_X1 port map( B1 => n10838, B2 => n10575, A => n10510, ZN => 
                           n10514);
   U1641 : NOR2_X1 port map( A1 => n10511, A2 => DATA2(13), ZN => n10741);
   U1642 : NOR2_X1 port map( A1 => DATA1(13), A2 => n10914, ZN => n10669);
   U1643 : OAI21_X1 port map( B1 => n10741, B2 => n10669, A => n10556, ZN => 
                           n10513);
   U1644 : NAND3_X1 port map( A1 => DATA2(13), A2 => DATA1(13), A3 => n10578, 
                           ZN => n10512);
   U1645 : OAI211_X1 port map( C1 => n10514, C2 => n10559, A => n10513, B => 
                           n10512, ZN => n10519);
   U1646 : AOI222_X1 port map( A1 => n10526, A2 => n10848, B1 => n10529, B2 => 
                           n10527, C1 => n10530, C2 => n10846, ZN => n10517);
   U1647 : INV_X1 port map( A => n10542, ZN => n10540);
   U1648 : NAND2_X1 port map( A1 => n10540, A2 => n10535, ZN => n10534);
   U1649 : OAI211_X1 port map( C1 => n10541, C2 => n10515, A => n10895, B => 
                           n10521, ZN => n10516);
   U1650 : OAI22_X1 port map( A1 => n10517, A2 => n10591, B1 => n10534, B2 => 
                           n10516, ZN => n10518);
   U1651 : AOI211_X1 port map( C1 => n10583, C2 => dataout_mul_13_port, A => 
                           n10519, B => n10518, ZN => n10520);
   U1652 : OAI221_X1 port map( B1 => n10523, B2 => n10522, C1 => n10523, C2 => 
                           n10521, A => n10520, ZN => OUTALU(13));
   U1653 : AOI222_X1 port map( A1 => n10553, A2 => n10554, B1 => n10575, B2 => 
                           n10525, C1 => n10524, C2 => n10576, ZN => n10546);
   U1654 : AOI22_X1 port map( A1 => n10848, A2 => n10528, B1 => n10527, B2 => 
                           n10526, ZN => n10533);
   U1655 : AOI22_X1 port map( A1 => n10531, A2 => n10530, B1 => n10846, B2 => 
                           n10529, ZN => n10532);
   U1656 : AOI21_X1 port map( B1 => n10533, B2 => n10532, A => n10591, ZN => 
                           n10539);
   U1657 : OAI22_X1 port map( A1 => n10744, A2 => DATA2(12), B1 => n10915, B2 
                           => DATA1(12), ZN => n10665);
   U1658 : INV_X1 port map( A => n10665, ZN => n10738);
   U1659 : OAI211_X1 port map( C1 => n10540, C2 => n10535, A => n10586, B => 
                           n10534, ZN => n10537);
   U1660 : NAND3_X1 port map( A1 => DATA2(12), A2 => DATA1(12), A3 => n10578, 
                           ZN => n10536);
   U1661 : OAI211_X1 port map( C1 => n10738, C2 => n10594, A => n10537, B => 
                           n10536, ZN => n10538);
   U1662 : AOI211_X1 port map( C1 => n10583, C2 => dataout_mul_12_port, A => 
                           n10539, B => n10538, ZN => n10545);
   U1663 : INV_X1 port map( A => n10541, ZN => n10543);
   U1664 : OAI221_X1 port map( B1 => n10543, B2 => n10542, C1 => n10541, C2 => 
                           n10540, A => n10548, ZN => n10544);
   U1665 : OAI211_X1 port map( C1 => n10546, C2 => n10559, A => n10545, B => 
                           n10544, ZN => OUTALU(12));
   U1666 : INV_X1 port map( A => n10551, ZN => n10549);
   U1667 : XNOR2_X1 port map( A => n10549, B => n10547, ZN => n10566);
   U1668 : INV_X1 port map( A => n10552, ZN => n10550);
   U1669 : INV_X1 port map( A => n10548, ZN => n10572);
   U1670 : AOI221_X1 port map( B1 => n10552, B2 => n10551, C1 => n10550, C2 => 
                           n10549, A => n10572, ZN => n10562);
   U1671 : AOI22_X1 port map( A1 => n10554, A2 => n10575, B1 => n10576, B2 => 
                           n10553, ZN => n10560);
   U1672 : NAND3_X1 port map( A1 => DATA2(11), A2 => n11228, A3 => n10578, ZN 
                           => n10558);
   U1673 : NOR2_X1 port map( A1 => DATA2(11), A2 => n10555, ZN => n10666);
   U1674 : NAND2_X1 port map( A1 => n10555, A2 => DATA2(11), ZN => n10737);
   U1675 : INV_X1 port map( A => n10737, ZN => n10627);
   U1676 : OAI21_X1 port map( B1 => n10666, B2 => n10627, A => n10556, ZN => 
                           n10557);
   U1677 : OAI211_X1 port map( C1 => n10560, C2 => n10559, A => n10558, B => 
                           n10557, ZN => n10561);
   U1678 : AOI211_X1 port map( C1 => n10583, C2 => dataout_mul_11_port, A => 
                           n10562, B => n10561, ZN => n10564);
   U1679 : NAND3_X1 port map( A1 => n10885, A2 => n10858, A3 => n10568, ZN => 
                           n10563);
   U1680 : OAI211_X1 port map( C1 => n10566, C2 => n10565, A => n10564, B => 
                           n10563, ZN => OUTALU(11));
   U1681 : AOI22_X1 port map( A1 => n10569, A2 => n10568, B1 => n10858, B2 => 
                           n10567, ZN => n10592);
   U1682 : NOR2_X1 port map( A1 => n10571, A2 => n10570, ZN => n10584);
   U1683 : AOI211_X1 port map( C1 => n10584, C2 => n10574, A => n10573, B => 
                           n10572, ZN => n10582);
   U1684 : OAI22_X1 port map( A1 => n10628, A2 => DATA2(10), B1 => n10917, B2 
                           => DATA1(10), ZN => n10734);
   U1685 : INV_X1 port map( A => n10734, ZN => n10662);
   U1686 : NAND3_X1 port map( A1 => n10577, A2 => n10576, A3 => n10575, ZN => 
                           n10580);
   U1687 : NAND3_X1 port map( A1 => DATA2(10), A2 => DATA1(10), A3 => n10578, 
                           ZN => n10579);
   U1688 : OAI211_X1 port map( C1 => n10662, C2 => n10594, A => n10580, B => 
                           n10579, ZN => n10581);
   U1689 : AOI211_X1 port map( C1 => n10583, C2 => dataout_mul_10_port, A => 
                           n10582, B => n10581, ZN => n10590);
   U1690 : INV_X1 port map( A => n10584, ZN => n10587);
   U1691 : OAI211_X1 port map( C1 => n10588, C2 => n10587, A => n10586, B => 
                           n10585, ZN => n10589);
   U1692 : OAI211_X1 port map( C1 => n10592, C2 => n10591, A => n10590, B => 
                           n10589, ZN => OUTALU(10));
   U1693 : OAI21_X1 port map( B1 => DATA1(0), B2 => DATA2_I_0_port, A => n10593
                           , ZN => n10598);
   U1694 : OAI22_X1 port map( A1 => n10929, A2 => n10645, B1 => DATA1(0), B2 =>
                           DATA2(0), ZN => n10610);
   U1695 : OR2_X1 port map( A1 => n10594, A2 => n10610, ZN => n10595);
   U1696 : OAI21_X1 port map( B1 => n10596, B2 => n10598, A => n10595, ZN => 
                           n10597);
   U1697 : AOI21_X1 port map( B1 => n10599, B2 => n10598, A => n10597, ZN => 
                           n10893);
   U1698 : OAI21_X1 port map( B1 => n10929, B2 => n10601, A => n10600, ZN => 
                           n10603);
   U1699 : AOI22_X1 port map( A1 => DATA1(0), A2 => n10603, B1 => n10602, B2 =>
                           dataout_mul_0_port, ZN => n10892);
   U1700 : NOR4_X1 port map( A1 => n10607, A2 => n10606, A3 => n10605, A4 => 
                           n10604, ZN => n10608);
   U1701 : NAND4_X1 port map( A1 => FUNC(2), A2 => n10610, A3 => n10609, A4 => 
                           n10608, ZN => n10641);
   U1702 : INV_X1 port map( A => n10611, ZN => n10615);
   U1703 : NOR4_X1 port map( A1 => n10615, A2 => n10614, A3 => n10613, A4 => 
                           n10612, ZN => n10639);
   U1704 : OR2_X1 port map( A1 => n10741, A2 => n10746, ZN => n10673);
   U1705 : NOR2_X1 port map( A1 => n10616, A2 => n10764, ZN => n10688);
   U1706 : INV_X1 port map( A => n10688, ZN => n10619);
   U1707 : NOR4_X1 port map( A1 => n10673, A2 => n10619, A3 => n10618, A4 => 
                           n10617, ZN => n10638);
   U1708 : NOR2_X1 port map( A1 => n10669, A2 => n10620, ZN => n10748);
   U1709 : INV_X1 port map( A => n10682, ZN => n10621);
   U1710 : NOR2_X1 port map( A1 => n10686, A2 => n10621, ZN => n10766);
   U1711 : NAND4_X1 port map( A1 => n10738, A2 => n10748, A3 => n10622, A4 => 
                           n10766, ZN => n10636);
   U1712 : INV_X1 port map( A => n10719, ZN => n10625);
   U1713 : INV_X1 port map( A => n10649, ZN => n10623);
   U1714 : NAND2_X1 port map( A1 => n10623, A2 => n10652, ZN => n10722);
   U1715 : AOI21_X1 port map( B1 => DATA1(10), B2 => n10917, A => n10666, ZN =>
                           n10624);
   U1716 : INV_X1 port map( A => n10624, ZN => n10739);
   U1717 : OR4_X1 port map( A1 => n10625, A2 => n10722, A3 => n10727, A4 => 
                           n10739, ZN => n10635);
   U1718 : INV_X1 port map( A => n10701, ZN => n10788);
   U1719 : INV_X1 port map( A => n10716, ZN => n10626);
   U1720 : NAND2_X1 port map( A1 => n10626, A2 => n10721, ZN => n10653);
   U1721 : INV_X1 port map( A => n10653, ZN => n10630);
   U1722 : AOI21_X1 port map( B1 => DATA2(10), B2 => n10628, A => n10627, ZN =>
                           n10668);
   U1723 : NAND4_X1 port map( A1 => n10788, A2 => n10630, A3 => n10629, A4 => 
                           n10668, ZN => n10634);
   U1724 : INV_X1 port map( A => n10631, ZN => n10632);
   U1725 : OR4_X1 port map( A1 => n10763, A2 => n10690, A3 => n10632, A4 => 
                           n10698, ZN => n10633);
   U1726 : NOR4_X1 port map( A1 => n10636, A2 => n10635, A3 => n10634, A4 => 
                           n10633, ZN => n10637);
   U1727 : NAND3_X1 port map( A1 => n10639, A2 => n10638, A3 => n10637, ZN => 
                           n10640);
   U1728 : NOR4_X1 port map( A1 => n10643, A2 => n10642, A3 => n10641, A4 => 
                           n10640, ZN => n10709);
   U1729 : NOR2_X1 port map( A1 => n10755, A2 => n10745, ZN => n10677);
   U1730 : NOR2_X1 port map( A1 => DATA2(6), A2 => n10644, ZN => n10658);
   U1731 : NAND2_X1 port map( A1 => DATA2(0), A2 => n10645, ZN => n10647);
   U1732 : OAI21_X1 port map( B1 => n10648, B2 => n10647, A => n10646, ZN => 
                           n10651);
   U1733 : NOR2_X1 port map( A1 => DATA1(2), A2 => n10927, ZN => n10650);
   U1734 : AOI211_X1 port map( C1 => n10719, C2 => n10651, A => n10650, B => 
                           n10649, ZN => n10654);
   U1735 : OAI211_X1 port map( C1 => n10654, C2 => n10653, A => n10652, B => 
                           n10724, ZN => n10655);
   U1736 : NAND2_X1 port map( A1 => n10720, A2 => n10655, ZN => n10657);
   U1737 : INV_X1 port map( A => n10728, ZN => n10656);
   U1738 : OAI211_X1 port map( C1 => n10658, C2 => n10657, A => n10725, B => 
                           n10656, ZN => n10659);
   U1739 : OAI21_X1 port map( B1 => DATA2(8), B2 => n10710, A => n10659, ZN => 
                           n10661);
   U1740 : OAI22_X1 port map( A1 => n10711, A2 => n10661, B1 => n10660, B2 => 
                           n10919, ZN => n10663);
   U1741 : OAI211_X1 port map( C1 => n10664, C2 => n10663, A => n10662, B => 
                           n10736, ZN => n10667);
   U1742 : AOI211_X1 port map( C1 => n10668, C2 => n10667, A => n10666, B => 
                           n10665, ZN => n10670);
   U1743 : AOI211_X1 port map( C1 => DATA2(12), C2 => n10744, A => n10670, B =>
                           n10669, ZN => n10674);
   U1744 : INV_X1 port map( A => n10750, ZN => n10671);
   U1745 : OAI211_X1 port map( C1 => n10674, C2 => n10673, A => n10672, B => 
                           n10671, ZN => n10676);
   U1746 : AOI22_X1 port map( A1 => n10677, A2 => n10676, B1 => DATA2(16), B2 
                           => n10675, ZN => n10680);
   U1747 : INV_X1 port map( A => n10678, ZN => n10752);
   U1748 : AOI211_X1 port map( C1 => n10680, C2 => n10754, A => n10752, B => 
                           n10679, ZN => n10685);
   U1749 : NAND2_X1 port map( A1 => n10681, A2 => n10760, ZN => n10684);
   U1750 : OAI211_X1 port map( C1 => n10685, C2 => n10684, A => n10683, B => 
                           n10682, ZN => n10687);
   U1751 : AOI211_X1 port map( C1 => n10688, C2 => n10687, A => n10686, B => 
                           n10763, ZN => n10689);
   U1752 : AOI21_X1 port map( B1 => DATA2(22), B2 => n10768, A => n10689, ZN =>
                           n10692);
   U1753 : AOI211_X1 port map( C1 => n10692, C2 => n10769, A => n10691, B => 
                           n10690, ZN => n10693);
   U1754 : AOI21_X1 port map( B1 => DATA2(24), B2 => n10694, A => n10693, ZN =>
                           n10696);
   U1755 : INV_X1 port map( A => n10777, ZN => n10695);
   U1756 : AOI211_X1 port map( C1 => n10696, C2 => n10695, A => n10780, B => 
                           n10773, ZN => n10697);
   U1757 : AOI21_X1 port map( B1 => DATA2(26), B2 => n10778, A => n10697, ZN =>
                           n10699);
   U1758 : AOI211_X1 port map( C1 => n10699, C2 => n10783, A => n10779, B => 
                           n10698, ZN => n10700);
   U1759 : AOI21_X1 port map( B1 => DATA2(28), B2 => n10784, A => n10700, ZN =>
                           n10702);
   U1760 : AOI211_X1 port map( C1 => n10702, C2 => n10787, A => n10790, B => 
                           n10701, ZN => n10704);
   U1761 : AOI211_X1 port map( C1 => DATA2(30), C2 => n10793, A => n10704, B =>
                           n10703, ZN => n10705);
   U1762 : NOR4_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => n10706, A4 => 
                           n10705, ZN => n10708);
   U1763 : NOR4_X1 port map( A1 => FUNC(1), A2 => n10709, A3 => n10708, A4 => 
                           n10707, ZN => n10887);
   U1764 : NAND2_X1 port map( A1 => DATA1(24), A2 => n10903, ZN => n10776);
   U1765 : NOR2_X1 port map( A1 => DATA2(8), A2 => n10710, ZN => n10733);
   U1766 : INV_X1 port map( A => DATA2(6), ZN => n10923);
   U1767 : AOI21_X1 port map( B1 => DATA1(6), B2 => n10923, A => n10711, ZN => 
                           n10730);
   U1768 : NAND2_X1 port map( A1 => DATA1(0), A2 => n10929, ZN => n10713);
   U1769 : OAI21_X1 port map( B1 => n10714, B2 => n10713, A => n10712, ZN => 
                           n10718);
   U1770 : NOR2_X1 port map( A1 => DATA2(2), A2 => n10715, ZN => n10717);
   U1771 : AOI211_X1 port map( C1 => n10719, C2 => n10718, A => n10717, B => 
                           n10716, ZN => n10723);
   U1772 : OAI211_X1 port map( C1 => n10723, C2 => n10722, A => n10721, B => 
                           n10720, ZN => n10726);
   U1773 : NAND3_X1 port map( A1 => n10726, A2 => n10725, A3 => n10724, ZN => 
                           n10729);
   U1774 : AOI211_X1 port map( C1 => n10730, C2 => n10729, A => n10728, B => 
                           n10727, ZN => n10732);
   U1775 : OAI21_X1 port map( B1 => n10733, B2 => n10732, A => n10731, ZN => 
                           n10735);
   U1776 : AOI21_X1 port map( B1 => n10736, B2 => n10735, A => n10734, ZN => 
                           n10740);
   U1777 : OAI211_X1 port map( C1 => n10740, C2 => n10739, A => n10738, B => 
                           n10737, ZN => n10743);
   U1778 : INV_X1 port map( A => n10741, ZN => n10742);
   U1779 : OAI211_X1 port map( C1 => DATA2(12), C2 => n10744, A => n10743, B =>
                           n10742, ZN => n10747);
   U1780 : AOI211_X1 port map( C1 => n10748, C2 => n10747, A => n10746, B => 
                           n10745, ZN => n10751);
   U1781 : NOR3_X1 port map( A1 => n10751, A2 => n10750, A3 => n10749, ZN => 
                           n10753);
   U1782 : AOI221_X1 port map( B1 => n10755, B2 => n10754, C1 => n10753, C2 => 
                           n10754, A => n10752, ZN => n10757);
   U1783 : OAI21_X1 port map( B1 => n10758, B2 => n10757, A => n10756, ZN => 
                           n10761);
   U1784 : OAI211_X1 port map( C1 => n10762, C2 => n10761, A => n10760, B => 
                           n10759, ZN => n10765);
   U1785 : AOI211_X1 port map( C1 => n10766, C2 => n10765, A => n10764, B => 
                           n10763, ZN => n10772);
   U1786 : OAI21_X1 port map( B1 => DATA2(22), B2 => n10768, A => n10767, ZN =>
                           n10771);
   U1787 : OAI211_X1 port map( C1 => n10772, C2 => n10771, A => n10770, B => 
                           n10769, ZN => n10775);
   U1788 : INV_X1 port map( A => n10773, ZN => n10774);
   U1789 : OAI221_X1 port map( B1 => n10777, B2 => n10776, C1 => n10777, C2 => 
                           n10775, A => n10774, ZN => n10782);
   U1790 : NAND2_X1 port map( A1 => DATA2(26), A2 => n10778, ZN => n10781);
   U1791 : AOI211_X1 port map( C1 => n10782, C2 => n10781, A => n10780, B => 
                           n10779, ZN => n10786);
   U1792 : OAI21_X1 port map( B1 => DATA1(28), B2 => n10899, A => n10783, ZN =>
                           n10785);
   U1793 : OAI22_X1 port map( A1 => n10786, A2 => n10785, B1 => DATA2(28), B2 
                           => n10784, ZN => n10789);
   U1794 : OAI211_X1 port map( C1 => n10790, C2 => n10789, A => n10788, B => 
                           n10787, ZN => n10792);
   U1795 : OAI211_X1 port map( C1 => DATA2(30), C2 => n10793, A => n10792, B =>
                           n10791, ZN => n10794);
   U1796 : OAI221_X1 port map( B1 => FUNC(2), B2 => n10795, C1 => FUNC(2), C2 
                           => n10794, A => FUNC(3), ZN => n10886);
   U1797 : AOI22_X1 port map( A1 => n10799, A2 => n10798, B1 => n10797, B2 => 
                           n10796, ZN => n10862);
   U1798 : INV_X1 port map( A => n10800, ZN => n10856);
   U1799 : INV_X1 port map( A => n10801, ZN => n10837);
   U1800 : AOI22_X1 port map( A1 => n10803, A2 => DATA1(1), B1 => n10802, B2 =>
                           DATA1(0), ZN => n10807);
   U1801 : NAND4_X1 port map( A1 => n10807, A2 => n10806, A3 => n10805, A4 => 
                           n10804, ZN => n10809);
   U1802 : AOI222_X1 port map( A1 => n10813, A2 => n10812, B1 => n10811, B2 => 
                           n10810, C1 => n10809, C2 => n10808, ZN => n10816);
   U1803 : OAI22_X1 port map( A1 => n10817, A2 => n10816, B1 => n10815, B2 => 
                           n10814, ZN => n10823);
   U1804 : OAI22_X1 port map( A1 => n10821, A2 => n10820, B1 => n10819, B2 => 
                           n10818, ZN => n10822);
   U1805 : AOI211_X1 port map( C1 => n10825, C2 => n10824, A => n10823, B => 
                           n10822, ZN => n10827);
   U1806 : OAI22_X1 port map( A1 => n10829, A2 => n10828, B1 => n10827, B2 => 
                           n10826, ZN => n10836);
   U1807 : INV_X1 port map( A => n10830, ZN => n10833);
   U1808 : OAI22_X1 port map( A1 => n10834, A2 => n10833, B1 => n10832, B2 => 
                           n10831, ZN => n10835);
   U1809 : AOI211_X1 port map( C1 => n10838, C2 => n10837, A => n10836, B => 
                           n10835, ZN => n10841);
   U1810 : OAI222_X1 port map( A1 => n10844, A2 => n10843, B1 => n10842, B2 => 
                           n10841, C1 => n10840, C2 => n10839, ZN => n10847);
   U1811 : AOI22_X1 port map( A1 => n10848, A2 => n10847, B1 => n10846, B2 => 
                           n10845, ZN => n10854);
   U1812 : AOI22_X1 port map( A1 => n10852, A2 => n10851, B1 => n10850, B2 => 
                           n10849, ZN => n10853);
   U1813 : OAI211_X1 port map( C1 => n10856, C2 => n10855, A => n10854, B => 
                           n10853, ZN => n10857);
   U1814 : AOI22_X1 port map( A1 => n10860, A2 => n10859, B1 => n10858, B2 => 
                           n10857, ZN => n10861);
   U1815 : OAI211_X1 port map( C1 => n10864, C2 => n10863, A => n10862, B => 
                           n10861, ZN => n10871);
   U1816 : INV_X1 port map( A => n10865, ZN => n10867);
   U1817 : AOI222_X1 port map( A1 => n10871, A2 => n10870, B1 => n10869, B2 => 
                           n10868, C1 => n10867, C2 => n10866, ZN => n10883);
   U1818 : AOI22_X1 port map( A1 => n10875, A2 => n10874, B1 => n10873, B2 => 
                           n10872, ZN => n10881);
   U1819 : AOI22_X1 port map( A1 => n10879, A2 => n10878, B1 => n10877, B2 => 
                           n10876, ZN => n10880);
   U1820 : OAI211_X1 port map( C1 => n10883, C2 => n10882, A => n10881, B => 
                           n10880, ZN => n10884);
   U1821 : AOI22_X1 port map( A1 => n10887, A2 => n10886, B1 => n10885, B2 => 
                           n10884, ZN => n10891);
   U1822 : NAND4_X1 port map( A1 => FUNC(2), A2 => FUNC(3), A3 => n10889, A4 =>
                           n10888, ZN => n10890);
   U1823 : NAND4_X1 port map( A1 => n10893, A2 => n10892, A3 => n10891, A4 => 
                           n10890, ZN => OUTALU(0));
   U1824 : NAND2_X1 port map( A1 => n10895, A2 => n10894, ZN => n10931);
   U1825 : CLKBUF_X1 port map( A => n10931, Z => n10921);
   U1826 : NAND2_X1 port map( A1 => FUNC(3), A2 => n10895, ZN => n10930);
   U1827 : CLKBUF_X1 port map( A => n10930, Z => n10920);
   U1828 : AOI22_X1 port map( A1 => DATA2(31), A2 => n10921, B1 => n10920, B2 
                           => n10896, ZN => N2548);
   U1829 : AOI22_X1 port map( A1 => DATA2(30), A2 => n10931, B1 => n10930, B2 
                           => n10897, ZN => N2547);
   U1830 : INV_X1 port map( A => DATA2(29), ZN => n10898);
   U1831 : AOI22_X1 port map( A1 => DATA2(29), A2 => n10921, B1 => n10920, B2 
                           => n10898, ZN => N2546);
   U1832 : AOI22_X1 port map( A1 => DATA2(28), A2 => n10931, B1 => n10930, B2 
                           => n10899, ZN => N2545);
   U1833 : INV_X1 port map( A => DATA2(27), ZN => n10900);
   U1834 : AOI22_X1 port map( A1 => DATA2(27), A2 => n10921, B1 => n10920, B2 
                           => n10900, ZN => N2544);
   U1835 : INV_X1 port map( A => DATA2(26), ZN => n10901);
   U1836 : AOI22_X1 port map( A1 => DATA2(26), A2 => n10931, B1 => n10930, B2 
                           => n10901, ZN => N2543);
   U1837 : AOI22_X1 port map( A1 => DATA2(25), A2 => n10921, B1 => n10920, B2 
                           => n10902, ZN => N2542);
   U1838 : AOI22_X1 port map( A1 => DATA2(24), A2 => n10931, B1 => n10930, B2 
                           => n10903, ZN => N2541);
   U1839 : AOI22_X1 port map( A1 => DATA2(23), A2 => n10921, B1 => n10920, B2 
                           => n10904, ZN => N2540);
   U1840 : AOI22_X1 port map( A1 => DATA2(22), A2 => n10931, B1 => n10930, B2 
                           => n10905, ZN => N2539);
   U1841 : AOI22_X1 port map( A1 => DATA2(21), A2 => n10931, B1 => n10930, B2 
                           => n10906, ZN => N2538);
   U1842 : AOI22_X1 port map( A1 => DATA2(20), A2 => n10931, B1 => n10930, B2 
                           => n10907, ZN => N2537);
   U1843 : INV_X1 port map( A => DATA2(19), ZN => n10908);
   U1844 : AOI22_X1 port map( A1 => DATA2(19), A2 => n10921, B1 => n10920, B2 
                           => n10908, ZN => N2536);
   U1845 : AOI22_X1 port map( A1 => DATA2(18), A2 => n10921, B1 => n10920, B2 
                           => n10909, ZN => N2535);
   U1846 : AOI22_X1 port map( A1 => DATA2(17), A2 => n10921, B1 => n10920, B2 
                           => n10910, ZN => N2534);
   U1847 : INV_X1 port map( A => DATA2(16), ZN => n10911);
   U1848 : AOI22_X1 port map( A1 => DATA2(16), A2 => n10921, B1 => n10920, B2 
                           => n10911, ZN => N2533);
   U1849 : AOI22_X1 port map( A1 => DATA2(15), A2 => n10921, B1 => n10920, B2 
                           => n10912, ZN => N2532);
   U1850 : INV_X1 port map( A => DATA2(14), ZN => n10913);
   U1851 : AOI22_X1 port map( A1 => DATA2(14), A2 => n10921, B1 => n10920, B2 
                           => n10913, ZN => N2531);
   U1852 : AOI22_X1 port map( A1 => DATA2(13), A2 => n10921, B1 => n10920, B2 
                           => n10914, ZN => N2530);
   U1853 : AOI22_X1 port map( A1 => DATA2(12), A2 => n10921, B1 => n10920, B2 
                           => n10915, ZN => N2529);
   U1854 : AOI22_X1 port map( A1 => DATA2(11), A2 => n10921, B1 => n10920, B2 
                           => n10916, ZN => N2528);
   U1855 : AOI22_X1 port map( A1 => DATA2(10), A2 => n10921, B1 => n10920, B2 
                           => n10917, ZN => N2527);
   U1856 : AOI22_X1 port map( A1 => DATA2(9), A2 => n10921, B1 => n10920, B2 =>
                           n10918, ZN => N2526);
   U1857 : AOI22_X1 port map( A1 => DATA2(8), A2 => n10921, B1 => n10920, B2 =>
                           n10919, ZN => N2525);
   U1858 : AOI22_X1 port map( A1 => DATA2(7), A2 => n10931, B1 => n10930, B2 =>
                           n10922, ZN => N2524);
   U1859 : AOI22_X1 port map( A1 => DATA2(6), A2 => n10931, B1 => n10930, B2 =>
                           n10923, ZN => N2523);
   U1860 : AOI22_X1 port map( A1 => DATA2(5), A2 => n10931, B1 => n10930, B2 =>
                           n10924, ZN => N2522);
   U1861 : AOI22_X1 port map( A1 => DATA2(4), A2 => n10931, B1 => n10930, B2 =>
                           n10925, ZN => N2521);
   U1862 : AOI22_X1 port map( A1 => DATA2(3), A2 => n10931, B1 => n10930, B2 =>
                           n10926, ZN => N2520);
   U1863 : AOI22_X1 port map( A1 => DATA2(2), A2 => n10931, B1 => n10930, B2 =>
                           n10927, ZN => N2519);
   U1864 : AOI22_X1 port map( A1 => DATA2(1), A2 => n10931, B1 => n10930, B2 =>
                           n10928, ZN => N2518);
   U1865 : AOI22_X1 port map( A1 => DATA2(0), A2 => n10931, B1 => n10930, B2 =>
                           n10929, ZN => N2517);
   U1866 : NOR2_X1 port map( A1 => n10932, A2 => n2024, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1867 : NAND2_X1 port map( A1 => n10973, A2 => data2_mul_3_port, ZN => 
                           n10936);
   U1868 : INV_X1 port map( A => data2_mul_3_port, ZN => n10969);
   U1869 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n10969, ZN => n10968);
   U1870 : INV_X1 port map( A => n10933, ZN => n10934);
   U1871 : NOR2_X1 port map( A1 => n10934, A2 => n10969, ZN => n10971);
   U1872 : NOR2_X1 port map( A1 => data2_mul_3_port, A2 => n10934, ZN => n10961
                           );
   U1873 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n10971, B1 => data1_mul_1_port, B2 => n10961, 
                           ZN => n10935);
   U1874 : OAI221_X1 port map( B1 => n2024, B2 => n10936, C1 => n2024, C2 => 
                           n10968, A => n10935, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1875 : INV_X1 port map( A => n10936, ZN => n10970);
   U1876 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n10961, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n10970, ZN => n10938);
   U1877 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n10971, ZN => n10937);
   U1878 : OAI211_X1 port map( C1 => n2023, C2 => n10968, A => n10938, B => 
                           n10937, ZN => boothmul_pipelined_i_mux_out_1_4_port)
                           ;
   U1879 : CLKBUF_X1 port map( A => n10961, Z => n10965);
   U1880 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n10970, B1 => n10965, B2 => data1_mul_3_port, 
                           ZN => n10940);
   U1881 : CLKBUF_X1 port map( A => n10971, Z => n10962);
   U1882 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n10939);
   U1883 : OAI211_X1 port map( C1 => n10968, C2 => n2021, A => n10940, B => 
                           n10939, ZN => boothmul_pipelined_i_mux_out_1_5_port)
                           ;
   U1884 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n10965, B2 => data1_mul_4_port, ZN => n10942);
   U1885 : NAND2_X1 port map( A1 => n10971, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n10941);
   U1886 : OAI211_X1 port map( C1 => n2020, C2 => n10968, A => n10942, B => 
                           n10941, ZN => boothmul_pipelined_i_mux_out_1_6_port)
                           ;
   U1887 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n10965, B2 => data1_mul_5_port, ZN => n10944);
   U1888 : NAND2_X1 port map( A1 => n10971, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n10943);
   U1889 : OAI211_X1 port map( C1 => n2018, C2 => n10968, A => n10944, B => 
                           n10943, ZN => boothmul_pipelined_i_mux_out_1_7_port)
                           ;
   U1890 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n10965, B2 => data1_mul_6_port, ZN => n10946);
   U1891 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n10945);
   U1892 : OAI211_X1 port map( C1 => n2016, C2 => n10968, A => n10946, B => 
                           n10945, ZN => boothmul_pipelined_i_mux_out_1_8_port)
                           ;
   U1893 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n10961, B2 => data1_mul_7_port, ZN => n10948);
   U1894 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n10947);
   U1895 : OAI211_X1 port map( C1 => n2014, C2 => n10968, A => n10948, B => 
                           n10947, ZN => boothmul_pipelined_i_mux_out_1_9_port)
                           ;
   U1896 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n10961, B2 => data1_mul_8_port, ZN => n10950);
   U1897 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n10949);
   U1898 : OAI211_X1 port map( C1 => n2012, C2 => n10968, A => n10950, B => 
                           n10949, ZN => boothmul_pipelined_i_mux_out_1_10_port
                           );
   U1899 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n10965, B2 => data1_mul_9_port, ZN => n10952);
   U1900 : NAND2_X1 port map( A1 => n10971, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n10951);
   U1901 : OAI211_X1 port map( C1 => n2010, C2 => n10968, A => n10952, B => 
                           n10951, ZN => boothmul_pipelined_i_mux_out_1_11_port
                           );
   U1902 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n10961, B2 => data1_mul_10_port, ZN => n10954);
   U1903 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n10953);
   U1904 : OAI211_X1 port map( C1 => n2008, C2 => n10968, A => n10954, B => 
                           n10953, ZN => boothmul_pipelined_i_mux_out_1_12_port
                           );
   U1905 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n10965, B2 => data1_mul_11_port, ZN => n10956);
   U1906 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n10955);
   U1907 : OAI211_X1 port map( C1 => n2006, C2 => n10968, A => n10956, B => 
                           n10955, ZN => boothmul_pipelined_i_mux_out_1_13_port
                           );
   U1908 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n10965, B2 => data1_mul_12_port, ZN => n10958);
   U1909 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n10957);
   U1910 : OAI211_X1 port map( C1 => n2004, C2 => n10968, A => n10958, B => 
                           n10957, ZN => boothmul_pipelined_i_mux_out_1_14_port
                           );
   U1911 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n10961, B2 => data1_mul_13_port, ZN => n10960);
   U1912 : NAND2_X1 port map( A1 => n10971, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n10959);
   U1913 : OAI211_X1 port map( C1 => n2002, C2 => n10968, A => n10960, B => 
                           n10959, ZN => boothmul_pipelined_i_mux_out_1_15_port
                           );
   U1914 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n10961, B2 => data1_mul_14_port, ZN => n10964);
   U1915 : NAND2_X1 port map( A1 => n10962, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n10963);
   U1916 : OAI211_X1 port map( C1 => n2000, C2 => n10968, A => n10964, B => 
                           n10963, ZN => boothmul_pipelined_i_mux_out_1_16_port
                           );
   U1917 : AOI22_X1 port map( A1 => n10970, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n10965, B2 => data1_mul_15_port, ZN => n10967);
   U1918 : NAND2_X1 port map( A1 => n10971, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n10966);
   U1919 : OAI211_X1 port map( C1 => n1998, C2 => n10968, A => n10967, B => 
                           n10966, ZN => boothmul_pipelined_i_mux_out_1_17_port
                           );
   U1920 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n10969, ZN => 
                           n10974);
   U1921 : AOI22_X1 port map( A1 => n10971, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n10970, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n10972);
   U1922 : OAI21_X1 port map( B1 => n10974, B2 => n10973, A => n10972, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1923 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n11013);
   U1924 : NAND2_X1 port map( A1 => n11013, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n10977);
   U1925 : NAND3_X1 port map( A1 => n3076, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n11009);
   U1926 : NOR2_X1 port map( A1 => n3076, A2 => n10975, ZN => n10990);
   U1927 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n10975, ZN => n11003);
   U1928 : CLKBUF_X1 port map( A => n11003, Z => n11006);
   U1929 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n10990, B1 => data1_mul_1_port, B2 => n11006, 
                           ZN => n10976);
   U1930 : OAI221_X1 port map( B1 => n2024, B2 => n10977, C1 => n2024, C2 => 
                           n11009, A => n10976, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1931 : INV_X1 port map( A => n10977, ZN => n11011);
   U1932 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n11003, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n11011, ZN => n10979);
   U1933 : CLKBUF_X1 port map( A => n10990, Z => n11010);
   U1934 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n11010, ZN => n10978);
   U1935 : OAI211_X1 port map( C1 => n11009, C2 => n2023, A => n10979, B => 
                           n10978, ZN => boothmul_pipelined_i_mux_out_2_6_port)
                           ;
   U1936 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n11011, B1 => data1_mul_3_port, B2 => n11006, 
                           ZN => n10981);
   U1937 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n10990, ZN => n10980);
   U1938 : OAI211_X1 port map( C1 => n11009, C2 => n2021, A => n10981, B => 
                           n10980, ZN => boothmul_pipelined_i_mux_out_2_7_port)
                           ;
   U1939 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n11011, B1 => data1_mul_4_port, B2 => n11006, 
                           ZN => n10983);
   U1940 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n10990, ZN => n10982);
   U1941 : OAI211_X1 port map( C1 => n11009, C2 => n2020, A => n10983, B => 
                           n10982, ZN => boothmul_pipelined_i_mux_out_2_8_port)
                           ;
   U1942 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n11011, B1 => data1_mul_5_port, B2 => n11003, 
                           ZN => n10985);
   U1943 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n10990, ZN => n10984);
   U1944 : OAI211_X1 port map( C1 => n11009, C2 => n2018, A => n10985, B => 
                           n10984, ZN => boothmul_pipelined_i_mux_out_2_9_port)
                           ;
   U1945 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n11011, B1 => data1_mul_6_port, B2 => n11006, 
                           ZN => n10987);
   U1946 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n10990, ZN => n10986);
   U1947 : OAI211_X1 port map( C1 => n11009, C2 => n2016, A => n10987, B => 
                           n10986, ZN => boothmul_pipelined_i_mux_out_2_10_port
                           );
   U1948 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n11011, B1 => data1_mul_7_port, B2 => n11003, 
                           ZN => n10989);
   U1949 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n10990, ZN => n10988);
   U1950 : OAI211_X1 port map( C1 => n11009, C2 => n2014, A => n10989, B => 
                           n10988, ZN => boothmul_pipelined_i_mux_out_2_11_port
                           );
   U1951 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n11011, B1 => data1_mul_8_port, B2 => n11006, 
                           ZN => n10992);
   U1952 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n10990, ZN => n10991);
   U1953 : OAI211_X1 port map( C1 => n11009, C2 => n2012, A => n10992, B => 
                           n10991, ZN => boothmul_pipelined_i_mux_out_2_12_port
                           );
   U1954 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n11011, B1 => data1_mul_9_port, B2 => n11006, 
                           ZN => n10994);
   U1955 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n11010, ZN => n10993);
   U1956 : OAI211_X1 port map( C1 => n11009, C2 => n2010, A => n10994, B => 
                           n10993, ZN => boothmul_pipelined_i_mux_out_2_13_port
                           );
   U1957 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n11011, B1 => data1_mul_10_port, B2 => n11003,
                           ZN => n10996);
   U1958 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n11010, ZN => n10995);
   U1959 : OAI211_X1 port map( C1 => n11009, C2 => n2008, A => n10996, B => 
                           n10995, ZN => boothmul_pipelined_i_mux_out_2_14_port
                           );
   U1960 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n11011, B1 => data1_mul_11_port, B2 => n11003,
                           ZN => n10998);
   U1961 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n11010, ZN => n10997);
   U1962 : OAI211_X1 port map( C1 => n11009, C2 => n2006, A => n10998, B => 
                           n10997, ZN => boothmul_pipelined_i_mux_out_2_15_port
                           );
   U1963 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n11011, B1 => data1_mul_12_port, B2 => n11006,
                           ZN => n11000);
   U1964 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n11010, ZN => n10999);
   U1965 : OAI211_X1 port map( C1 => n11009, C2 => n2004, A => n11000, B => 
                           n10999, ZN => boothmul_pipelined_i_mux_out_2_16_port
                           );
   U1966 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n11011, B1 => data1_mul_13_port, B2 => n11003,
                           ZN => n11002);
   U1967 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n11010, ZN => n11001);
   U1968 : OAI211_X1 port map( C1 => n11009, C2 => n2002, A => n11002, B => 
                           n11001, ZN => boothmul_pipelined_i_mux_out_2_17_port
                           );
   U1969 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n11011, B1 => data1_mul_14_port, B2 => n11003,
                           ZN => n11005);
   U1970 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n11010, ZN => n11004);
   U1971 : OAI211_X1 port map( C1 => n11009, C2 => n2000, A => n11005, B => 
                           n11004, ZN => boothmul_pipelined_i_mux_out_2_18_port
                           );
   U1972 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n11011, B1 => data1_mul_15_port, B2 => n11006,
                           ZN => n11008);
   U1973 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n11010, ZN => n11007);
   U1974 : OAI211_X1 port map( C1 => n11009, C2 => n1998, A => n11008, B => 
                           n11007, ZN => boothmul_pipelined_i_mux_out_2_19_port
                           );
   U1975 : NAND2_X1 port map( A1 => n3076, A2 => data1_mul_15_port, ZN => 
                           n11014);
   U1976 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n11011, B1 => n11010, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n11012);
   U1977 : OAI21_X1 port map( B1 => n11014, B2 => n11013, A => n11012, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1978 : NAND3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n11224);
   U1979 : NOR3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n11222);
   U1980 : INV_X1 port map( A => n11222, ZN => n11018);
   U1981 : INV_X1 port map( A => n11016, ZN => n11015);
   U1982 : NAND2_X1 port map( A1 => n3082, A2 => n11015, ZN => n11225);
   U1983 : INV_X1 port map( A => n11225, ZN => n11044);
   U1984 : NOR2_X1 port map( A1 => n3082, A2 => n11016, ZN => n11048);
   U1985 : CLKBUF_X1 port map( A => n11048, Z => n11221);
   U1986 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n11017);
   U1987 : OAI221_X1 port map( B1 => n3077, B2 => n11224, C1 => n3077, C2 => 
                           n11018, A => n11017, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1988 : INV_X1 port map( A => n11224, ZN => n11047);
   U1989 : CLKBUF_X1 port map( A => n11222, Z => n11043);
   U1990 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_3_60_port, A2
                           => n11047, B1 => n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n11020);
   U1991 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => 
                           n11048, B2 => 
                           boothmul_pipelined_i_muxes_in_3_175_port, ZN => 
                           n11019);
   U1992 : NAND2_X1 port map( A1 => n11020, A2 => n11019, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1993 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => 
                           n11222, B2 => 
                           boothmul_pipelined_i_muxes_in_3_175_port, ZN => 
                           n11022);
   U1994 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => 
                           n11048, B2 => 
                           boothmul_pipelined_i_muxes_in_3_174_port, ZN => 
                           n11021);
   U1995 : NAND2_X1 port map( A1 => n11022, A2 => n11021, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1996 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => 
                           n11222, B2 => 
                           boothmul_pipelined_i_muxes_in_3_174_port, ZN => 
                           n11024);
   U1997 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => 
                           n11048, B2 => 
                           boothmul_pipelined_i_muxes_in_3_173_port, ZN => 
                           n11023);
   U1998 : NAND2_X1 port map( A1 => n11024, A2 => n11023, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1999 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_173_port, ZN => 
                           n11026);
   U2000 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_172_port, ZN => 
                           n11025);
   U2001 : NAND2_X1 port map( A1 => n11026, A2 => n11025, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U2002 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_172_port, ZN => 
                           n11028);
   U2003 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => 
                           n11048, B2 => 
                           boothmul_pipelined_i_muxes_in_3_171_port, ZN => 
                           n11027);
   U2004 : NAND2_X1 port map( A1 => n11028, A2 => n11027, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U2005 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_171_port, ZN => 
                           n11030);
   U2006 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_170_port, ZN => 
                           n11029);
   U2007 : NAND2_X1 port map( A1 => n11030, A2 => n11029, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U2008 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_170_port, ZN => 
                           n11032);
   U2009 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_169_port, ZN => 
                           n11031);
   U2010 : NAND2_X1 port map( A1 => n11032, A2 => n11031, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U2011 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_169_port, ZN => 
                           n11034);
   U2012 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_168_port, ZN => 
                           n11033);
   U2013 : NAND2_X1 port map( A1 => n11034, A2 => n11033, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U2014 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_168_port, ZN => 
                           n11036);
   U2015 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => 
                           n11048, B2 => 
                           boothmul_pipelined_i_muxes_in_3_167_port, ZN => 
                           n11035);
   U2016 : NAND2_X1 port map( A1 => n11036, A2 => n11035, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U2017 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_167_port, ZN => 
                           n11038);
   U2018 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_166_port, ZN => 
                           n11037);
   U2019 : NAND2_X1 port map( A1 => n11038, A2 => n11037, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U2020 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_166_port, ZN => 
                           n11040);
   U2021 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_165_port, ZN => 
                           n11039);
   U2022 : NAND2_X1 port map( A1 => n11040, A2 => n11039, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U2023 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => 
                           n11222, B2 => 
                           boothmul_pipelined_i_muxes_in_3_165_port, ZN => 
                           n11042);
   U2024 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_164_port, ZN => 
                           n11041);
   U2025 : NAND2_X1 port map( A1 => n11042, A2 => n11041, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U2026 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => 
                           n11043, B2 => 
                           boothmul_pipelined_i_muxes_in_3_164_port, ZN => 
                           n11046);
   U2027 : AOI22_X1 port map( A1 => n11044, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => 
                           n11048, B2 => 
                           boothmul_pipelined_i_muxes_in_3_163_port, ZN => 
                           n11045);
   U2028 : NAND2_X1 port map( A1 => n11046, A2 => n11045, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U2029 : AOI22_X1 port map( A1 => n11047, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => 
                           n11222, B2 => 
                           boothmul_pipelined_i_muxes_in_3_163_port, ZN => 
                           n11050);
   U2030 : NAND2_X1 port map( A1 => n11048, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, ZN => 
                           n11049);
   U2031 : OAI211_X1 port map( C1 => n7164, C2 => n11225, A => n11050, B => 
                           n11049, ZN => boothmul_pipelined_i_mux_out_3_21_port
                           );
   U2032 : NAND3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n11209);
   U2033 : NOR3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n11207);
   U2034 : INV_X1 port map( A => n11207, ZN => n11054);
   U2035 : INV_X1 port map( A => n11052, ZN => n11051);
   U2036 : NAND2_X1 port map( A1 => n3078, A2 => n11051, ZN => n11210);
   U2037 : INV_X1 port map( A => n11210, ZN => n11080);
   U2038 : NOR2_X1 port map( A1 => n3078, A2 => n11052, ZN => n11084);
   U2039 : CLKBUF_X1 port map( A => n11084, Z => n11206);
   U2040 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n11053);
   U2041 : OAI221_X1 port map( B1 => n5121, B2 => n11209, C1 => n5121, C2 => 
                           n11054, A => n11053, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U2042 : INV_X1 port map( A => n11209, ZN => n11083);
   U2043 : CLKBUF_X1 port map( A => n11207, Z => n11079);
   U2044 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_64_port, A2
                           => n11083, B1 => n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n11056);
   U2045 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => 
                           n11084, B2 => 
                           boothmul_pipelined_i_muxes_in_4_189_port, ZN => 
                           n11055);
   U2046 : NAND2_X1 port map( A1 => n11056, A2 => n11055, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U2047 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => 
                           n11207, B2 => 
                           boothmul_pipelined_i_muxes_in_4_189_port, ZN => 
                           n11058);
   U2048 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => 
                           n11084, B2 => 
                           boothmul_pipelined_i_muxes_in_4_188_port, ZN => 
                           n11057);
   U2049 : NAND2_X1 port map( A1 => n11058, A2 => n11057, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U2050 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => 
                           n11207, B2 => 
                           boothmul_pipelined_i_muxes_in_4_188_port, ZN => 
                           n11060);
   U2051 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => 
                           n11084, B2 => 
                           boothmul_pipelined_i_muxes_in_4_187_port, ZN => 
                           n11059);
   U2052 : NAND2_X1 port map( A1 => n11060, A2 => n11059, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2053 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_187_port, ZN => 
                           n11062);
   U2054 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_186_port, ZN => 
                           n11061);
   U2055 : NAND2_X1 port map( A1 => n11062, A2 => n11061, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2056 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_186_port, ZN => 
                           n11064);
   U2057 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => 
                           n11084, B2 => 
                           boothmul_pipelined_i_muxes_in_4_185_port, ZN => 
                           n11063);
   U2058 : NAND2_X1 port map( A1 => n11064, A2 => n11063, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2059 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_185_port, ZN => 
                           n11066);
   U2060 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_184_port, ZN => 
                           n11065);
   U2061 : NAND2_X1 port map( A1 => n11066, A2 => n11065, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2062 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_184_port, ZN => 
                           n11068);
   U2063 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_183_port, ZN => 
                           n11067);
   U2064 : NAND2_X1 port map( A1 => n11068, A2 => n11067, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2065 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_183_port, ZN => 
                           n11070);
   U2066 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_182_port, ZN => 
                           n11069);
   U2067 : NAND2_X1 port map( A1 => n11070, A2 => n11069, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2068 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_182_port, ZN => 
                           n11072);
   U2069 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => 
                           n11084, B2 => 
                           boothmul_pipelined_i_muxes_in_4_181_port, ZN => 
                           n11071);
   U2070 : NAND2_X1 port map( A1 => n11072, A2 => n11071, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2071 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_181_port, ZN => 
                           n11074);
   U2072 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_180_port, ZN => 
                           n11073);
   U2073 : NAND2_X1 port map( A1 => n11074, A2 => n11073, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2074 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_180_port, ZN => 
                           n11076);
   U2075 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_179_port, ZN => 
                           n11075);
   U2076 : NAND2_X1 port map( A1 => n11076, A2 => n11075, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2077 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => 
                           n11207, B2 => 
                           boothmul_pipelined_i_muxes_in_4_179_port, ZN => 
                           n11078);
   U2078 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_178_port, ZN => 
                           n11077);
   U2079 : NAND2_X1 port map( A1 => n11078, A2 => n11077, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2080 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => 
                           n11079, B2 => 
                           boothmul_pipelined_i_muxes_in_4_178_port, ZN => 
                           n11082);
   U2081 : AOI22_X1 port map( A1 => n11080, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => 
                           n11084, B2 => 
                           boothmul_pipelined_i_muxes_in_4_177_port, ZN => 
                           n11081);
   U2082 : NAND2_X1 port map( A1 => n11082, A2 => n11081, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2083 : AOI22_X1 port map( A1 => n11083, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => 
                           n11207, B2 => 
                           boothmul_pipelined_i_muxes_in_4_177_port, ZN => 
                           n11086);
   U2084 : NAND2_X1 port map( A1 => n11084, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, ZN => 
                           n11085);
   U2085 : OAI211_X1 port map( C1 => n5127, C2 => n11210, A => n11086, B => 
                           n11085, ZN => boothmul_pipelined_i_mux_out_4_23_port
                           );
   U2086 : NAND3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n11214);
   U2087 : NOR3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n11212);
   U2088 : INV_X1 port map( A => n11212, ZN => n11090);
   U2089 : INV_X1 port map( A => n11088, ZN => n11087);
   U2090 : NAND2_X1 port map( A1 => n3079, A2 => n11087, ZN => n11215);
   U2091 : INV_X1 port map( A => n11215, ZN => n11116);
   U2092 : NOR2_X1 port map( A1 => n3079, A2 => n11088, ZN => n11120);
   U2093 : CLKBUF_X1 port map( A => n11120, Z => n11211);
   U2094 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n11089);
   U2095 : OAI221_X1 port map( B1 => n5122, B2 => n11214, C1 => n5122, C2 => 
                           n11090, A => n11089, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2096 : INV_X1 port map( A => n11214, ZN => n11119);
   U2097 : CLKBUF_X1 port map( A => n11212, Z => n11115);
   U2098 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_5_68_port, A2
                           => n11119, B1 => n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n11092);
   U2099 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => 
                           n11120, B2 => 
                           boothmul_pipelined_i_muxes_in_5_203_port, ZN => 
                           n11091);
   U2100 : NAND2_X1 port map( A1 => n11092, A2 => n11091, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2101 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => 
                           n11212, B2 => 
                           boothmul_pipelined_i_muxes_in_5_203_port, ZN => 
                           n11094);
   U2102 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => 
                           n11120, B2 => 
                           boothmul_pipelined_i_muxes_in_5_202_port, ZN => 
                           n11093);
   U2103 : NAND2_X1 port map( A1 => n11094, A2 => n11093, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2104 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => 
                           n11212, B2 => 
                           boothmul_pipelined_i_muxes_in_5_202_port, ZN => 
                           n11096);
   U2105 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => 
                           n11120, B2 => 
                           boothmul_pipelined_i_muxes_in_5_201_port, ZN => 
                           n11095);
   U2106 : NAND2_X1 port map( A1 => n11096, A2 => n11095, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2107 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_201_port, ZN => 
                           n11098);
   U2108 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_200_port, ZN => 
                           n11097);
   U2109 : NAND2_X1 port map( A1 => n11098, A2 => n11097, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2110 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_200_port, ZN => 
                           n11100);
   U2111 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => 
                           n11120, B2 => 
                           boothmul_pipelined_i_muxes_in_5_199_port, ZN => 
                           n11099);
   U2112 : NAND2_X1 port map( A1 => n11100, A2 => n11099, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2113 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_199_port, ZN => 
                           n11102);
   U2114 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_198_port, ZN => 
                           n11101);
   U2115 : NAND2_X1 port map( A1 => n11102, A2 => n11101, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2116 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_198_port, ZN => 
                           n11104);
   U2117 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_197_port, ZN => 
                           n11103);
   U2118 : NAND2_X1 port map( A1 => n11104, A2 => n11103, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2119 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_197_port, ZN => 
                           n11106);
   U2120 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_196_port, ZN => 
                           n11105);
   U2121 : NAND2_X1 port map( A1 => n11106, A2 => n11105, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2122 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_196_port, ZN => 
                           n11108);
   U2123 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => 
                           n11120, B2 => 
                           boothmul_pipelined_i_muxes_in_5_195_port, ZN => 
                           n11107);
   U2124 : NAND2_X1 port map( A1 => n11108, A2 => n11107, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2125 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_195_port, ZN => 
                           n11110);
   U2126 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_194_port, ZN => 
                           n11109);
   U2127 : NAND2_X1 port map( A1 => n11110, A2 => n11109, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2128 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_194_port, ZN => 
                           n11112);
   U2129 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_193_port, ZN => 
                           n11111);
   U2130 : NAND2_X1 port map( A1 => n11112, A2 => n11111, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2131 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => 
                           n11212, B2 => 
                           boothmul_pipelined_i_muxes_in_5_193_port, ZN => 
                           n11114);
   U2132 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_192_port, ZN => 
                           n11113);
   U2133 : NAND2_X1 port map( A1 => n11114, A2 => n11113, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2134 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => 
                           n11115, B2 => 
                           boothmul_pipelined_i_muxes_in_5_192_port, ZN => 
                           n11118);
   U2135 : AOI22_X1 port map( A1 => n11116, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => 
                           n11120, B2 => 
                           boothmul_pipelined_i_muxes_in_5_191_port, ZN => 
                           n11117);
   U2136 : NAND2_X1 port map( A1 => n11118, A2 => n11117, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2137 : AOI22_X1 port map( A1 => n11119, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => 
                           n11212, B2 => 
                           boothmul_pipelined_i_muxes_in_5_191_port, ZN => 
                           n11122);
   U2138 : NAND2_X1 port map( A1 => n11120, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, ZN => 
                           n11121);
   U2139 : OAI211_X1 port map( C1 => n5128, C2 => n11215, A => n11122, B => 
                           n11121, ZN => boothmul_pipelined_i_mux_out_5_25_port
                           );
   U2140 : NAND3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n11219);
   U2141 : NOR3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n11217);
   U2142 : INV_X1 port map( A => n11217, ZN => n11126);
   U2143 : INV_X1 port map( A => n11124, ZN => n11123);
   U2144 : NAND2_X1 port map( A1 => n3080, A2 => n11123, ZN => n11220);
   U2145 : INV_X1 port map( A => n11220, ZN => n11152);
   U2146 : NOR2_X1 port map( A1 => n3080, A2 => n11124, ZN => n11156);
   U2147 : CLKBUF_X1 port map( A => n11156, Z => n11216);
   U2148 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n11125);
   U2149 : OAI221_X1 port map( B1 => n5123, B2 => n11219, C1 => n5123, C2 => 
                           n11126, A => n11125, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2150 : INV_X1 port map( A => n11219, ZN => n11155);
   U2151 : CLKBUF_X1 port map( A => n11217, Z => n11151);
   U2152 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_6_72_port, A2
                           => n11155, B1 => n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n11128);
   U2153 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => 
                           n11156, B2 => 
                           boothmul_pipelined_i_muxes_in_6_217_port, ZN => 
                           n11127);
   U2154 : NAND2_X1 port map( A1 => n11128, A2 => n11127, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2155 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => 
                           n11217, B2 => 
                           boothmul_pipelined_i_muxes_in_6_217_port, ZN => 
                           n11130);
   U2156 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => 
                           n11156, B2 => 
                           boothmul_pipelined_i_muxes_in_6_216_port, ZN => 
                           n11129);
   U2157 : NAND2_X1 port map( A1 => n11130, A2 => n11129, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2158 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => 
                           n11217, B2 => 
                           boothmul_pipelined_i_muxes_in_6_216_port, ZN => 
                           n11132);
   U2159 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => 
                           n11156, B2 => 
                           boothmul_pipelined_i_muxes_in_6_215_port, ZN => 
                           n11131);
   U2160 : NAND2_X1 port map( A1 => n11132, A2 => n11131, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2161 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_215_port, ZN => 
                           n11134);
   U2162 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_214_port, ZN => 
                           n11133);
   U2163 : NAND2_X1 port map( A1 => n11134, A2 => n11133, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2164 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_214_port, ZN => 
                           n11136);
   U2165 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => 
                           n11156, B2 => 
                           boothmul_pipelined_i_muxes_in_6_213_port, ZN => 
                           n11135);
   U2166 : NAND2_X1 port map( A1 => n11136, A2 => n11135, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2167 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_213_port, ZN => 
                           n11138);
   U2168 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_212_port, ZN => 
                           n11137);
   U2169 : NAND2_X1 port map( A1 => n11138, A2 => n11137, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2170 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_212_port, ZN => 
                           n11140);
   U2171 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_211_port, ZN => 
                           n11139);
   U2172 : NAND2_X1 port map( A1 => n11140, A2 => n11139, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2173 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_211_port, ZN => 
                           n11142);
   U2174 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_210_port, ZN => 
                           n11141);
   U2175 : NAND2_X1 port map( A1 => n11142, A2 => n11141, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2176 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_210_port, ZN => 
                           n11144);
   U2177 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => 
                           n11156, B2 => 
                           boothmul_pipelined_i_muxes_in_6_209_port, ZN => 
                           n11143);
   U2178 : NAND2_X1 port map( A1 => n11144, A2 => n11143, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2179 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_209_port, ZN => 
                           n11146);
   U2180 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_208_port, ZN => 
                           n11145);
   U2181 : NAND2_X1 port map( A1 => n11146, A2 => n11145, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2182 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_208_port, ZN => 
                           n11148);
   U2183 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_207_port, ZN => 
                           n11147);
   U2184 : NAND2_X1 port map( A1 => n11148, A2 => n11147, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2185 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => 
                           n11217, B2 => 
                           boothmul_pipelined_i_muxes_in_6_207_port, ZN => 
                           n11150);
   U2186 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_206_port, ZN => 
                           n11149);
   U2187 : NAND2_X1 port map( A1 => n11150, A2 => n11149, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2188 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => 
                           n11151, B2 => 
                           boothmul_pipelined_i_muxes_in_6_206_port, ZN => 
                           n11154);
   U2189 : AOI22_X1 port map( A1 => n11152, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => 
                           n11156, B2 => 
                           boothmul_pipelined_i_muxes_in_6_205_port, ZN => 
                           n11153);
   U2190 : NAND2_X1 port map( A1 => n11154, A2 => n11153, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2191 : AOI22_X1 port map( A1 => n11155, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => 
                           n11217, B2 => 
                           boothmul_pipelined_i_muxes_in_6_205_port, ZN => 
                           n11158);
   U2192 : NAND2_X1 port map( A1 => n11156, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, ZN => 
                           n11157);
   U2193 : OAI211_X1 port map( C1 => n5129, C2 => n11220, A => n11158, B => 
                           n11157, ZN => boothmul_pipelined_i_mux_out_6_27_port
                           );
   U2194 : NOR2_X1 port map( A1 => n11159, A2 => n11226, ZN => n11176);
   U2195 : INV_X1 port map( A => n11176, ZN => n11163);
   U2196 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           A3 => n7165, ZN => n11199);
   U2197 : INV_X1 port map( A => n11199, ZN => n11162);
   U2198 : NOR2_X1 port map( A1 => n11160, A2 => n11226, ZN => n11193);
   U2199 : CLKBUF_X1 port map( A => n11193, Z => n11197);
   U2200 : NOR2_X1 port map( A1 => n7165, A2 => n11160, ZN => n11177);
   U2201 : CLKBUF_X1 port map( A => n11177, Z => n11198);
   U2202 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_76_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n11161);
   U2203 : OAI221_X1 port map( B1 => n5134, B2 => n11163, C1 => n5134, C2 => 
                           n11162, A => n11161, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2204 : CLKBUF_X1 port map( A => n11199, Z => n11192);
   U2205 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_7_76_port, A2
                           => n11176, B1 => n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n11165);
   U2206 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_231_port, ZN => 
                           n11164);
   U2207 : NAND2_X1 port map( A1 => n11165, A2 => n11164, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2208 : CLKBUF_X1 port map( A => n11176, Z => n11196);
   U2209 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => 
                           n11199, B2 => 
                           boothmul_pipelined_i_muxes_in_7_231_port, ZN => 
                           n11167);
   U2210 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_230_port, ZN => 
                           n11166);
   U2211 : NAND2_X1 port map( A1 => n11167, A2 => n11166, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2212 : AOI22_X1 port map( A1 => n11176, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => 
                           n11199, B2 => 
                           boothmul_pipelined_i_muxes_in_7_230_port, ZN => 
                           n11169);
   U2213 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_229_port, ZN => 
                           n11168);
   U2214 : NAND2_X1 port map( A1 => n11169, A2 => n11168, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2215 : AOI22_X1 port map( A1 => n11176, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_229_port, ZN => 
                           n11171);
   U2216 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_228_port, ZN => 
                           n11170);
   U2217 : NAND2_X1 port map( A1 => n11171, A2 => n11170, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2218 : AOI22_X1 port map( A1 => n11176, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_228_port, ZN => 
                           n11173);
   U2219 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_227_port, ZN => 
                           n11172);
   U2220 : NAND2_X1 port map( A1 => n11173, A2 => n11172, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2221 : AOI22_X1 port map( A1 => n11176, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_227_port, ZN => 
                           n11175);
   U2222 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_226_port, ZN => 
                           n11174);
   U2223 : NAND2_X1 port map( A1 => n11175, A2 => n11174, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2224 : AOI22_X1 port map( A1 => n11176, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_226_port, ZN => 
                           n11179);
   U2225 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => 
                           n11177, B2 => 
                           boothmul_pipelined_i_muxes_in_7_225_port, ZN => 
                           n11178);
   U2226 : NAND2_X1 port map( A1 => n11179, A2 => n11178, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2227 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_225_port, ZN => 
                           n11181);
   U2228 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_224_port, ZN => 
                           n11180);
   U2229 : NAND2_X1 port map( A1 => n11181, A2 => n11180, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2230 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => 
                           n11199, B2 => 
                           boothmul_pipelined_i_muxes_in_7_224_port, ZN => 
                           n11183);
   U2231 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_223_port, ZN => 
                           n11182);
   U2232 : NAND2_X1 port map( A1 => n11183, A2 => n11182, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2233 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_223_port, ZN => 
                           n11185);
   U2234 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_222_port, ZN => 
                           n11184);
   U2235 : NAND2_X1 port map( A1 => n11185, A2 => n11184, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2236 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_222_port, ZN => 
                           n11187);
   U2237 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_221_port, ZN => 
                           n11186);
   U2238 : NAND2_X1 port map( A1 => n11187, A2 => n11186, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2239 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_221_port, ZN => 
                           n11189);
   U2240 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_220_port, ZN => 
                           n11188);
   U2241 : NAND2_X1 port map( A1 => n11189, A2 => n11188, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2242 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => 
                           n11199, B2 => 
                           boothmul_pipelined_i_muxes_in_7_220_port, ZN => 
                           n11191);
   U2243 : AOI22_X1 port map( A1 => n11197, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_219_port, ZN => 
                           n11190);
   U2244 : NAND2_X1 port map( A1 => n11191, A2 => n11190, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2245 : AOI22_X1 port map( A1 => n11196, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => 
                           n11192, B2 => 
                           boothmul_pipelined_i_muxes_in_7_219_port, ZN => 
                           n11195);
   U2246 : AOI22_X1 port map( A1 => n11193, A2 => 
                           boothmul_pipelined_i_muxes_in_7_62_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, ZN => 
                           n11194);
   U2247 : NAND2_X1 port map( A1 => n11195, A2 => n11194, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2248 : OAI21_X1 port map( B1 => n11197, B2 => n11196, A => 
                           boothmul_pipelined_i_muxes_in_7_62_port, ZN => 
                           n11201);
   U2249 : AOI22_X1 port map( A1 => n11199, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n11198, B2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, ZN => 
                           n11200);
   U2250 : NAND2_X1 port map( A1 => n11201, A2 => n11200, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2251 : AOI22_X1 port map( A1 => n11203, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n11202, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n11204);
   U2252 : OAI21_X1 port map( B1 => n11205, B2 => n1993, A => n11204, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2253 : AOI22_X1 port map( A1 => n11207, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, B1 => 
                           n11206, B2 => 
                           boothmul_pipelined_i_muxes_in_4_175_port, ZN => 
                           n11208);
   U2254 : OAI221_X1 port map( B1 => n5127, B2 => n11210, C1 => n5127, C2 => 
                           n11209, A => n11208, ZN => n1997);
   U2255 : AOI22_X1 port map( A1 => n11212, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, B1 => 
                           n11211, B2 => 
                           boothmul_pipelined_i_muxes_in_5_189_port, ZN => 
                           n11213);
   U2256 : OAI221_X1 port map( B1 => n5128, B2 => n11215, C1 => n5128, C2 => 
                           n11214, A => n11213, ZN => n1996);
   U2257 : AOI22_X1 port map( A1 => n11217, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, B1 => 
                           n11216, B2 => 
                           boothmul_pipelined_i_muxes_in_6_203_port, ZN => 
                           n11218);
   U2258 : OAI221_X1 port map( B1 => n5129, B2 => n11220, C1 => n5129, C2 => 
                           n11219, A => n11218, ZN => n1995);
   U2259 : AOI22_X1 port map( A1 => n11222, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, B1 => 
                           n11221, B2 => 
                           boothmul_pipelined_i_muxes_in_3_161_port, ZN => 
                           n11223);
   U2260 : OAI221_X1 port map( B1 => n7164, B2 => n11225, C1 => n7164, C2 => 
                           n11224, A => n11223, ZN => n1991);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, 
      n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, 
      n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, 
      n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, 
      n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, 
      n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, 
      n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, 
      n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, 
      n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, 
      n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, 
      n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, 
      n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, 
      n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, 
      n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, 
      n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, 
      n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, 
      n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, 
      n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, 
      n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, 
      n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, 
      n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, 
      n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, 
      n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, 
      n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, 
      n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, 
      n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, 
      n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, 
      n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, 
      n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, 
      n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, 
      n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, 
      n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, 
      n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, 
      n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, 
      n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, 
      n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, 
      n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, 
      n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, 
      n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, 
      n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, 
      n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, 
      n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, 
      n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, 
      n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, 
      n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, 
      n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, 
      n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, 
      n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, 
      n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, 
      n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, 
      n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, 
      n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, 
      n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, 
      n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, 
      n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, 
      n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, 
      n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, 
      n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, 
      n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, 
      n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, 
      n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, 
      n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, 
      n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, 
      n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, 
      n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, 
      n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, 
      n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, 
      n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, 
      n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, 
      n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, 
      n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, 
      n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, 
      n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, 
      n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, 
      n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, 
      n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, 
      n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, 
      n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, 
      n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, 
      n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, 
      n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, 
      n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, 
      n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, 
      n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, 
      n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, 
      n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, 
      n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, 
      n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, 
      n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, 
      n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, 
      n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, 
      n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, 
      n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, 
      n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, 
      n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, 
      n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, 
      n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, 
      n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, 
      n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, 
      n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, 
      n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, 
      n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, 
      n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, 
      n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, 
      n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, 
      n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, 
      n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, 
      n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, 
      n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, 
      n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, 
      n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, 
      n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, 
      n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, 
      n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, 
      n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, 
      n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, 
      n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, 
      n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, 
      n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, 
      n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, 
      n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, 
      n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, 
      n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, 
      n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, 
      n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, 
      n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, 
      n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, 
      n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, 
      n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, 
      n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, 
      n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, 
      n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, 
      n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, 
      n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, 
      n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, 
      n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, 
      n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, 
      n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, 
      n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, 
      n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, 
      n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, 
      n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, 
      n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, 
      n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, 
      n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, 
      n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, 
      n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, 
      n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, 
      n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, 
      n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, 
      n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, 
      n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, 
      n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, 
      n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, 
      n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, 
      n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, 
      n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, 
      n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, 
      n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, 
      n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, 
      n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, 
      n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, 
      n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, 
      n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, 
      n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, 
      n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, 
      n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, 
      n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, 
      n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, 
      n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, 
      n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, 
      n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, 
      n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, 
      n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, 
      n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, 
      n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, 
      n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, 
      n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, 
      n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, 
      n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, 
      n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, 
      n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, 
      n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, 
      n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, 
      n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, 
      n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, 
      n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, 
      n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, 
      n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, 
      n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, 
      n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, 
      n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, 
      n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, 
      n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, 
      n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, 
      n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, 
      n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, 
      n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, 
      n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, 
      n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, 
      n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, 
      n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, 
      n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, 
      n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, 
      n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, 
      n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, 
      n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, 
      n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, 
      n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, 
      n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, 
      n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, 
      n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, 
      n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, 
      n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, 
      n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, 
      n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, 
      n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, 
      n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, 
      n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, 
      n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, 
      n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, 
      n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, 
      n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, 
      n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, 
      n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, 
      n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, 
      n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, 
      n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, 
      n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, 
      n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, 
      n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, 
      n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, 
      n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, 
      n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, 
      n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, 
      n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, 
      n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, 
      n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, 
      n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, 
      n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, 
      n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, 
      n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, 
      n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, 
      n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, 
      n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, 
      n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, 
      n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, 
      n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, 
      n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, 
      n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, 
      n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, 
      n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, 
      n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, 
      n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, 
      n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, 
      n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, 
      n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, 
      n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, 
      n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, 
      n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, 
      n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, 
      n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, 
      n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, 
      n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, 
      n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, 
      n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, 
      n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, 
      n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, 
      n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, 
      n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, 
      n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, 
      n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, 
      n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, 
      n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, 
      n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, 
      n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, 
      n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, 
      n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, 
      n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, 
      n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, 
      n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, 
      n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, 
      n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, 
      n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, 
      n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, 
      n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, 
      n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, 
      n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, 
      n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, 
      n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, 
      n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, 
      n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, 
      n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, 
      n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, 
      n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, 
      n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, 
      n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, 
      n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, 
      n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, 
      n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, 
      n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, 
      n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, 
      n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, 
      n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, 
      n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, 
      n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, 
      n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, 
      n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, 
      n16775, n16776, n16777, n16778, n16779, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412 : std_logic;

begin
   
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n15763);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n15764);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n15765);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n16034);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n15766);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n16035);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n15767);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n15768);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n15769);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n15770);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n16036);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n16037);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n16038);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n15771);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n16039);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n15772);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n15773);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n16040);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n16041);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n15774);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n16042);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n15775);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n16043);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n15776);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n15777);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n16044);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n15778);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n15779);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n15780);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n16045);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n15781);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n16046);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n16515);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n16276);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n15782);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n15783);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n16277);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n16516);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n16278);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n16279);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n16047);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n16280);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n16517);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n15784);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n16518);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n16281);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n16519);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n16048);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n15785);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n15786);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n15787);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n16282);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n16049);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n15788);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n16050);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n16051);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n15789);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n15790);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n16052);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n16283);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n16053);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n15791);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n16054);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n16284);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n16055);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n15792);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n16285);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n16056);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n16057);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n16058);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n16059);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n15793);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n16286);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n16060);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n15794);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n16061);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n15795);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n16062);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n16063);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n15796);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n16520);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n15797);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n15798);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n16064);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n15799);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n16065);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n15800);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n15801);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n16066);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n15802);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n15803);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n16067);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n16287);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n16521);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n16288);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n16068);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n16289);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n16522);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n16069);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n16070);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n16071);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n15804);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n15805);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n16523);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n16072);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n16073);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n16524);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n16525);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n15806);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n16074);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n16526);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n16527);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n16528);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n16529);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n16530);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n15807);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n15808);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n16531);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n15809);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n16532);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n16533);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n16075);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n16534);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n16076);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n15810);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n16290);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n15811);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n16077);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n15812);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n15813);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n15814);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n16291);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n15815);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n15816);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n16078);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n16079);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n16535);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n15817);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n15818);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n16292);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n16536);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n15819);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n15820);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n16080);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n15821);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n16293);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n16081);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n16294);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n16537);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n16082);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n16538);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n16083);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n15822);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n16295);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n16539);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n16540);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n16296);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n16297);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n16541);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n16298);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n16542);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n16543);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n16544);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n16299);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n16545);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n16300);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n16546);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n16547);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n16548);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n16549);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n15823);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n16301);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n16302);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n16303);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n15824);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n16304);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n16305);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n16550);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n16306);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n16551);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n16307);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n16552);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n16308);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n16553);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n16554);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n16555);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n16084);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n16309);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n16556);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n16085);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n16557);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n16310);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n15825);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n16086);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n16558);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n16559);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n16560);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n16311);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n16312);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n16087);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n15826);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n16313);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n16561);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n15827);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n15828);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n16562);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n16314);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n16563);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n16088);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n16089);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n16315);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n16090);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n16316);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n16317);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n16564);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n16318);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n16319);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n16320);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n16321);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n15829);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n16565);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n16566);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n16322);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n16567);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n16568);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n16569);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n16570);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n16323);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n16324);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n16571);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n16572);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n16325);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n16326);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n16573);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n16327);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n16574);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n16575);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n16576);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n16328);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n16329);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n16577);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n16330);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n16578);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n16579);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n16580);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n16331);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n16332);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n16333);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n16581);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n16582);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n16334);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n16583);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n16091);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n16092);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n16093);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n15830);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n16094);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n16095);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n16096);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n16097);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n16098);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n15831);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n15832);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n16099);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n16100);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n16101);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n15833);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n15834);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n15835);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n16102);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n16103);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n16104);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n15836);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n15837);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n15838);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n15839);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n16105);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n16106);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n16107);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n16108);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n15840);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n16109);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n15841);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n16110);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n15842);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n16111);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n15843);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n15844);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n15845);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n16335);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n16112);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n16336);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n15846);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n16113);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n16114);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n15847);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n15848);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n15849);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n16337);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n15850);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n16115);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n16584);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n16116);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n16585);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n16338);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n15851);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n16117);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n16339);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n15852);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n16118);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n15853);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n16119);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n16120);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n15854);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n16121);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n15855);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n16340);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n15856);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n15857);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n16341);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n16122);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n15858);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n15859);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n16123);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n15860);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n16124);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n15861);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n16586);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n15862);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n16125);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n16126);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n16127);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n15863);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n15864);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n15865);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n15866);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n16128);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n16129);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n16130);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n16131);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n16132);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n15867);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n16133);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n15868);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n16134);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n16587);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n16135);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n16588);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n16589);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n15869);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n16590);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n16136);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n16342);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n16591);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n16343);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n16137);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n16138);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n16592);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n16344);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n15870);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n16593);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n16345);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n16139);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n16594);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n16346);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n16140);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n16347);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n15871);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n16141);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n15872);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n16348);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n16595);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n16596);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n16142);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n16349);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n16597);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n16598);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n16143);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n16599);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n16600);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n16144);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n16350);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n16145);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n16601);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n16602);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n15873);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n15874);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n15875);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n16351);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n16603);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n16604);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n16146);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n16352);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n16605);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n16353);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n16147);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n16148);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n15876);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n15877);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n16149);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n16606);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n16354);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n15878);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n15879);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n16355);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n16356);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n15880);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n16357);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n15881);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n16358);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n15882);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n16150);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n16607);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n16608);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n16359);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n16609);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n16360);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n16361);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n16610);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n16611);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n16612);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n16362);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n16613);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n16363);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n16614);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n15883);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n16364);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n16365);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n16615);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n16616);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n16366);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n16367);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n16617);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n16618);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n16368);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n16151);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n16619);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n16369);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n16370);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n16371);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n16372);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n16620);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n16373);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n15884);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n15885);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n16621);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n16374);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n15886);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n16152);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n16153);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n16622);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n16375);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n16376);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n15887);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n16154);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n16377);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n16155);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n16378);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n16156);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n16379);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n16380);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n16381);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n16623);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n16382);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n15888);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n16624);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n16625);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n16383);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n15889);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n16626);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n16627);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n15890);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n16384);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n15891);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n16628);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n16385);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n16386);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n16387);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n16629);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n16630);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n16388);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n16631);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n16389);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n16390);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n16632);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n16391);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n16392);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n16633);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n16393);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n16634);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n16635);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n16636);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n16637);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n16394);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n16638);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n16639);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n16395);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n16640);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n16641);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n16642);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n16396);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n16397);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n16643);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n16644);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n16645);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n16398);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n16399);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n16400);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n16026);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n15892);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n15893);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n15894);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n16157);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n16158);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n16159);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n16646);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n15895);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n15896);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n16647);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n16160);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n16161);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n16648);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n16162);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n16163);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n16164);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n15897);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n16165);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n16166);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n16167);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n15898);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n16649);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n16168);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n16650);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n15899);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n16169);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n15900);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n16170);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n16171);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n15901);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n15902);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n16027);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n16172);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n15903);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n16651);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n15904);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n15905);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n15906);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n16401);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n16652);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n16653);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n16654);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n16655);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n16173);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n16174);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n16656);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n16402);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n16403);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n15907);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n16175);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n16404);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n16657);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n16405);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n15908);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n15909);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n16176);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n15910);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n15911);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n16658);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n16177);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n16659);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n16406);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n16407);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n15756);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n16178);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n15912);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n16179);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n16180);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n16181);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n15913);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n15914);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n15915);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n15916);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n16182);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n16408);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n15917);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n16183);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n16409);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n16410);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n16184);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n16660);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n16185);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n15918);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n16411);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n16186);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n16661);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n15919);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n15920);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n15921);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n16412);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n15922);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n15923);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n15924);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n16187);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n16188);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n16271);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n16413);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n16662);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n16189);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n16663);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n15925);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n16664);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n16190);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n15926);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n16665);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n16191);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n15927);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n16666);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n15928);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n15929);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n16192);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n15930);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n15931);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n16667);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n16414);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n16415);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n16416);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n16417);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n16193);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n16194);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n16195);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n16196);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n16418);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n16419);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n15932);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n16668);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n15933);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n16028);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n15934);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n16197);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n15935);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n15936);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n15937);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n15938);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n16669);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n16198);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n16420);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n15939);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n15940);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n16199);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n15941);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n15942);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n16670);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n15943);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n16200);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n15944);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n16201);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n15945);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n16202);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n16203);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n16421);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n16204);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n15946);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n15947);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n15948);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n15949);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n15950);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n16205);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n15951);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n15757);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n16206);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n16207);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n15952);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n16208);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n16671);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n16422);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n15953);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n16423);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n15954);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n15955);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n16672);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n15956);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n15957);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n16209);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n15958);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n15959);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n16424);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n16673);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n15960);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n15961);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n15962);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n16210);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n16211);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n16674);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n15963);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n16675);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n16676);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n16212);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n15964);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n16425);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n15965);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n16272);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n15966);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n16426);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n16677);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n16213);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n16427);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n16428);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n15967);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n16678);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n16429);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n16214);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n16215);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n16430);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n16431);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n16432);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n16679);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n16680);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n16681);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n16433);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n16682);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n16216);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n15968);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n16434);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n16683);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n16684);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n16685);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n16435);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n16686);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n16436);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n16437);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n16687);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n16688);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n16273);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n16438);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n16689);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n16439);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n16440);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n16441);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n16690);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n16691);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n16442);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n16692);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n16443);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n16444);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n16693);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n16445);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n16694);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n16446);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n16695);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n16447);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n16448);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n16449);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n16450);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n16696);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n16451);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n16452);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n16453);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n16454);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n16455);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n16697);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n16698);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n16699);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n16700);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n16701);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n16029);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n15969);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n15970);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n15971);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n16217);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n15972);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n16218);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n15973);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n16219);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n16220);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n15974);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n15975);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n16221);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n15976);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n16222);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n15977);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n16223);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n15978);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n15979);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n15980);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n16224);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n15981);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n15982);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n15983);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n15984);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n16456);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n16225);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n16226);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n16702);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n16227);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n15985);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n16228);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n16030);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n16457);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n16703);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n16704);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n16458);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n16229);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n16230);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n16231);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n16232);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n16459);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n16705);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n16233);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n16234);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n16460);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n15986);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n15987);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n16461);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n16235);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n16706);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n15988);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n15989);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n16707);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n16236);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n16462);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n16237);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n16708);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n16238);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n16239);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n16709);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n15990);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n15991);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n16463);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n15758);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n16710);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n16464);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n16711);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n16712);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n16465);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n16466);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n15992);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n16467);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n16240);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n16713);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n16468);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n16469);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n16714);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n16715);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n15993);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n16716);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n16717);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n16241);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n16718);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n16719);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n16720);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n16721);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n16242);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n16470);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n16722);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n16723);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n15994);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n16243);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n16471);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n16244);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n16724);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n15759);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n16725);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n16726);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n16727);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n16472);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n16728);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n16729);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n16730);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n16245);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n16731);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n16473);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n16732);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n16733);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n16246);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n16474);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n16734);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n16475);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n16476);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n16735);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n16736);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n16477);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n16478);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n15995);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n16737);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n15996);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n16479);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n15997);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n16247);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n16480);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n16738);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n16481);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n16739);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n16274);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n16740);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n16482);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n16483);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n16484);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n16741);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n16485);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n16742);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n16743);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n15998);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n16486);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n16744);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n16487);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n16745);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n16746);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n16747);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n15999);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n16748);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n16488);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n16749);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n16750);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n16751);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n16752);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n16753);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n16489);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n16754);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n16755);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n16490);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n16000);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n16756);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n16757);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n16758);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n16031);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n16491);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n16759);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n16492);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n16493);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n16760);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n16001);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n16494);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n16761);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n16762);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n16495);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n16763);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n16496);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n16497);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n16498);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n16764);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n16765);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n16002);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n16499);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n16766);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n16767);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n16500);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n16501);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n16768);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n16502);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n16769);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n16503);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n16770);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n16504);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n16505);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n16506);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n16248);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n15760);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n16249);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n16003);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n16250);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n16251);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n16252);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n16253);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n16004);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n16005);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n16006);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n16254);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n16007);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n16008);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n16255);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n16009);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n16256);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n16010);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n16257);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n16011);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n16012);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n16013);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n16258);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n16014);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n16015);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n16259);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n16260);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n16016);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n16017);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n16018);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n16261);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n16262);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n16019);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n16275);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n16771);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n16263);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n16020);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n16507);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n16508);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n16772);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n16773);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n16509);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n16264);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n16021);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n16022);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n16510);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n16774);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n16265);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n16023);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n16775);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n16776);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n16024);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n16266);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n16267);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n16268);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n16269);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n16511);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n16512);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n16270);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n16777);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n16513);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n16778);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n16779);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n16025);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n16514);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1349);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1350);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1351);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1352);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1353);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1354);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1355);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1356);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1357);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1358);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1359);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1360);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1361);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1362);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1363);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1364);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1365);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1366);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1367);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1368);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1369);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1370);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1371);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1372);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1373);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1374);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1375);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1376);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1377);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1378);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1379);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1380);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1381);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1382);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1383);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1384);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1385);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1386);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1387);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1388);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1389);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1390);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1391);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1392);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1393);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1394);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1395);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1396);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1397);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1398);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1399);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1400);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1401);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1402);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1403);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1404);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1405);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1406);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1407);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1408);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1409);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1410);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1411);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1412);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n16032);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n15761);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n16033);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n15762);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n14003);
   U4 : CLKBUF_X1 port map( A => RESET_BAR, Z => n14004);
   U5 : CLKBUF_X1 port map( A => RESET_BAR, Z => n14005);
   U6 : NAND2_X2 port map( A1 => n14004, A2 => n14180, ZN => n14192);
   U7 : NAND2_X2 port map( A1 => n14003, A2 => n14148, ZN => n14150);
   U8 : NAND2_X2 port map( A1 => n14003, A2 => n14144, ZN => n14146);
   U9 : NAND2_X2 port map( A1 => n14003, A2 => n14140, ZN => n14142);
   U10 : NAND2_X2 port map( A1 => n14003, A2 => n14136, ZN => n14138);
   U11 : NAND2_X2 port map( A1 => n14005, A2 => n14132, ZN => n14134);
   U12 : NAND2_X2 port map( A1 => n14003, A2 => n14128, ZN => n14130);
   U13 : NAND2_X2 port map( A1 => n14003, A2 => n14058, ZN => n14060);
   U14 : NAND2_X2 port map( A1 => n14003, A2 => n14055, ZN => n14057);
   U15 : NAND2_X2 port map( A1 => n14003, A2 => n14052, ZN => n14054);
   U16 : NAND2_X2 port map( A1 => n14003, A2 => n14049, ZN => n14051);
   U17 : NAND2_X2 port map( A1 => n14003, A2 => n14046, ZN => n14048);
   U18 : NAND2_X2 port map( A1 => n14003, A2 => n14043, ZN => n14045);
   U19 : NAND2_X2 port map( A1 => n14003, A2 => n14122, ZN => n14124);
   U20 : NAND2_X2 port map( A1 => n14005, A2 => n14117, ZN => n14119);
   U21 : NAND2_X2 port map( A1 => n14004, A2 => n14114, ZN => n14116);
   U22 : NAND2_X2 port map( A1 => n14004, A2 => n14111, ZN => n14113);
   U23 : NAND2_X2 port map( A1 => n14003, A2 => n14094, ZN => n14106);
   U24 : NAND2_X2 port map( A1 => n14005, A2 => n14070, ZN => n14072);
   U25 : NAND2_X2 port map( A1 => n14004, A2 => n14067, ZN => n14069);
   U26 : NAND2_X2 port map( A1 => n14003, A2 => n14036, ZN => n14038);
   U27 : NAND2_X2 port map( A1 => n14005, A2 => n14030, ZN => n14032);
   U28 : NAND2_X2 port map( A1 => n14003, A2 => n14026, ZN => n14028);
   U29 : INV_X1 port map( A => ADD_WR(4), ZN => n14126);
   U30 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n14029, ZN => n14135);
   U31 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n14066, ZN => n14035);
   U32 : CLKBUF_X1 port map( A => n14973, Z => n14920);
   U33 : CLKBUF_X1 port map( A => n15755, Z => n15700);
   U34 : NAND2_X1 port map( A1 => n14004, A2 => n14152, ZN => n14155);
   U35 : CLKBUF_X1 port map( A => n14122, Z => n14123);
   U36 : NAND2_X1 port map( A1 => n14004, A2 => n14107, ZN => n14110);
   U37 : NAND2_X1 port map( A1 => n14004, A2 => n14062, ZN => n14065);
   U38 : CLKBUF_X1 port map( A => n14089, Z => n14175);
   U39 : CLKBUF_X1 port map( A => n14074, Z => n14160);
   U40 : NAND2_X1 port map( A1 => n14005, A2 => n14039, ZN => n14042);
   U41 : NAND2_X1 port map( A1 => n14005, A2 => n14021, ZN => n14024);
   U42 : NAND2_X1 port map( A1 => n14004, A2 => n14014, ZN => n14017);
   U43 : CLKBUF_X1 port map( A => n14011, Z => n14012);
   U44 : CLKBUF_X1 port map( A => n14008, Z => n14009);
   U45 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n14127);
   U46 : INV_X1 port map( A => ADD_WR(3), ZN => n14006);
   U47 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n14006, ZN => n14066)
                           ;
   U48 : NAND2_X1 port map( A1 => n14127, A2 => n14035, ZN => n14008);
   U49 : NAND2_X1 port map( A1 => n14005, A2 => n14009, ZN => n14010);
   U50 : CLKBUF_X1 port map( A => n14010, Z => n14007);
   U51 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(31), ZN => n14158);
   U52 : CLKBUF_X1 port map( A => n14158, Z => n14121);
   U53 : OAI22_X1 port map( A1 => n16032, A2 => n14007, B1 => n14121, B2 => 
                           n14009, ZN => n2166);
   U54 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(30), ZN => n14073);
   U55 : OAI22_X1 port map( A1 => n15761, A2 => n14010, B1 => n14009, B2 => 
                           n14073, ZN => n2165);
   U56 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(29), ZN => n14074);
   U57 : OAI22_X1 port map( A1 => n16033, A2 => n14007, B1 => n14009, B2 => 
                           n14074, ZN => n2164);
   U58 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(28), ZN => n14075);
   U59 : OAI22_X1 port map( A1 => n15762, A2 => n14010, B1 => n14009, B2 => 
                           n14075, ZN => n2163);
   U60 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(27), ZN => n14076);
   U61 : OAI22_X1 port map( A1 => n15763, A2 => n14007, B1 => n14009, B2 => 
                           n14076, ZN => n2162);
   U62 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(26), ZN => n14077);
   U63 : OAI22_X1 port map( A1 => n15764, A2 => n14010, B1 => n14009, B2 => 
                           n14077, ZN => n2161);
   U64 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(25), ZN => n14078);
   U65 : OAI22_X1 port map( A1 => n15765, A2 => n14007, B1 => n14009, B2 => 
                           n14078, ZN => n2160);
   U66 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(24), ZN => n14079);
   U67 : OAI22_X1 port map( A1 => n16034, A2 => n14010, B1 => n14009, B2 => 
                           n14079, ZN => n2159);
   U68 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(23), ZN => n14080);
   U69 : OAI22_X1 port map( A1 => n15766, A2 => n14007, B1 => n14008, B2 => 
                           n14080, ZN => n2158);
   U70 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(22), ZN => n14081);
   U71 : OAI22_X1 port map( A1 => n16035, A2 => n14010, B1 => n14008, B2 => 
                           n14081, ZN => n2157);
   U72 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(21), ZN => n14082);
   U73 : OAI22_X1 port map( A1 => n15767, A2 => n14010, B1 => n14008, B2 => 
                           n14082, ZN => n2156);
   U74 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(20), ZN => n14083);
   U75 : OAI22_X1 port map( A1 => n15768, A2 => n14010, B1 => n14008, B2 => 
                           n14083, ZN => n2155);
   U76 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(19), ZN => n14084);
   U77 : OAI22_X1 port map( A1 => n15769, A2 => n14007, B1 => n14008, B2 => 
                           n14084, ZN => n2154);
   U78 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(18), ZN => n14085);
   U79 : OAI22_X1 port map( A1 => n15770, A2 => n14007, B1 => n14008, B2 => 
                           n14085, ZN => n2153);
   U80 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(17), ZN => n14086);
   U81 : OAI22_X1 port map( A1 => n16036, A2 => n14007, B1 => n14008, B2 => 
                           n14086, ZN => n2152);
   U82 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(16), ZN => n14087);
   U83 : OAI22_X1 port map( A1 => n16037, A2 => n14007, B1 => n14008, B2 => 
                           n14087, ZN => n2151);
   U84 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(15), ZN => n14088);
   U85 : OAI22_X1 port map( A1 => n16038, A2 => n14007, B1 => n14009, B2 => 
                           n14088, ZN => n2150);
   U86 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(14), ZN => n14089);
   U87 : OAI22_X1 port map( A1 => n15771, A2 => n14007, B1 => n14008, B2 => 
                           n14089, ZN => n2149);
   U88 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(13), ZN => n14090);
   U89 : OAI22_X1 port map( A1 => n16039, A2 => n14007, B1 => n14009, B2 => 
                           n14090, ZN => n2148);
   U90 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(12), ZN => n14091);
   U91 : OAI22_X1 port map( A1 => n15772, A2 => n14007, B1 => n14008, B2 => 
                           n14091, ZN => n2147);
   U92 : NAND2_X1 port map( A1 => RESET_BAR, A2 => DATAIN(11), ZN => n14092);
   U93 : OAI22_X1 port map( A1 => n15773, A2 => n14007, B1 => n14008, B2 => 
                           n14092, ZN => n2146);
   U94 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(10), ZN => n14093);
   U95 : OAI22_X1 port map( A1 => n16040, A2 => n14007, B1 => n14008, B2 => 
                           n14093, ZN => n2145);
   U96 : NAND2_X1 port map( A1 => n14004, A2 => DATAIN(9), ZN => n14095);
   U97 : OAI22_X1 port map( A1 => n16041, A2 => n14007, B1 => n14009, B2 => 
                           n14095, ZN => n2144);
   U98 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(8), ZN => n14096);
   U99 : OAI22_X1 port map( A1 => n15774, A2 => n14007, B1 => n14008, B2 => 
                           n14096, ZN => n2143);
   U100 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(7), ZN => n14097);
   U101 : OAI22_X1 port map( A1 => n16042, A2 => n14010, B1 => n14009, B2 => 
                           n14097, ZN => n2142);
   U102 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(6), ZN => n14098);
   U103 : OAI22_X1 port map( A1 => n15775, A2 => n14010, B1 => n14008, B2 => 
                           n14098, ZN => n2141);
   U104 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(5), ZN => n14099);
   U105 : OAI22_X1 port map( A1 => n16043, A2 => n14010, B1 => n14009, B2 => 
                           n14099, ZN => n2140);
   U106 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(4), ZN => n14100);
   U107 : OAI22_X1 port map( A1 => n15776, A2 => n14010, B1 => n14008, B2 => 
                           n14100, ZN => n2139);
   U108 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(3), ZN => n14101);
   U109 : OAI22_X1 port map( A1 => n15777, A2 => n14010, B1 => n14009, B2 => 
                           n14101, ZN => n2138);
   U110 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(2), ZN => n14102);
   U111 : OAI22_X1 port map( A1 => n16044, A2 => n14010, B1 => n14008, B2 => 
                           n14102, ZN => n2137);
   U112 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(1), ZN => n14103);
   U113 : OAI22_X1 port map( A1 => n15778, A2 => n14010, B1 => n14009, B2 => 
                           n14103, ZN => n2136);
   U114 : NAND2_X1 port map( A1 => n14005, A2 => DATAIN(0), ZN => n14105);
   U115 : OAI22_X1 port map( A1 => n15779, A2 => n14010, B1 => n14009, B2 => 
                           n14105, ZN => n2135);
   U116 : INV_X1 port map( A => ADD_WR(0), ZN => n14025);
   U117 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n14025, ZN 
                           => n14131);
   U118 : NAND2_X1 port map( A1 => n14035, A2 => n14131, ZN => n14011);
   U119 : NAND2_X2 port map( A1 => n14004, A2 => n14011, ZN => n14013);
   U120 : OAI22_X1 port map( A1 => n15780, A2 => n14013, B1 => n14158, B2 => 
                           n14012, ZN => n2134);
   U121 : OAI22_X1 port map( A1 => n16045, A2 => n14013, B1 => n14073, B2 => 
                           n14011, ZN => n2133);
   U122 : OAI22_X1 port map( A1 => n15781, A2 => n14013, B1 => n14074, B2 => 
                           n14012, ZN => n2132);
   U123 : OAI22_X1 port map( A1 => n16046, A2 => n14013, B1 => n14075, B2 => 
                           n14011, ZN => n2131);
   U124 : OAI22_X1 port map( A1 => n16515, A2 => n14013, B1 => n14076, B2 => 
                           n14012, ZN => n2130);
   U125 : OAI22_X1 port map( A1 => n16276, A2 => n14013, B1 => n14077, B2 => 
                           n14011, ZN => n2129);
   U126 : OAI22_X1 port map( A1 => n15782, A2 => n14013, B1 => n14078, B2 => 
                           n14012, ZN => n2128);
   U127 : OAI22_X1 port map( A1 => n15783, A2 => n14013, B1 => n14079, B2 => 
                           n14011, ZN => n2127);
   U128 : OAI22_X1 port map( A1 => n16277, A2 => n14013, B1 => n14080, B2 => 
                           n14012, ZN => n2126);
   U129 : OAI22_X1 port map( A1 => n16516, A2 => n14013, B1 => n14081, B2 => 
                           n14011, ZN => n2125);
   U130 : OAI22_X1 port map( A1 => n16278, A2 => n14013, B1 => n14082, B2 => 
                           n14011, ZN => n2124);
   U131 : OAI22_X1 port map( A1 => n16279, A2 => n14013, B1 => n14083, B2 => 
                           n14012, ZN => n2123);
   U132 : OAI22_X1 port map( A1 => n16047, A2 => n14013, B1 => n14084, B2 => 
                           n14011, ZN => n2122);
   U133 : OAI22_X1 port map( A1 => n16280, A2 => n14013, B1 => n14085, B2 => 
                           n14012, ZN => n2121);
   U134 : OAI22_X1 port map( A1 => n16517, A2 => n14013, B1 => n14086, B2 => 
                           n14011, ZN => n2120);
   U135 : OAI22_X1 port map( A1 => n15784, A2 => n14013, B1 => n14087, B2 => 
                           n14012, ZN => n2119);
   U136 : OAI22_X1 port map( A1 => n16518, A2 => n14013, B1 => n14088, B2 => 
                           n14011, ZN => n2118);
   U137 : OAI22_X1 port map( A1 => n16281, A2 => n14013, B1 => n14089, B2 => 
                           n14011, ZN => n2117);
   U138 : OAI22_X1 port map( A1 => n16519, A2 => n14013, B1 => n14090, B2 => 
                           n14011, ZN => n2116);
   U139 : OAI22_X1 port map( A1 => n16048, A2 => n14013, B1 => n14091, B2 => 
                           n14011, ZN => n2115);
   U140 : OAI22_X1 port map( A1 => n15785, A2 => n14013, B1 => n14092, B2 => 
                           n14011, ZN => n2114);
   U141 : OAI22_X1 port map( A1 => n15786, A2 => n14013, B1 => n14093, B2 => 
                           n14011, ZN => n2113);
   U142 : OAI22_X1 port map( A1 => n15787, A2 => n14013, B1 => n14095, B2 => 
                           n14011, ZN => n2112);
   U143 : OAI22_X1 port map( A1 => n16282, A2 => n14013, B1 => n14096, B2 => 
                           n14012, ZN => n2111);
   U144 : OAI22_X1 port map( A1 => n16049, A2 => n14013, B1 => n14097, B2 => 
                           n14012, ZN => n2110);
   U145 : OAI22_X1 port map( A1 => n15788, A2 => n14013, B1 => n14098, B2 => 
                           n14012, ZN => n2109);
   U146 : OAI22_X1 port map( A1 => n16050, A2 => n14013, B1 => n14099, B2 => 
                           n14012, ZN => n2108);
   U147 : OAI22_X1 port map( A1 => n16051, A2 => n14013, B1 => n14100, B2 => 
                           n14012, ZN => n2107);
   U148 : OAI22_X1 port map( A1 => n15789, A2 => n14013, B1 => n14101, B2 => 
                           n14012, ZN => n2106);
   U149 : OAI22_X1 port map( A1 => n15790, A2 => n14013, B1 => n14102, B2 => 
                           n14012, ZN => n2105);
   U150 : OAI22_X1 port map( A1 => n16052, A2 => n14013, B1 => n14103, B2 => 
                           n14012, ZN => n2104);
   U151 : OAI22_X1 port map( A1 => n16283, A2 => n14013, B1 => n14105, B2 => 
                           n14012, ZN => n2103);
   U152 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n14025, ZN => n14029);
   U153 : NAND2_X1 port map( A1 => n14035, A2 => n14135, ZN => n14014);
   U154 : CLKBUF_X1 port map( A => n14017, Z => n14015);
   U155 : CLKBUF_X1 port map( A => n14014, Z => n14016);
   U156 : OAI22_X1 port map( A1 => n16053, A2 => n14015, B1 => n14121, B2 => 
                           n14016, ZN => n2102);
   U157 : OAI22_X1 port map( A1 => n15791, A2 => n14017, B1 => n14073, B2 => 
                           n14014, ZN => n2101);
   U158 : OAI22_X1 port map( A1 => n16054, A2 => n14015, B1 => n14074, B2 => 
                           n14016, ZN => n2100);
   U159 : OAI22_X1 port map( A1 => n16284, A2 => n14017, B1 => n14075, B2 => 
                           n14014, ZN => n2099);
   U160 : OAI22_X1 port map( A1 => n16055, A2 => n14015, B1 => n14076, B2 => 
                           n14016, ZN => n2098);
   U161 : OAI22_X1 port map( A1 => n15792, A2 => n14017, B1 => n14077, B2 => 
                           n14014, ZN => n2097);
   U162 : OAI22_X1 port map( A1 => n16285, A2 => n14015, B1 => n14078, B2 => 
                           n14016, ZN => n2096);
   U163 : OAI22_X1 port map( A1 => n16056, A2 => n14017, B1 => n14079, B2 => 
                           n14014, ZN => n2095);
   U164 : OAI22_X1 port map( A1 => n16057, A2 => n14015, B1 => n14080, B2 => 
                           n14016, ZN => n2094);
   U165 : OAI22_X1 port map( A1 => n16058, A2 => n14017, B1 => n14081, B2 => 
                           n14014, ZN => n2093);
   U166 : OAI22_X1 port map( A1 => n16059, A2 => n14017, B1 => n14082, B2 => 
                           n14014, ZN => n2092);
   U167 : OAI22_X1 port map( A1 => n15793, A2 => n14017, B1 => n14083, B2 => 
                           n14016, ZN => n2091);
   U168 : OAI22_X1 port map( A1 => n16286, A2 => n14015, B1 => n14084, B2 => 
                           n14014, ZN => n2090);
   U169 : OAI22_X1 port map( A1 => n16060, A2 => n14015, B1 => n14085, B2 => 
                           n14016, ZN => n2089);
   U170 : OAI22_X1 port map( A1 => n15794, A2 => n14015, B1 => n14086, B2 => 
                           n14014, ZN => n2088);
   U171 : OAI22_X1 port map( A1 => n16061, A2 => n14015, B1 => n14087, B2 => 
                           n14016, ZN => n2087);
   U172 : OAI22_X1 port map( A1 => n15795, A2 => n14015, B1 => n14088, B2 => 
                           n14014, ZN => n2086);
   U173 : OAI22_X1 port map( A1 => n16062, A2 => n14015, B1 => n14089, B2 => 
                           n14014, ZN => n2085);
   U174 : OAI22_X1 port map( A1 => n16063, A2 => n14015, B1 => n14090, B2 => 
                           n14014, ZN => n2084);
   U175 : OAI22_X1 port map( A1 => n15796, A2 => n14015, B1 => n14091, B2 => 
                           n14014, ZN => n2083);
   U176 : OAI22_X1 port map( A1 => n16520, A2 => n14015, B1 => n14092, B2 => 
                           n14014, ZN => n2082);
   U177 : OAI22_X1 port map( A1 => n15797, A2 => n14015, B1 => n14093, B2 => 
                           n14014, ZN => n2081);
   U178 : OAI22_X1 port map( A1 => n15798, A2 => n14015, B1 => n14095, B2 => 
                           n14014, ZN => n2080);
   U179 : OAI22_X1 port map( A1 => n16064, A2 => n14015, B1 => n14096, B2 => 
                           n14016, ZN => n2079);
   U180 : OAI22_X1 port map( A1 => n15799, A2 => n14017, B1 => n14097, B2 => 
                           n14016, ZN => n2078);
   U181 : OAI22_X1 port map( A1 => n16065, A2 => n14017, B1 => n14098, B2 => 
                           n14016, ZN => n2077);
   U182 : OAI22_X1 port map( A1 => n15800, A2 => n14017, B1 => n14099, B2 => 
                           n14016, ZN => n2076);
   U183 : OAI22_X1 port map( A1 => n15801, A2 => n14017, B1 => n14100, B2 => 
                           n14016, ZN => n2075);
   U184 : OAI22_X1 port map( A1 => n16066, A2 => n14017, B1 => n14101, B2 => 
                           n14016, ZN => n2074);
   U185 : OAI22_X1 port map( A1 => n15802, A2 => n14017, B1 => n14102, B2 => 
                           n14016, ZN => n2073);
   U186 : OAI22_X1 port map( A1 => n15803, A2 => n14017, B1 => n14103, B2 => 
                           n14016, ZN => n2072);
   U187 : OAI22_X1 port map( A1 => n16067, A2 => n14017, B1 => n14105, B2 => 
                           n14016, ZN => n2071);
   U188 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n14033);
   U189 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n14033, ZN => n14139);
   U190 : NAND2_X1 port map( A1 => n14035, A2 => n14139, ZN => n14018);
   U191 : NAND2_X2 port map( A1 => n14003, A2 => n14018, ZN => n14020);
   U192 : CLKBUF_X1 port map( A => n14018, Z => n14019);
   U193 : OAI22_X1 port map( A1 => n16287, A2 => n14020, B1 => n14158, B2 => 
                           n14019, ZN => n2070);
   U194 : OAI22_X1 port map( A1 => n16521, A2 => n14020, B1 => n14073, B2 => 
                           n14018, ZN => n2069);
   U195 : OAI22_X1 port map( A1 => n16288, A2 => n14020, B1 => n14074, B2 => 
                           n14019, ZN => n2068);
   U196 : OAI22_X1 port map( A1 => n16068, A2 => n14020, B1 => n14075, B2 => 
                           n14018, ZN => n2067);
   U197 : OAI22_X1 port map( A1 => n16289, A2 => n14020, B1 => n14076, B2 => 
                           n14019, ZN => n2066);
   U198 : OAI22_X1 port map( A1 => n16522, A2 => n14020, B1 => n14077, B2 => 
                           n14018, ZN => n2065);
   U199 : OAI22_X1 port map( A1 => n16069, A2 => n14020, B1 => n14078, B2 => 
                           n14019, ZN => n2064);
   U200 : OAI22_X1 port map( A1 => n16070, A2 => n14020, B1 => n14079, B2 => 
                           n14018, ZN => n2063);
   U201 : OAI22_X1 port map( A1 => n16071, A2 => n14020, B1 => n14080, B2 => 
                           n14019, ZN => n2062);
   U202 : OAI22_X1 port map( A1 => n15804, A2 => n14020, B1 => n14081, B2 => 
                           n14018, ZN => n2061);
   U203 : OAI22_X1 port map( A1 => n15805, A2 => n14020, B1 => n14082, B2 => 
                           n14018, ZN => n2060);
   U204 : OAI22_X1 port map( A1 => n16523, A2 => n14020, B1 => n14083, B2 => 
                           n14019, ZN => n2059);
   U205 : OAI22_X1 port map( A1 => n16072, A2 => n14020, B1 => n14084, B2 => 
                           n14018, ZN => n2058);
   U206 : OAI22_X1 port map( A1 => n16073, A2 => n14020, B1 => n14085, B2 => 
                           n14019, ZN => n2057);
   U207 : OAI22_X1 port map( A1 => n16524, A2 => n14020, B1 => n14086, B2 => 
                           n14018, ZN => n2056);
   U208 : OAI22_X1 port map( A1 => n16525, A2 => n14020, B1 => n14087, B2 => 
                           n14019, ZN => n2055);
   U209 : OAI22_X1 port map( A1 => n15806, A2 => n14020, B1 => n14088, B2 => 
                           n14018, ZN => n2054);
   U210 : OAI22_X1 port map( A1 => n16074, A2 => n14020, B1 => n14089, B2 => 
                           n14018, ZN => n2053);
   U211 : OAI22_X1 port map( A1 => n16526, A2 => n14020, B1 => n14090, B2 => 
                           n14018, ZN => n2052);
   U212 : OAI22_X1 port map( A1 => n16527, A2 => n14020, B1 => n14091, B2 => 
                           n14018, ZN => n2051);
   U213 : OAI22_X1 port map( A1 => n16528, A2 => n14020, B1 => n14092, B2 => 
                           n14018, ZN => n2050);
   U214 : OAI22_X1 port map( A1 => n16529, A2 => n14020, B1 => n14093, B2 => 
                           n14018, ZN => n2049);
   U215 : OAI22_X1 port map( A1 => n16530, A2 => n14020, B1 => n14095, B2 => 
                           n14018, ZN => n2048);
   U216 : OAI22_X1 port map( A1 => n15807, A2 => n14020, B1 => n14096, B2 => 
                           n14019, ZN => n2047);
   U217 : OAI22_X1 port map( A1 => n15808, A2 => n14020, B1 => n14097, B2 => 
                           n14019, ZN => n2046);
   U218 : OAI22_X1 port map( A1 => n16531, A2 => n14020, B1 => n14098, B2 => 
                           n14019, ZN => n2045);
   U219 : OAI22_X1 port map( A1 => n15809, A2 => n14020, B1 => n14099, B2 => 
                           n14019, ZN => n2044);
   U220 : OAI22_X1 port map( A1 => n16532, A2 => n14020, B1 => n14100, B2 => 
                           n14019, ZN => n2043);
   U221 : OAI22_X1 port map( A1 => n16533, A2 => n14020, B1 => n14101, B2 => 
                           n14019, ZN => n2042);
   U222 : OAI22_X1 port map( A1 => n16075, A2 => n14020, B1 => n14102, B2 => 
                           n14019, ZN => n2041);
   U223 : OAI22_X1 port map( A1 => n16534, A2 => n14020, B1 => n14103, B2 => 
                           n14019, ZN => n2040);
   U224 : OAI22_X1 port map( A1 => n16076, A2 => n14020, B1 => n14105, B2 => 
                           n14019, ZN => n2039);
   U225 : INV_X1 port map( A => ADD_WR(2), ZN => n14034);
   U226 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n14034, ZN 
                           => n14143);
   U227 : NAND2_X1 port map( A1 => n14035, A2 => n14143, ZN => n14021);
   U228 : CLKBUF_X1 port map( A => n14024, Z => n14022);
   U229 : CLKBUF_X1 port map( A => n14021, Z => n14023);
   U230 : OAI22_X1 port map( A1 => n15810, A2 => n14022, B1 => n14121, B2 => 
                           n14023, ZN => n2038);
   U231 : OAI22_X1 port map( A1 => n16290, A2 => n14024, B1 => n14073, B2 => 
                           n14021, ZN => n2037);
   U232 : OAI22_X1 port map( A1 => n15811, A2 => n14022, B1 => n14074, B2 => 
                           n14023, ZN => n2036);
   U233 : OAI22_X1 port map( A1 => n16077, A2 => n14024, B1 => n14075, B2 => 
                           n14021, ZN => n2035);
   U234 : OAI22_X1 port map( A1 => n15812, A2 => n14022, B1 => n14076, B2 => 
                           n14023, ZN => n2034);
   U235 : OAI22_X1 port map( A1 => n15813, A2 => n14024, B1 => n14077, B2 => 
                           n14021, ZN => n2033);
   U236 : OAI22_X1 port map( A1 => n15814, A2 => n14022, B1 => n14078, B2 => 
                           n14023, ZN => n2032);
   U237 : OAI22_X1 port map( A1 => n16291, A2 => n14024, B1 => n14079, B2 => 
                           n14021, ZN => n2031);
   U238 : OAI22_X1 port map( A1 => n15815, A2 => n14022, B1 => n14080, B2 => 
                           n14023, ZN => n2030);
   U239 : OAI22_X1 port map( A1 => n15816, A2 => n14024, B1 => n14081, B2 => 
                           n14021, ZN => n2029);
   U240 : OAI22_X1 port map( A1 => n16078, A2 => n14024, B1 => n14082, B2 => 
                           n14021, ZN => n2028);
   U241 : OAI22_X1 port map( A1 => n16079, A2 => n14024, B1 => n14083, B2 => 
                           n14023, ZN => n2027);
   U242 : OAI22_X1 port map( A1 => n16535, A2 => n14022, B1 => n14084, B2 => 
                           n14021, ZN => n2026);
   U243 : OAI22_X1 port map( A1 => n15817, A2 => n14022, B1 => n14085, B2 => 
                           n14023, ZN => n2025);
   U244 : OAI22_X1 port map( A1 => n15818, A2 => n14022, B1 => n14086, B2 => 
                           n14021, ZN => n2024);
   U245 : OAI22_X1 port map( A1 => n16292, A2 => n14022, B1 => n14087, B2 => 
                           n14023, ZN => n2023);
   U246 : OAI22_X1 port map( A1 => n16536, A2 => n14022, B1 => n14088, B2 => 
                           n14021, ZN => n2022);
   U247 : OAI22_X1 port map( A1 => n15819, A2 => n14022, B1 => n14089, B2 => 
                           n14021, ZN => n2021);
   U248 : OAI22_X1 port map( A1 => n15820, A2 => n14022, B1 => n14090, B2 => 
                           n14021, ZN => n2020);
   U249 : OAI22_X1 port map( A1 => n16080, A2 => n14022, B1 => n14091, B2 => 
                           n14021, ZN => n2019);
   U250 : OAI22_X1 port map( A1 => n15821, A2 => n14022, B1 => n14092, B2 => 
                           n14021, ZN => n2018);
   U251 : OAI22_X1 port map( A1 => n16293, A2 => n14022, B1 => n14093, B2 => 
                           n14021, ZN => n2017);
   U252 : OAI22_X1 port map( A1 => n16081, A2 => n14022, B1 => n14095, B2 => 
                           n14021, ZN => n2016);
   U253 : OAI22_X1 port map( A1 => n16294, A2 => n14022, B1 => n14096, B2 => 
                           n14023, ZN => n2015);
   U254 : OAI22_X1 port map( A1 => n16537, A2 => n14024, B1 => n14097, B2 => 
                           n14023, ZN => n2014);
   U255 : OAI22_X1 port map( A1 => n16082, A2 => n14024, B1 => n14098, B2 => 
                           n14023, ZN => n2013);
   U256 : OAI22_X1 port map( A1 => n16538, A2 => n14024, B1 => n14099, B2 => 
                           n14023, ZN => n2012);
   U257 : OAI22_X1 port map( A1 => n16083, A2 => n14024, B1 => n14100, B2 => 
                           n14023, ZN => n2011);
   U258 : OAI22_X1 port map( A1 => n15822, A2 => n14024, B1 => n14101, B2 => 
                           n14023, ZN => n2010);
   U259 : OAI22_X1 port map( A1 => n16295, A2 => n14024, B1 => n14102, B2 => 
                           n14023, ZN => n2009);
   U260 : OAI22_X1 port map( A1 => n16539, A2 => n14024, B1 => n14103, B2 => 
                           n14023, ZN => n2008);
   U261 : OAI22_X1 port map( A1 => n16540, A2 => n14024, B1 => n14105, B2 => 
                           n14023, ZN => n2007);
   U262 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n14025, A3 => n14034, ZN => 
                           n14147);
   U263 : NAND2_X1 port map( A1 => n14035, A2 => n14147, ZN => n14026);
   U264 : CLKBUF_X1 port map( A => n14026, Z => n14027);
   U265 : OAI22_X1 port map( A1 => n16296, A2 => n14028, B1 => n14158, B2 => 
                           n14027, ZN => n2006);
   U266 : OAI22_X1 port map( A1 => n16297, A2 => n14028, B1 => n14073, B2 => 
                           n14026, ZN => n2005);
   U267 : OAI22_X1 port map( A1 => n16541, A2 => n14028, B1 => n14074, B2 => 
                           n14027, ZN => n2004);
   U268 : OAI22_X1 port map( A1 => n16298, A2 => n14028, B1 => n14075, B2 => 
                           n14026, ZN => n2003);
   U269 : OAI22_X1 port map( A1 => n16542, A2 => n14028, B1 => n14076, B2 => 
                           n14027, ZN => n2002);
   U270 : OAI22_X1 port map( A1 => n16543, A2 => n14028, B1 => n14077, B2 => 
                           n14026, ZN => n2001);
   U271 : OAI22_X1 port map( A1 => n16544, A2 => n14028, B1 => n14078, B2 => 
                           n14027, ZN => n2000);
   U272 : OAI22_X1 port map( A1 => n16299, A2 => n14028, B1 => n14079, B2 => 
                           n14026, ZN => n1999);
   U273 : OAI22_X1 port map( A1 => n16545, A2 => n14028, B1 => n14080, B2 => 
                           n14027, ZN => n1998);
   U274 : OAI22_X1 port map( A1 => n16300, A2 => n14028, B1 => n14081, B2 => 
                           n14026, ZN => n1997);
   U275 : OAI22_X1 port map( A1 => n16546, A2 => n14028, B1 => n14082, B2 => 
                           n14026, ZN => n1996);
   U276 : OAI22_X1 port map( A1 => n16547, A2 => n14028, B1 => n14083, B2 => 
                           n14027, ZN => n1995);
   U277 : OAI22_X1 port map( A1 => n16548, A2 => n14028, B1 => n14084, B2 => 
                           n14026, ZN => n1994);
   U278 : OAI22_X1 port map( A1 => n16549, A2 => n14028, B1 => n14085, B2 => 
                           n14027, ZN => n1993);
   U279 : OAI22_X1 port map( A1 => n15823, A2 => n14028, B1 => n14086, B2 => 
                           n14026, ZN => n1992);
   U280 : OAI22_X1 port map( A1 => n16301, A2 => n14028, B1 => n14087, B2 => 
                           n14027, ZN => n1991);
   U281 : OAI22_X1 port map( A1 => n16302, A2 => n14028, B1 => n14088, B2 => 
                           n14026, ZN => n1990);
   U282 : OAI22_X1 port map( A1 => n16303, A2 => n14028, B1 => n14089, B2 => 
                           n14026, ZN => n1989);
   U283 : OAI22_X1 port map( A1 => n15824, A2 => n14028, B1 => n14090, B2 => 
                           n14026, ZN => n1988);
   U284 : OAI22_X1 port map( A1 => n16304, A2 => n14028, B1 => n14091, B2 => 
                           n14026, ZN => n1987);
   U285 : OAI22_X1 port map( A1 => n16305, A2 => n14028, B1 => n14092, B2 => 
                           n14026, ZN => n1986);
   U286 : OAI22_X1 port map( A1 => n16550, A2 => n14028, B1 => n14093, B2 => 
                           n14026, ZN => n1985);
   U287 : OAI22_X1 port map( A1 => n16306, A2 => n14028, B1 => n14095, B2 => 
                           n14026, ZN => n1984);
   U288 : OAI22_X1 port map( A1 => n16551, A2 => n14028, B1 => n14096, B2 => 
                           n14027, ZN => n1983);
   U289 : OAI22_X1 port map( A1 => n16307, A2 => n14028, B1 => n14097, B2 => 
                           n14027, ZN => n1982);
   U290 : OAI22_X1 port map( A1 => n16552, A2 => n14028, B1 => n14098, B2 => 
                           n14027, ZN => n1981);
   U291 : OAI22_X1 port map( A1 => n16308, A2 => n14028, B1 => n14099, B2 => 
                           n14027, ZN => n1980);
   U292 : OAI22_X1 port map( A1 => n16553, A2 => n14028, B1 => n14100, B2 => 
                           n14027, ZN => n1979);
   U293 : OAI22_X1 port map( A1 => n16554, A2 => n14028, B1 => n14101, B2 => 
                           n14027, ZN => n1978);
   U294 : OAI22_X1 port map( A1 => n16555, A2 => n14028, B1 => n14102, B2 => 
                           n14027, ZN => n1977);
   U295 : OAI22_X1 port map( A1 => n16084, A2 => n14028, B1 => n14103, B2 => 
                           n14027, ZN => n1976);
   U296 : OAI22_X1 port map( A1 => n16309, A2 => n14028, B1 => n14105, B2 => 
                           n14027, ZN => n1975);
   U297 : NOR2_X1 port map( A1 => n14034, A2 => n14029, ZN => n14151);
   U298 : NAND2_X1 port map( A1 => n14035, A2 => n14151, ZN => n14030);
   U299 : CLKBUF_X1 port map( A => n14030, Z => n14031);
   U300 : OAI22_X1 port map( A1 => n16556, A2 => n14032, B1 => n14121, B2 => 
                           n14031, ZN => n1974);
   U301 : OAI22_X1 port map( A1 => n16085, A2 => n14032, B1 => n14073, B2 => 
                           n14030, ZN => n1973);
   U302 : OAI22_X1 port map( A1 => n16557, A2 => n14032, B1 => n14074, B2 => 
                           n14031, ZN => n1972);
   U303 : OAI22_X1 port map( A1 => n16310, A2 => n14032, B1 => n14075, B2 => 
                           n14030, ZN => n1971);
   U304 : OAI22_X1 port map( A1 => n15825, A2 => n14032, B1 => n14076, B2 => 
                           n14031, ZN => n1970);
   U305 : OAI22_X1 port map( A1 => n16086, A2 => n14032, B1 => n14077, B2 => 
                           n14030, ZN => n1969);
   U306 : OAI22_X1 port map( A1 => n16558, A2 => n14032, B1 => n14078, B2 => 
                           n14031, ZN => n1968);
   U307 : OAI22_X1 port map( A1 => n16559, A2 => n14032, B1 => n14079, B2 => 
                           n14030, ZN => n1967);
   U308 : OAI22_X1 port map( A1 => n16560, A2 => n14032, B1 => n14080, B2 => 
                           n14031, ZN => n1966);
   U309 : OAI22_X1 port map( A1 => n16311, A2 => n14032, B1 => n14081, B2 => 
                           n14030, ZN => n1965);
   U310 : OAI22_X1 port map( A1 => n16312, A2 => n14032, B1 => n14082, B2 => 
                           n14030, ZN => n1964);
   U311 : OAI22_X1 port map( A1 => n16087, A2 => n14032, B1 => n14083, B2 => 
                           n14031, ZN => n1963);
   U312 : OAI22_X1 port map( A1 => n15826, A2 => n14032, B1 => n14084, B2 => 
                           n14030, ZN => n1962);
   U313 : OAI22_X1 port map( A1 => n16313, A2 => n14032, B1 => n14085, B2 => 
                           n14031, ZN => n1961);
   U314 : OAI22_X1 port map( A1 => n16561, A2 => n14032, B1 => n14086, B2 => 
                           n14030, ZN => n1960);
   U315 : OAI22_X1 port map( A1 => n15827, A2 => n14032, B1 => n14087, B2 => 
                           n14031, ZN => n1959);
   U316 : OAI22_X1 port map( A1 => n15828, A2 => n14032, B1 => n14088, B2 => 
                           n14030, ZN => n1958);
   U317 : OAI22_X1 port map( A1 => n16562, A2 => n14032, B1 => n14089, B2 => 
                           n14030, ZN => n1957);
   U318 : OAI22_X1 port map( A1 => n16314, A2 => n14032, B1 => n14090, B2 => 
                           n14030, ZN => n1956);
   U319 : OAI22_X1 port map( A1 => n16563, A2 => n14032, B1 => n14091, B2 => 
                           n14030, ZN => n1955);
   U320 : OAI22_X1 port map( A1 => n16088, A2 => n14032, B1 => n14092, B2 => 
                           n14030, ZN => n1954);
   U321 : OAI22_X1 port map( A1 => n16089, A2 => n14032, B1 => n14093, B2 => 
                           n14030, ZN => n1953);
   U322 : OAI22_X1 port map( A1 => n16315, A2 => n14032, B1 => n14095, B2 => 
                           n14030, ZN => n1952);
   U323 : OAI22_X1 port map( A1 => n16090, A2 => n14032, B1 => n14096, B2 => 
                           n14031, ZN => n1951);
   U324 : OAI22_X1 port map( A1 => n16316, A2 => n14032, B1 => n14097, B2 => 
                           n14031, ZN => n1950);
   U325 : OAI22_X1 port map( A1 => n16317, A2 => n14032, B1 => n14098, B2 => 
                           n14031, ZN => n1949);
   U326 : OAI22_X1 port map( A1 => n16564, A2 => n14032, B1 => n14099, B2 => 
                           n14031, ZN => n1948);
   U327 : OAI22_X1 port map( A1 => n16318, A2 => n14032, B1 => n14100, B2 => 
                           n14031, ZN => n1947);
   U328 : OAI22_X1 port map( A1 => n16319, A2 => n14032, B1 => n14101, B2 => 
                           n14031, ZN => n1946);
   U329 : OAI22_X1 port map( A1 => n16320, A2 => n14032, B1 => n14102, B2 => 
                           n14031, ZN => n1945);
   U330 : OAI22_X1 port map( A1 => n16321, A2 => n14032, B1 => n14103, B2 => 
                           n14031, ZN => n1944);
   U331 : OAI22_X1 port map( A1 => n15829, A2 => n14032, B1 => n14105, B2 => 
                           n14031, ZN => n1943);
   U332 : NOR2_X1 port map( A1 => n14034, A2 => n14033, ZN => n14157);
   U333 : NAND2_X1 port map( A1 => n14035, A2 => n14157, ZN => n14036);
   U334 : CLKBUF_X1 port map( A => n14036, Z => n14037);
   U335 : OAI22_X1 port map( A1 => n16565, A2 => n14038, B1 => n14158, B2 => 
                           n14037, ZN => n1942);
   U336 : OAI22_X1 port map( A1 => n16566, A2 => n14038, B1 => n14073, B2 => 
                           n14036, ZN => n1941);
   U337 : OAI22_X1 port map( A1 => n16322, A2 => n14038, B1 => n14074, B2 => 
                           n14037, ZN => n1940);
   U338 : OAI22_X1 port map( A1 => n16567, A2 => n14038, B1 => n14075, B2 => 
                           n14036, ZN => n1939);
   U339 : OAI22_X1 port map( A1 => n16568, A2 => n14038, B1 => n14076, B2 => 
                           n14037, ZN => n1938);
   U340 : OAI22_X1 port map( A1 => n16569, A2 => n14038, B1 => n14077, B2 => 
                           n14036, ZN => n1937);
   U341 : OAI22_X1 port map( A1 => n16570, A2 => n14038, B1 => n14078, B2 => 
                           n14037, ZN => n1936);
   U342 : OAI22_X1 port map( A1 => n16323, A2 => n14038, B1 => n14079, B2 => 
                           n14036, ZN => n1935);
   U343 : OAI22_X1 port map( A1 => n16324, A2 => n14038, B1 => n14080, B2 => 
                           n14037, ZN => n1934);
   U344 : OAI22_X1 port map( A1 => n16571, A2 => n14038, B1 => n14081, B2 => 
                           n14036, ZN => n1933);
   U345 : OAI22_X1 port map( A1 => n16572, A2 => n14038, B1 => n14082, B2 => 
                           n14036, ZN => n1932);
   U346 : OAI22_X1 port map( A1 => n16325, A2 => n14038, B1 => n14083, B2 => 
                           n14037, ZN => n1931);
   U347 : OAI22_X1 port map( A1 => n16326, A2 => n14038, B1 => n14084, B2 => 
                           n14036, ZN => n1930);
   U348 : OAI22_X1 port map( A1 => n16573, A2 => n14038, B1 => n14085, B2 => 
                           n14037, ZN => n1929);
   U349 : OAI22_X1 port map( A1 => n16327, A2 => n14038, B1 => n14086, B2 => 
                           n14036, ZN => n1928);
   U350 : OAI22_X1 port map( A1 => n16574, A2 => n14038, B1 => n14087, B2 => 
                           n14037, ZN => n1927);
   U351 : OAI22_X1 port map( A1 => n16575, A2 => n14038, B1 => n14088, B2 => 
                           n14036, ZN => n1926);
   U352 : OAI22_X1 port map( A1 => n16576, A2 => n14038, B1 => n14089, B2 => 
                           n14036, ZN => n1925);
   U353 : OAI22_X1 port map( A1 => n16328, A2 => n14038, B1 => n14090, B2 => 
                           n14036, ZN => n1924);
   U354 : OAI22_X1 port map( A1 => n16329, A2 => n14038, B1 => n14091, B2 => 
                           n14036, ZN => n1923);
   U355 : OAI22_X1 port map( A1 => n16577, A2 => n14038, B1 => n14092, B2 => 
                           n14036, ZN => n1922);
   U356 : OAI22_X1 port map( A1 => n16330, A2 => n14038, B1 => n14093, B2 => 
                           n14036, ZN => n1921);
   U357 : OAI22_X1 port map( A1 => n16578, A2 => n14038, B1 => n14095, B2 => 
                           n14036, ZN => n1920);
   U358 : OAI22_X1 port map( A1 => n16579, A2 => n14038, B1 => n14096, B2 => 
                           n14037, ZN => n1919);
   U359 : OAI22_X1 port map( A1 => n16580, A2 => n14038, B1 => n14097, B2 => 
                           n14037, ZN => n1918);
   U360 : OAI22_X1 port map( A1 => n16331, A2 => n14038, B1 => n14098, B2 => 
                           n14037, ZN => n1917);
   U361 : OAI22_X1 port map( A1 => n16332, A2 => n14038, B1 => n14099, B2 => 
                           n14037, ZN => n1916);
   U362 : OAI22_X1 port map( A1 => n16333, A2 => n14038, B1 => n14100, B2 => 
                           n14037, ZN => n1915);
   U363 : OAI22_X1 port map( A1 => n16581, A2 => n14038, B1 => n14101, B2 => 
                           n14037, ZN => n1914);
   U364 : OAI22_X1 port map( A1 => n16582, A2 => n14038, B1 => n14102, B2 => 
                           n14037, ZN => n1913);
   U365 : OAI22_X1 port map( A1 => n16334, A2 => n14038, B1 => n14103, B2 => 
                           n14037, ZN => n1912);
   U366 : OAI22_X1 port map( A1 => n16583, A2 => n14038, B1 => n14105, B2 => 
                           n14037, ZN => n1911);
   U367 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(3), ZN => 
                           n14125);
   U368 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n14125, ZN => n14061);
   U369 : NAND2_X1 port map( A1 => n14127, A2 => n14061, ZN => n14039);
   U370 : CLKBUF_X1 port map( A => n14042, Z => n14040);
   U371 : CLKBUF_X1 port map( A => n14039, Z => n14041);
   U372 : OAI22_X1 port map( A1 => n16091, A2 => n14040, B1 => n14121, B2 => 
                           n14041, ZN => n1910);
   U373 : OAI22_X1 port map( A1 => n16092, A2 => n14042, B1 => n14073, B2 => 
                           n14039, ZN => n1909);
   U374 : OAI22_X1 port map( A1 => n16093, A2 => n14040, B1 => n14074, B2 => 
                           n14041, ZN => n1908);
   U375 : OAI22_X1 port map( A1 => n15830, A2 => n14042, B1 => n14075, B2 => 
                           n14039, ZN => n1907);
   U376 : OAI22_X1 port map( A1 => n16094, A2 => n14040, B1 => n14076, B2 => 
                           n14041, ZN => n1906);
   U377 : OAI22_X1 port map( A1 => n16095, A2 => n14042, B1 => n14077, B2 => 
                           n14039, ZN => n1905);
   U378 : OAI22_X1 port map( A1 => n16096, A2 => n14040, B1 => n14078, B2 => 
                           n14041, ZN => n1904);
   U379 : OAI22_X1 port map( A1 => n16097, A2 => n14042, B1 => n14079, B2 => 
                           n14039, ZN => n1903);
   U380 : OAI22_X1 port map( A1 => n16098, A2 => n14040, B1 => n14080, B2 => 
                           n14041, ZN => n1902);
   U381 : OAI22_X1 port map( A1 => n15831, A2 => n14042, B1 => n14081, B2 => 
                           n14039, ZN => n1901);
   U382 : OAI22_X1 port map( A1 => n15832, A2 => n14042, B1 => n14082, B2 => 
                           n14039, ZN => n1900);
   U383 : OAI22_X1 port map( A1 => n16099, A2 => n14042, B1 => n14083, B2 => 
                           n14041, ZN => n1899);
   U384 : OAI22_X1 port map( A1 => n16100, A2 => n14040, B1 => n14084, B2 => 
                           n14039, ZN => n1898);
   U385 : OAI22_X1 port map( A1 => n16101, A2 => n14040, B1 => n14085, B2 => 
                           n14041, ZN => n1897);
   U386 : OAI22_X1 port map( A1 => n15833, A2 => n14040, B1 => n14086, B2 => 
                           n14039, ZN => n1896);
   U387 : OAI22_X1 port map( A1 => n15834, A2 => n14040, B1 => n14087, B2 => 
                           n14041, ZN => n1895);
   U388 : OAI22_X1 port map( A1 => n15835, A2 => n14040, B1 => n14088, B2 => 
                           n14039, ZN => n1894);
   U389 : OAI22_X1 port map( A1 => n16102, A2 => n14040, B1 => n14089, B2 => 
                           n14039, ZN => n1893);
   U390 : OAI22_X1 port map( A1 => n16103, A2 => n14040, B1 => n14090, B2 => 
                           n14039, ZN => n1892);
   U391 : OAI22_X1 port map( A1 => n16104, A2 => n14040, B1 => n14091, B2 => 
                           n14039, ZN => n1891);
   U392 : OAI22_X1 port map( A1 => n15836, A2 => n14040, B1 => n14092, B2 => 
                           n14039, ZN => n1890);
   U393 : OAI22_X1 port map( A1 => n15837, A2 => n14040, B1 => n14093, B2 => 
                           n14039, ZN => n1889);
   U394 : OAI22_X1 port map( A1 => n15838, A2 => n14040, B1 => n14095, B2 => 
                           n14039, ZN => n1888);
   U395 : OAI22_X1 port map( A1 => n15839, A2 => n14040, B1 => n14096, B2 => 
                           n14041, ZN => n1887);
   U396 : OAI22_X1 port map( A1 => n16105, A2 => n14042, B1 => n14097, B2 => 
                           n14041, ZN => n1886);
   U397 : OAI22_X1 port map( A1 => n16106, A2 => n14042, B1 => n14098, B2 => 
                           n14041, ZN => n1885);
   U398 : OAI22_X1 port map( A1 => n16107, A2 => n14042, B1 => n14099, B2 => 
                           n14041, ZN => n1884);
   U399 : OAI22_X1 port map( A1 => n16108, A2 => n14042, B1 => n14100, B2 => 
                           n14041, ZN => n1883);
   U400 : OAI22_X1 port map( A1 => n15840, A2 => n14042, B1 => n14101, B2 => 
                           n14041, ZN => n1882);
   U401 : OAI22_X1 port map( A1 => n16109, A2 => n14042, B1 => n14102, B2 => 
                           n14041, ZN => n1881);
   U402 : OAI22_X1 port map( A1 => n15841, A2 => n14042, B1 => n14103, B2 => 
                           n14041, ZN => n1880);
   U403 : OAI22_X1 port map( A1 => n16110, A2 => n14042, B1 => n14105, B2 => 
                           n14041, ZN => n1879);
   U404 : NAND2_X1 port map( A1 => n14131, A2 => n14061, ZN => n14043);
   U405 : CLKBUF_X1 port map( A => n14043, Z => n14044);
   U406 : OAI22_X1 port map( A1 => n15842, A2 => n14045, B1 => n14158, B2 => 
                           n14044, ZN => n1878);
   U407 : OAI22_X1 port map( A1 => n16111, A2 => n14045, B1 => n14073, B2 => 
                           n14043, ZN => n1877);
   U408 : OAI22_X1 port map( A1 => n15843, A2 => n14045, B1 => n14074, B2 => 
                           n14044, ZN => n1876);
   U409 : OAI22_X1 port map( A1 => n15844, A2 => n14045, B1 => n14075, B2 => 
                           n14043, ZN => n1875);
   U410 : OAI22_X1 port map( A1 => n15845, A2 => n14045, B1 => n14076, B2 => 
                           n14044, ZN => n1874);
   U411 : OAI22_X1 port map( A1 => n16335, A2 => n14045, B1 => n14077, B2 => 
                           n14043, ZN => n1873);
   U412 : OAI22_X1 port map( A1 => n16112, A2 => n14045, B1 => n14078, B2 => 
                           n14044, ZN => n1872);
   U413 : OAI22_X1 port map( A1 => n16336, A2 => n14045, B1 => n14079, B2 => 
                           n14043, ZN => n1871);
   U414 : OAI22_X1 port map( A1 => n15846, A2 => n14045, B1 => n14080, B2 => 
                           n14044, ZN => n1870);
   U415 : OAI22_X1 port map( A1 => n16113, A2 => n14045, B1 => n14081, B2 => 
                           n14043, ZN => n1869);
   U416 : OAI22_X1 port map( A1 => n16114, A2 => n14045, B1 => n14082, B2 => 
                           n14043, ZN => n1868);
   U417 : OAI22_X1 port map( A1 => n15847, A2 => n14045, B1 => n14083, B2 => 
                           n14044, ZN => n1867);
   U418 : OAI22_X1 port map( A1 => n15848, A2 => n14045, B1 => n14084, B2 => 
                           n14043, ZN => n1866);
   U419 : OAI22_X1 port map( A1 => n15849, A2 => n14045, B1 => n14085, B2 => 
                           n14044, ZN => n1865);
   U420 : OAI22_X1 port map( A1 => n16337, A2 => n14045, B1 => n14086, B2 => 
                           n14043, ZN => n1864);
   U421 : OAI22_X1 port map( A1 => n15850, A2 => n14045, B1 => n14087, B2 => 
                           n14044, ZN => n1863);
   U422 : OAI22_X1 port map( A1 => n16115, A2 => n14045, B1 => n14088, B2 => 
                           n14043, ZN => n1862);
   U423 : OAI22_X1 port map( A1 => n16584, A2 => n14045, B1 => n14089, B2 => 
                           n14043, ZN => n1861);
   U424 : OAI22_X1 port map( A1 => n16116, A2 => n14045, B1 => n14090, B2 => 
                           n14043, ZN => n1860);
   U425 : OAI22_X1 port map( A1 => n16585, A2 => n14045, B1 => n14091, B2 => 
                           n14043, ZN => n1859);
   U426 : OAI22_X1 port map( A1 => n16338, A2 => n14045, B1 => n14092, B2 => 
                           n14043, ZN => n1858);
   U427 : OAI22_X1 port map( A1 => n15851, A2 => n14045, B1 => n14093, B2 => 
                           n14043, ZN => n1857);
   U428 : OAI22_X1 port map( A1 => n16117, A2 => n14045, B1 => n14095, B2 => 
                           n14043, ZN => n1856);
   U429 : OAI22_X1 port map( A1 => n16339, A2 => n14045, B1 => n14096, B2 => 
                           n14044, ZN => n1855);
   U430 : OAI22_X1 port map( A1 => n15852, A2 => n14045, B1 => n14097, B2 => 
                           n14044, ZN => n1854);
   U431 : OAI22_X1 port map( A1 => n16118, A2 => n14045, B1 => n14098, B2 => 
                           n14044, ZN => n1853);
   U432 : OAI22_X1 port map( A1 => n15853, A2 => n14045, B1 => n14099, B2 => 
                           n14044, ZN => n1852);
   U433 : OAI22_X1 port map( A1 => n16119, A2 => n14045, B1 => n14100, B2 => 
                           n14044, ZN => n1851);
   U434 : OAI22_X1 port map( A1 => n16120, A2 => n14045, B1 => n14101, B2 => 
                           n14044, ZN => n1850);
   U435 : OAI22_X1 port map( A1 => n15854, A2 => n14045, B1 => n14102, B2 => 
                           n14044, ZN => n1849);
   U436 : OAI22_X1 port map( A1 => n16121, A2 => n14045, B1 => n14103, B2 => 
                           n14044, ZN => n1848);
   U437 : OAI22_X1 port map( A1 => n15855, A2 => n14045, B1 => n14105, B2 => 
                           n14044, ZN => n1847);
   U438 : NAND2_X1 port map( A1 => n14135, A2 => n14061, ZN => n14046);
   U439 : CLKBUF_X1 port map( A => n14046, Z => n14047);
   U440 : OAI22_X1 port map( A1 => n16340, A2 => n14048, B1 => n14158, B2 => 
                           n14047, ZN => n1846);
   U441 : OAI22_X1 port map( A1 => n15856, A2 => n14048, B1 => n14073, B2 => 
                           n14046, ZN => n1845);
   U442 : OAI22_X1 port map( A1 => n15857, A2 => n14048, B1 => n14074, B2 => 
                           n14047, ZN => n1844);
   U443 : OAI22_X1 port map( A1 => n16341, A2 => n14048, B1 => n14075, B2 => 
                           n14046, ZN => n1843);
   U444 : OAI22_X1 port map( A1 => n16122, A2 => n14048, B1 => n14076, B2 => 
                           n14047, ZN => n1842);
   U445 : OAI22_X1 port map( A1 => n15858, A2 => n14048, B1 => n14077, B2 => 
                           n14046, ZN => n1841);
   U446 : OAI22_X1 port map( A1 => n15859, A2 => n14048, B1 => n14078, B2 => 
                           n14047, ZN => n1840);
   U447 : OAI22_X1 port map( A1 => n16123, A2 => n14048, B1 => n14079, B2 => 
                           n14046, ZN => n1839);
   U448 : OAI22_X1 port map( A1 => n15860, A2 => n14048, B1 => n14080, B2 => 
                           n14047, ZN => n1838);
   U449 : OAI22_X1 port map( A1 => n16124, A2 => n14048, B1 => n14081, B2 => 
                           n14046, ZN => n1837);
   U450 : OAI22_X1 port map( A1 => n15861, A2 => n14048, B1 => n14082, B2 => 
                           n14046, ZN => n1836);
   U451 : OAI22_X1 port map( A1 => n16586, A2 => n14048, B1 => n14083, B2 => 
                           n14047, ZN => n1835);
   U452 : OAI22_X1 port map( A1 => n15862, A2 => n14048, B1 => n14084, B2 => 
                           n14046, ZN => n1834);
   U453 : OAI22_X1 port map( A1 => n16125, A2 => n14048, B1 => n14085, B2 => 
                           n14047, ZN => n1833);
   U454 : OAI22_X1 port map( A1 => n16126, A2 => n14048, B1 => n14086, B2 => 
                           n14046, ZN => n1832);
   U455 : OAI22_X1 port map( A1 => n16127, A2 => n14048, B1 => n14087, B2 => 
                           n14047, ZN => n1831);
   U456 : OAI22_X1 port map( A1 => n15863, A2 => n14048, B1 => n14088, B2 => 
                           n14046, ZN => n1830);
   U457 : OAI22_X1 port map( A1 => n15864, A2 => n14048, B1 => n14089, B2 => 
                           n14046, ZN => n1829);
   U458 : OAI22_X1 port map( A1 => n15865, A2 => n14048, B1 => n14090, B2 => 
                           n14046, ZN => n1828);
   U459 : OAI22_X1 port map( A1 => n15866, A2 => n14048, B1 => n14091, B2 => 
                           n14046, ZN => n1827);
   U460 : OAI22_X1 port map( A1 => n16128, A2 => n14048, B1 => n14092, B2 => 
                           n14046, ZN => n1826);
   U461 : OAI22_X1 port map( A1 => n16129, A2 => n14048, B1 => n14093, B2 => 
                           n14046, ZN => n1825);
   U462 : OAI22_X1 port map( A1 => n16130, A2 => n14048, B1 => n14095, B2 => 
                           n14046, ZN => n1824);
   U463 : OAI22_X1 port map( A1 => n16131, A2 => n14048, B1 => n14096, B2 => 
                           n14047, ZN => n1823);
   U464 : OAI22_X1 port map( A1 => n16132, A2 => n14048, B1 => n14097, B2 => 
                           n14047, ZN => n1822);
   U465 : OAI22_X1 port map( A1 => n15867, A2 => n14048, B1 => n14098, B2 => 
                           n14047, ZN => n1821);
   U466 : OAI22_X1 port map( A1 => n16133, A2 => n14048, B1 => n14099, B2 => 
                           n14047, ZN => n1820);
   U467 : OAI22_X1 port map( A1 => n15868, A2 => n14048, B1 => n14100, B2 => 
                           n14047, ZN => n1819);
   U468 : OAI22_X1 port map( A1 => n16134, A2 => n14048, B1 => n14101, B2 => 
                           n14047, ZN => n1818);
   U469 : OAI22_X1 port map( A1 => n16587, A2 => n14048, B1 => n14102, B2 => 
                           n14047, ZN => n1817);
   U470 : OAI22_X1 port map( A1 => n16135, A2 => n14048, B1 => n14103, B2 => 
                           n14047, ZN => n1816);
   U471 : OAI22_X1 port map( A1 => n16588, A2 => n14048, B1 => n14105, B2 => 
                           n14047, ZN => n1815);
   U472 : NAND2_X1 port map( A1 => n14139, A2 => n14061, ZN => n14049);
   U473 : CLKBUF_X1 port map( A => n14049, Z => n14050);
   U474 : OAI22_X1 port map( A1 => n16589, A2 => n14051, B1 => n14158, B2 => 
                           n14050, ZN => n1814);
   U475 : CLKBUF_X1 port map( A => n14073, Z => n14159);
   U476 : OAI22_X1 port map( A1 => n15869, A2 => n14051, B1 => n14159, B2 => 
                           n14049, ZN => n1813);
   U477 : OAI22_X1 port map( A1 => n16590, A2 => n14051, B1 => n14160, B2 => 
                           n14050, ZN => n1812);
   U478 : CLKBUF_X1 port map( A => n14075, Z => n14161);
   U479 : OAI22_X1 port map( A1 => n16136, A2 => n14051, B1 => n14161, B2 => 
                           n14049, ZN => n1811);
   U480 : CLKBUF_X1 port map( A => n14076, Z => n14162);
   U481 : OAI22_X1 port map( A1 => n16342, A2 => n14051, B1 => n14162, B2 => 
                           n14050, ZN => n1810);
   U482 : CLKBUF_X1 port map( A => n14077, Z => n14163);
   U483 : OAI22_X1 port map( A1 => n16591, A2 => n14051, B1 => n14163, B2 => 
                           n14049, ZN => n1809);
   U484 : CLKBUF_X1 port map( A => n14078, Z => n14164);
   U485 : OAI22_X1 port map( A1 => n16343, A2 => n14051, B1 => n14164, B2 => 
                           n14050, ZN => n1808);
   U486 : CLKBUF_X1 port map( A => n14079, Z => n14165);
   U487 : OAI22_X1 port map( A1 => n16137, A2 => n14051, B1 => n14165, B2 => 
                           n14049, ZN => n1807);
   U488 : CLKBUF_X1 port map( A => n14080, Z => n14166);
   U489 : OAI22_X1 port map( A1 => n16138, A2 => n14051, B1 => n14166, B2 => 
                           n14050, ZN => n1806);
   U490 : CLKBUF_X1 port map( A => n14081, Z => n14167);
   U491 : OAI22_X1 port map( A1 => n16592, A2 => n14051, B1 => n14167, B2 => 
                           n14049, ZN => n1805);
   U492 : CLKBUF_X1 port map( A => n14082, Z => n14168);
   U493 : OAI22_X1 port map( A1 => n16344, A2 => n14051, B1 => n14168, B2 => 
                           n14049, ZN => n1804);
   U494 : CLKBUF_X1 port map( A => n14083, Z => n14169);
   U495 : OAI22_X1 port map( A1 => n15870, A2 => n14051, B1 => n14169, B2 => 
                           n14050, ZN => n1803);
   U496 : CLKBUF_X1 port map( A => n14084, Z => n14170);
   U497 : OAI22_X1 port map( A1 => n16593, A2 => n14051, B1 => n14170, B2 => 
                           n14049, ZN => n1802);
   U498 : CLKBUF_X1 port map( A => n14085, Z => n14171);
   U499 : OAI22_X1 port map( A1 => n16345, A2 => n14051, B1 => n14171, B2 => 
                           n14050, ZN => n1801);
   U500 : CLKBUF_X1 port map( A => n14086, Z => n14172);
   U501 : OAI22_X1 port map( A1 => n16139, A2 => n14051, B1 => n14172, B2 => 
                           n14049, ZN => n1800);
   U502 : CLKBUF_X1 port map( A => n14087, Z => n14173);
   U503 : OAI22_X1 port map( A1 => n16594, A2 => n14051, B1 => n14173, B2 => 
                           n14050, ZN => n1799);
   U504 : CLKBUF_X1 port map( A => n14088, Z => n14174);
   U505 : OAI22_X1 port map( A1 => n16346, A2 => n14051, B1 => n14174, B2 => 
                           n14049, ZN => n1798);
   U506 : OAI22_X1 port map( A1 => n16140, A2 => n14051, B1 => n14175, B2 => 
                           n14049, ZN => n1797);
   U507 : CLKBUF_X1 port map( A => n14090, Z => n14176);
   U508 : OAI22_X1 port map( A1 => n16347, A2 => n14051, B1 => n14176, B2 => 
                           n14049, ZN => n1796);
   U509 : CLKBUF_X1 port map( A => n14091, Z => n14177);
   U510 : OAI22_X1 port map( A1 => n15871, A2 => n14051, B1 => n14177, B2 => 
                           n14049, ZN => n1795);
   U511 : CLKBUF_X1 port map( A => n14092, Z => n14178);
   U512 : OAI22_X1 port map( A1 => n16141, A2 => n14051, B1 => n14178, B2 => 
                           n14049, ZN => n1794);
   U513 : CLKBUF_X1 port map( A => n14093, Z => n14179);
   U514 : OAI22_X1 port map( A1 => n15872, A2 => n14051, B1 => n14179, B2 => 
                           n14049, ZN => n1793);
   U515 : CLKBUF_X1 port map( A => n14095, Z => n14181);
   U516 : OAI22_X1 port map( A1 => n16348, A2 => n14051, B1 => n14181, B2 => 
                           n14049, ZN => n1792);
   U517 : CLKBUF_X1 port map( A => n14096, Z => n14182);
   U518 : OAI22_X1 port map( A1 => n16595, A2 => n14051, B1 => n14182, B2 => 
                           n14050, ZN => n1791);
   U519 : CLKBUF_X1 port map( A => n14097, Z => n14183);
   U520 : OAI22_X1 port map( A1 => n16596, A2 => n14051, B1 => n14183, B2 => 
                           n14050, ZN => n1790);
   U521 : CLKBUF_X1 port map( A => n14098, Z => n14184);
   U522 : OAI22_X1 port map( A1 => n16142, A2 => n14051, B1 => n14184, B2 => 
                           n14050, ZN => n1789);
   U523 : CLKBUF_X1 port map( A => n14099, Z => n14185);
   U524 : OAI22_X1 port map( A1 => n16349, A2 => n14051, B1 => n14185, B2 => 
                           n14050, ZN => n1788);
   U525 : CLKBUF_X1 port map( A => n14100, Z => n14186);
   U526 : OAI22_X1 port map( A1 => n16597, A2 => n14051, B1 => n14186, B2 => 
                           n14050, ZN => n1787);
   U527 : CLKBUF_X1 port map( A => n14101, Z => n14187);
   U528 : OAI22_X1 port map( A1 => n16598, A2 => n14051, B1 => n14187, B2 => 
                           n14050, ZN => n1786);
   U529 : CLKBUF_X1 port map( A => n14102, Z => n14188);
   U530 : OAI22_X1 port map( A1 => n16143, A2 => n14051, B1 => n14188, B2 => 
                           n14050, ZN => n1785);
   U531 : CLKBUF_X1 port map( A => n14103, Z => n14189);
   U532 : OAI22_X1 port map( A1 => n16599, A2 => n14051, B1 => n14189, B2 => 
                           n14050, ZN => n1784);
   U533 : CLKBUF_X1 port map( A => n14105, Z => n14191);
   U534 : OAI22_X1 port map( A1 => n16600, A2 => n14051, B1 => n14191, B2 => 
                           n14050, ZN => n1783);
   U535 : NAND2_X1 port map( A1 => n14143, A2 => n14061, ZN => n14052);
   U536 : CLKBUF_X1 port map( A => n14052, Z => n14053);
   U537 : OAI22_X1 port map( A1 => n16144, A2 => n14054, B1 => n14121, B2 => 
                           n14053, ZN => n1782);
   U538 : OAI22_X1 port map( A1 => n16350, A2 => n14054, B1 => n14073, B2 => 
                           n14052, ZN => n1781);
   U539 : OAI22_X1 port map( A1 => n16145, A2 => n14054, B1 => n14074, B2 => 
                           n14053, ZN => n1780);
   U540 : OAI22_X1 port map( A1 => n16601, A2 => n14054, B1 => n14075, B2 => 
                           n14052, ZN => n1779);
   U541 : OAI22_X1 port map( A1 => n16602, A2 => n14054, B1 => n14076, B2 => 
                           n14053, ZN => n1778);
   U542 : OAI22_X1 port map( A1 => n15873, A2 => n14054, B1 => n14077, B2 => 
                           n14052, ZN => n1777);
   U543 : OAI22_X1 port map( A1 => n15874, A2 => n14054, B1 => n14078, B2 => 
                           n14053, ZN => n1776);
   U544 : OAI22_X1 port map( A1 => n15875, A2 => n14054, B1 => n14079, B2 => 
                           n14052, ZN => n1775);
   U545 : OAI22_X1 port map( A1 => n16351, A2 => n14054, B1 => n14080, B2 => 
                           n14053, ZN => n1774);
   U546 : OAI22_X1 port map( A1 => n16603, A2 => n14054, B1 => n14081, B2 => 
                           n14052, ZN => n1773);
   U547 : OAI22_X1 port map( A1 => n16604, A2 => n14054, B1 => n14082, B2 => 
                           n14052, ZN => n1772);
   U548 : OAI22_X1 port map( A1 => n16146, A2 => n14054, B1 => n14083, B2 => 
                           n14053, ZN => n1771);
   U549 : OAI22_X1 port map( A1 => n16352, A2 => n14054, B1 => n14084, B2 => 
                           n14052, ZN => n1770);
   U550 : OAI22_X1 port map( A1 => n16605, A2 => n14054, B1 => n14085, B2 => 
                           n14053, ZN => n1769);
   U551 : OAI22_X1 port map( A1 => n16353, A2 => n14054, B1 => n14086, B2 => 
                           n14052, ZN => n1768);
   U552 : OAI22_X1 port map( A1 => n16147, A2 => n14054, B1 => n14087, B2 => 
                           n14053, ZN => n1767);
   U553 : OAI22_X1 port map( A1 => n16148, A2 => n14054, B1 => n14088, B2 => 
                           n14052, ZN => n1766);
   U554 : OAI22_X1 port map( A1 => n15876, A2 => n14054, B1 => n14089, B2 => 
                           n14052, ZN => n1765);
   U555 : OAI22_X1 port map( A1 => n15877, A2 => n14054, B1 => n14090, B2 => 
                           n14052, ZN => n1764);
   U556 : OAI22_X1 port map( A1 => n16149, A2 => n14054, B1 => n14091, B2 => 
                           n14052, ZN => n1763);
   U557 : OAI22_X1 port map( A1 => n16606, A2 => n14054, B1 => n14092, B2 => 
                           n14052, ZN => n1762);
   U558 : OAI22_X1 port map( A1 => n16354, A2 => n14054, B1 => n14093, B2 => 
                           n14052, ZN => n1761);
   U559 : OAI22_X1 port map( A1 => n15878, A2 => n14054, B1 => n14095, B2 => 
                           n14052, ZN => n1760);
   U560 : OAI22_X1 port map( A1 => n15879, A2 => n14054, B1 => n14096, B2 => 
                           n14053, ZN => n1759);
   U561 : OAI22_X1 port map( A1 => n16355, A2 => n14054, B1 => n14097, B2 => 
                           n14053, ZN => n1758);
   U562 : OAI22_X1 port map( A1 => n16356, A2 => n14054, B1 => n14098, B2 => 
                           n14053, ZN => n1757);
   U563 : OAI22_X1 port map( A1 => n15880, A2 => n14054, B1 => n14099, B2 => 
                           n14053, ZN => n1756);
   U564 : OAI22_X1 port map( A1 => n16357, A2 => n14054, B1 => n14100, B2 => 
                           n14053, ZN => n1755);
   U565 : OAI22_X1 port map( A1 => n15881, A2 => n14054, B1 => n14101, B2 => 
                           n14053, ZN => n1754);
   U566 : OAI22_X1 port map( A1 => n16358, A2 => n14054, B1 => n14102, B2 => 
                           n14053, ZN => n1753);
   U567 : OAI22_X1 port map( A1 => n15882, A2 => n14054, B1 => n14103, B2 => 
                           n14053, ZN => n1752);
   U568 : OAI22_X1 port map( A1 => n16150, A2 => n14054, B1 => n14105, B2 => 
                           n14053, ZN => n1751);
   U569 : NAND2_X1 port map( A1 => n14147, A2 => n14061, ZN => n14055);
   U570 : CLKBUF_X1 port map( A => n14055, Z => n14056);
   U571 : OAI22_X1 port map( A1 => n16607, A2 => n14057, B1 => n14121, B2 => 
                           n14056, ZN => n1750);
   U572 : OAI22_X1 port map( A1 => n16608, A2 => n14057, B1 => n14159, B2 => 
                           n14055, ZN => n1749);
   U573 : OAI22_X1 port map( A1 => n16359, A2 => n14057, B1 => n14160, B2 => 
                           n14056, ZN => n1748);
   U574 : OAI22_X1 port map( A1 => n16609, A2 => n14057, B1 => n14161, B2 => 
                           n14055, ZN => n1747);
   U575 : OAI22_X1 port map( A1 => n16360, A2 => n14057, B1 => n14162, B2 => 
                           n14056, ZN => n1746);
   U576 : OAI22_X1 port map( A1 => n16361, A2 => n14057, B1 => n14163, B2 => 
                           n14055, ZN => n1745);
   U577 : OAI22_X1 port map( A1 => n16610, A2 => n14057, B1 => n14164, B2 => 
                           n14056, ZN => n1744);
   U578 : OAI22_X1 port map( A1 => n16611, A2 => n14057, B1 => n14165, B2 => 
                           n14055, ZN => n1743);
   U579 : OAI22_X1 port map( A1 => n16612, A2 => n14057, B1 => n14166, B2 => 
                           n14056, ZN => n1742);
   U580 : OAI22_X1 port map( A1 => n16362, A2 => n14057, B1 => n14167, B2 => 
                           n14055, ZN => n1741);
   U581 : OAI22_X1 port map( A1 => n16613, A2 => n14057, B1 => n14168, B2 => 
                           n14055, ZN => n1740);
   U582 : OAI22_X1 port map( A1 => n16363, A2 => n14057, B1 => n14169, B2 => 
                           n14056, ZN => n1739);
   U583 : OAI22_X1 port map( A1 => n16614, A2 => n14057, B1 => n14170, B2 => 
                           n14055, ZN => n1738);
   U584 : OAI22_X1 port map( A1 => n15883, A2 => n14057, B1 => n14171, B2 => 
                           n14056, ZN => n1737);
   U585 : OAI22_X1 port map( A1 => n16364, A2 => n14057, B1 => n14172, B2 => 
                           n14055, ZN => n1736);
   U586 : OAI22_X1 port map( A1 => n16365, A2 => n14057, B1 => n14173, B2 => 
                           n14056, ZN => n1735);
   U587 : OAI22_X1 port map( A1 => n16615, A2 => n14057, B1 => n14174, B2 => 
                           n14055, ZN => n1734);
   U588 : OAI22_X1 port map( A1 => n16616, A2 => n14057, B1 => n14175, B2 => 
                           n14055, ZN => n1733);
   U589 : OAI22_X1 port map( A1 => n16366, A2 => n14057, B1 => n14176, B2 => 
                           n14055, ZN => n1732);
   U590 : OAI22_X1 port map( A1 => n16367, A2 => n14057, B1 => n14177, B2 => 
                           n14055, ZN => n1731);
   U591 : OAI22_X1 port map( A1 => n16617, A2 => n14057, B1 => n14178, B2 => 
                           n14055, ZN => n1730);
   U592 : OAI22_X1 port map( A1 => n16618, A2 => n14057, B1 => n14179, B2 => 
                           n14055, ZN => n1729);
   U593 : OAI22_X1 port map( A1 => n16368, A2 => n14057, B1 => n14181, B2 => 
                           n14055, ZN => n1728);
   U594 : OAI22_X1 port map( A1 => n16151, A2 => n14057, B1 => n14182, B2 => 
                           n14056, ZN => n1727);
   U595 : OAI22_X1 port map( A1 => n16619, A2 => n14057, B1 => n14183, B2 => 
                           n14056, ZN => n1726);
   U596 : OAI22_X1 port map( A1 => n16369, A2 => n14057, B1 => n14184, B2 => 
                           n14056, ZN => n1725);
   U597 : OAI22_X1 port map( A1 => n16370, A2 => n14057, B1 => n14185, B2 => 
                           n14056, ZN => n1724);
   U598 : OAI22_X1 port map( A1 => n16371, A2 => n14057, B1 => n14186, B2 => 
                           n14056, ZN => n1723);
   U599 : OAI22_X1 port map( A1 => n16372, A2 => n14057, B1 => n14187, B2 => 
                           n14056, ZN => n1722);
   U600 : OAI22_X1 port map( A1 => n16620, A2 => n14057, B1 => n14188, B2 => 
                           n14056, ZN => n1721);
   U601 : OAI22_X1 port map( A1 => n16373, A2 => n14057, B1 => n14189, B2 => 
                           n14056, ZN => n1720);
   U602 : OAI22_X1 port map( A1 => n15884, A2 => n14057, B1 => n14191, B2 => 
                           n14056, ZN => n1719);
   U603 : NAND2_X1 port map( A1 => n14151, A2 => n14061, ZN => n14058);
   U604 : CLKBUF_X1 port map( A => n14058, Z => n14059);
   U605 : OAI22_X1 port map( A1 => n15885, A2 => n14060, B1 => n14121, B2 => 
                           n14059, ZN => n1718);
   U606 : OAI22_X1 port map( A1 => n16621, A2 => n14060, B1 => n14073, B2 => 
                           n14058, ZN => n1717);
   U607 : OAI22_X1 port map( A1 => n16374, A2 => n14060, B1 => n14074, B2 => 
                           n14059, ZN => n1716);
   U608 : OAI22_X1 port map( A1 => n15886, A2 => n14060, B1 => n14075, B2 => 
                           n14058, ZN => n1715);
   U609 : OAI22_X1 port map( A1 => n16152, A2 => n14060, B1 => n14076, B2 => 
                           n14059, ZN => n1714);
   U610 : OAI22_X1 port map( A1 => n16153, A2 => n14060, B1 => n14077, B2 => 
                           n14058, ZN => n1713);
   U611 : OAI22_X1 port map( A1 => n16622, A2 => n14060, B1 => n14078, B2 => 
                           n14059, ZN => n1712);
   U612 : OAI22_X1 port map( A1 => n16375, A2 => n14060, B1 => n14079, B2 => 
                           n14058, ZN => n1711);
   U613 : OAI22_X1 port map( A1 => n16376, A2 => n14060, B1 => n14080, B2 => 
                           n14059, ZN => n1710);
   U614 : OAI22_X1 port map( A1 => n15887, A2 => n14060, B1 => n14081, B2 => 
                           n14058, ZN => n1709);
   U615 : OAI22_X1 port map( A1 => n16154, A2 => n14060, B1 => n14082, B2 => 
                           n14058, ZN => n1708);
   U616 : OAI22_X1 port map( A1 => n16377, A2 => n14060, B1 => n14083, B2 => 
                           n14059, ZN => n1707);
   U617 : OAI22_X1 port map( A1 => n16155, A2 => n14060, B1 => n14084, B2 => 
                           n14058, ZN => n1706);
   U618 : OAI22_X1 port map( A1 => n16378, A2 => n14060, B1 => n14085, B2 => 
                           n14059, ZN => n1705);
   U619 : OAI22_X1 port map( A1 => n16156, A2 => n14060, B1 => n14086, B2 => 
                           n14058, ZN => n1704);
   U620 : OAI22_X1 port map( A1 => n16379, A2 => n14060, B1 => n14087, B2 => 
                           n14059, ZN => n1703);
   U621 : OAI22_X1 port map( A1 => n16380, A2 => n14060, B1 => n14088, B2 => 
                           n14058, ZN => n1702);
   U622 : OAI22_X1 port map( A1 => n16381, A2 => n14060, B1 => n14089, B2 => 
                           n14058, ZN => n1701);
   U623 : OAI22_X1 port map( A1 => n16623, A2 => n14060, B1 => n14090, B2 => 
                           n14058, ZN => n1700);
   U624 : OAI22_X1 port map( A1 => n16382, A2 => n14060, B1 => n14091, B2 => 
                           n14058, ZN => n1699);
   U625 : OAI22_X1 port map( A1 => n15888, A2 => n14060, B1 => n14092, B2 => 
                           n14058, ZN => n1698);
   U626 : OAI22_X1 port map( A1 => n16624, A2 => n14060, B1 => n14093, B2 => 
                           n14058, ZN => n1697);
   U627 : OAI22_X1 port map( A1 => n16625, A2 => n14060, B1 => n14095, B2 => 
                           n14058, ZN => n1696);
   U628 : OAI22_X1 port map( A1 => n16383, A2 => n14060, B1 => n14096, B2 => 
                           n14059, ZN => n1695);
   U629 : OAI22_X1 port map( A1 => n15889, A2 => n14060, B1 => n14097, B2 => 
                           n14059, ZN => n1694);
   U630 : OAI22_X1 port map( A1 => n16626, A2 => n14060, B1 => n14098, B2 => 
                           n14059, ZN => n1693);
   U631 : OAI22_X1 port map( A1 => n16627, A2 => n14060, B1 => n14099, B2 => 
                           n14059, ZN => n1692);
   U632 : OAI22_X1 port map( A1 => n15890, A2 => n14060, B1 => n14100, B2 => 
                           n14059, ZN => n1691);
   U633 : OAI22_X1 port map( A1 => n16384, A2 => n14060, B1 => n14101, B2 => 
                           n14059, ZN => n1690);
   U634 : OAI22_X1 port map( A1 => n15891, A2 => n14060, B1 => n14102, B2 => 
                           n14059, ZN => n1689);
   U635 : OAI22_X1 port map( A1 => n16628, A2 => n14060, B1 => n14103, B2 => 
                           n14059, ZN => n1688);
   U636 : OAI22_X1 port map( A1 => n16385, A2 => n14060, B1 => n14105, B2 => 
                           n14059, ZN => n1687);
   U637 : NAND2_X1 port map( A1 => n14157, A2 => n14061, ZN => n14062);
   U638 : CLKBUF_X1 port map( A => n14065, Z => n14063);
   U639 : CLKBUF_X1 port map( A => n14062, Z => n14064);
   U640 : OAI22_X1 port map( A1 => n16386, A2 => n14063, B1 => n14121, B2 => 
                           n14064, ZN => n1686);
   U641 : OAI22_X1 port map( A1 => n16387, A2 => n14065, B1 => n14159, B2 => 
                           n14062, ZN => n1685);
   U642 : OAI22_X1 port map( A1 => n16629, A2 => n14063, B1 => n14160, B2 => 
                           n14064, ZN => n1684);
   U643 : OAI22_X1 port map( A1 => n16630, A2 => n14065, B1 => n14161, B2 => 
                           n14062, ZN => n1683);
   U644 : OAI22_X1 port map( A1 => n16388, A2 => n14063, B1 => n14162, B2 => 
                           n14064, ZN => n1682);
   U645 : OAI22_X1 port map( A1 => n16631, A2 => n14065, B1 => n14163, B2 => 
                           n14062, ZN => n1681);
   U646 : OAI22_X1 port map( A1 => n16389, A2 => n14063, B1 => n14164, B2 => 
                           n14064, ZN => n1680);
   U647 : OAI22_X1 port map( A1 => n16390, A2 => n14065, B1 => n14165, B2 => 
                           n14062, ZN => n1679);
   U648 : OAI22_X1 port map( A1 => n16632, A2 => n14063, B1 => n14166, B2 => 
                           n14064, ZN => n1678);
   U649 : OAI22_X1 port map( A1 => n16391, A2 => n14065, B1 => n14167, B2 => 
                           n14062, ZN => n1677);
   U650 : OAI22_X1 port map( A1 => n16392, A2 => n14065, B1 => n14168, B2 => 
                           n14062, ZN => n1676);
   U651 : OAI22_X1 port map( A1 => n16633, A2 => n14065, B1 => n14169, B2 => 
                           n14064, ZN => n1675);
   U652 : OAI22_X1 port map( A1 => n16393, A2 => n14063, B1 => n14170, B2 => 
                           n14062, ZN => n1674);
   U653 : OAI22_X1 port map( A1 => n16634, A2 => n14063, B1 => n14171, B2 => 
                           n14064, ZN => n1673);
   U654 : OAI22_X1 port map( A1 => n16635, A2 => n14063, B1 => n14172, B2 => 
                           n14062, ZN => n1672);
   U655 : OAI22_X1 port map( A1 => n16636, A2 => n14063, B1 => n14173, B2 => 
                           n14064, ZN => n1671);
   U656 : OAI22_X1 port map( A1 => n16637, A2 => n14063, B1 => n14174, B2 => 
                           n14062, ZN => n1670);
   U657 : OAI22_X1 port map( A1 => n16394, A2 => n14063, B1 => n14175, B2 => 
                           n14062, ZN => n1669);
   U658 : OAI22_X1 port map( A1 => n16638, A2 => n14063, B1 => n14176, B2 => 
                           n14062, ZN => n1668);
   U659 : OAI22_X1 port map( A1 => n16639, A2 => n14063, B1 => n14177, B2 => 
                           n14062, ZN => n1667);
   U660 : OAI22_X1 port map( A1 => n16395, A2 => n14063, B1 => n14178, B2 => 
                           n14062, ZN => n1666);
   U661 : OAI22_X1 port map( A1 => n16640, A2 => n14063, B1 => n14179, B2 => 
                           n14062, ZN => n1665);
   U662 : OAI22_X1 port map( A1 => n16641, A2 => n14063, B1 => n14181, B2 => 
                           n14062, ZN => n1664);
   U663 : OAI22_X1 port map( A1 => n16642, A2 => n14063, B1 => n14182, B2 => 
                           n14064, ZN => n1663);
   U664 : OAI22_X1 port map( A1 => n16396, A2 => n14065, B1 => n14183, B2 => 
                           n14064, ZN => n1662);
   U665 : OAI22_X1 port map( A1 => n16397, A2 => n14065, B1 => n14184, B2 => 
                           n14064, ZN => n1661);
   U666 : OAI22_X1 port map( A1 => n16643, A2 => n14065, B1 => n14185, B2 => 
                           n14064, ZN => n1660);
   U667 : OAI22_X1 port map( A1 => n16644, A2 => n14065, B1 => n14186, B2 => 
                           n14064, ZN => n1659);
   U668 : OAI22_X1 port map( A1 => n16645, A2 => n14065, B1 => n14187, B2 => 
                           n14064, ZN => n1658);
   U669 : OAI22_X1 port map( A1 => n16398, A2 => n14065, B1 => n14188, B2 => 
                           n14064, ZN => n1657);
   U670 : OAI22_X1 port map( A1 => n16399, A2 => n14065, B1 => n14189, B2 => 
                           n14064, ZN => n1656);
   U671 : OAI22_X1 port map( A1 => n16400, A2 => n14065, B1 => n14191, B2 => 
                           n14064, ZN => n1655);
   U672 : NOR2_X1 port map( A1 => n14126, A2 => n14066, ZN => n14120);
   U673 : NAND2_X1 port map( A1 => n14127, A2 => n14120, ZN => n14067);
   U674 : CLKBUF_X1 port map( A => n14067, Z => n14068);
   U675 : OAI22_X1 port map( A1 => n16026, A2 => n14069, B1 => n14121, B2 => 
                           n14068, ZN => n1654);
   U676 : OAI22_X1 port map( A1 => n15892, A2 => n14069, B1 => n14073, B2 => 
                           n14067, ZN => n1653);
   U677 : OAI22_X1 port map( A1 => n15893, A2 => n14069, B1 => n14074, B2 => 
                           n14068, ZN => n1652);
   U678 : OAI22_X1 port map( A1 => n15894, A2 => n14069, B1 => n14075, B2 => 
                           n14067, ZN => n1651);
   U679 : OAI22_X1 port map( A1 => n16157, A2 => n14069, B1 => n14076, B2 => 
                           n14068, ZN => n1650);
   U680 : OAI22_X1 port map( A1 => n16158, A2 => n14069, B1 => n14077, B2 => 
                           n14067, ZN => n1649);
   U681 : OAI22_X1 port map( A1 => n16159, A2 => n14069, B1 => n14078, B2 => 
                           n14068, ZN => n1648);
   U682 : OAI22_X1 port map( A1 => n16646, A2 => n14069, B1 => n14079, B2 => 
                           n14067, ZN => n1647);
   U683 : OAI22_X1 port map( A1 => n15895, A2 => n14069, B1 => n14080, B2 => 
                           n14068, ZN => n1646);
   U684 : OAI22_X1 port map( A1 => n15896, A2 => n14069, B1 => n14081, B2 => 
                           n14067, ZN => n1645);
   U685 : OAI22_X1 port map( A1 => n16647, A2 => n14069, B1 => n14082, B2 => 
                           n14067, ZN => n1644);
   U686 : OAI22_X1 port map( A1 => n16160, A2 => n14069, B1 => n14083, B2 => 
                           n14068, ZN => n1643);
   U687 : OAI22_X1 port map( A1 => n16161, A2 => n14069, B1 => n14084, B2 => 
                           n14067, ZN => n1642);
   U688 : OAI22_X1 port map( A1 => n16648, A2 => n14069, B1 => n14085, B2 => 
                           n14068, ZN => n1641);
   U689 : OAI22_X1 port map( A1 => n16162, A2 => n14069, B1 => n14086, B2 => 
                           n14067, ZN => n1640);
   U690 : OAI22_X1 port map( A1 => n16163, A2 => n14069, B1 => n14087, B2 => 
                           n14068, ZN => n1639);
   U691 : OAI22_X1 port map( A1 => n16164, A2 => n14069, B1 => n14088, B2 => 
                           n14067, ZN => n1638);
   U692 : OAI22_X1 port map( A1 => n15897, A2 => n14069, B1 => n14089, B2 => 
                           n14067, ZN => n1637);
   U693 : OAI22_X1 port map( A1 => n16165, A2 => n14069, B1 => n14090, B2 => 
                           n14067, ZN => n1636);
   U694 : OAI22_X1 port map( A1 => n16166, A2 => n14069, B1 => n14091, B2 => 
                           n14067, ZN => n1635);
   U695 : OAI22_X1 port map( A1 => n16167, A2 => n14069, B1 => n14092, B2 => 
                           n14067, ZN => n1634);
   U696 : OAI22_X1 port map( A1 => n15898, A2 => n14069, B1 => n14093, B2 => 
                           n14067, ZN => n1633);
   U697 : OAI22_X1 port map( A1 => n16649, A2 => n14069, B1 => n14095, B2 => 
                           n14067, ZN => n1632);
   U698 : OAI22_X1 port map( A1 => n16168, A2 => n14069, B1 => n14096, B2 => 
                           n14068, ZN => n1631);
   U699 : OAI22_X1 port map( A1 => n16650, A2 => n14069, B1 => n14097, B2 => 
                           n14068, ZN => n1630);
   U700 : OAI22_X1 port map( A1 => n15899, A2 => n14069, B1 => n14098, B2 => 
                           n14068, ZN => n1629);
   U701 : OAI22_X1 port map( A1 => n16169, A2 => n14069, B1 => n14099, B2 => 
                           n14068, ZN => n1628);
   U702 : OAI22_X1 port map( A1 => n15900, A2 => n14069, B1 => n14100, B2 => 
                           n14068, ZN => n1627);
   U703 : OAI22_X1 port map( A1 => n16170, A2 => n14069, B1 => n14101, B2 => 
                           n14068, ZN => n1626);
   U704 : OAI22_X1 port map( A1 => n16171, A2 => n14069, B1 => n14102, B2 => 
                           n14068, ZN => n1625);
   U705 : OAI22_X1 port map( A1 => n15901, A2 => n14069, B1 => n14103, B2 => 
                           n14068, ZN => n1624);
   U706 : OAI22_X1 port map( A1 => n15902, A2 => n14069, B1 => n14105, B2 => 
                           n14068, ZN => n1623);
   U707 : NAND2_X1 port map( A1 => n14131, A2 => n14120, ZN => n14070);
   U708 : CLKBUF_X1 port map( A => n14070, Z => n14071);
   U709 : OAI22_X1 port map( A1 => n16027, A2 => n14072, B1 => n14121, B2 => 
                           n14071, ZN => n1622);
   U710 : OAI22_X1 port map( A1 => n16172, A2 => n14072, B1 => n14159, B2 => 
                           n14070, ZN => n1621);
   U711 : OAI22_X1 port map( A1 => n15903, A2 => n14072, B1 => n14160, B2 => 
                           n14071, ZN => n1620);
   U712 : OAI22_X1 port map( A1 => n16651, A2 => n14072, B1 => n14161, B2 => 
                           n14070, ZN => n1619);
   U713 : OAI22_X1 port map( A1 => n15904, A2 => n14072, B1 => n14162, B2 => 
                           n14071, ZN => n1618);
   U714 : OAI22_X1 port map( A1 => n15905, A2 => n14072, B1 => n14163, B2 => 
                           n14070, ZN => n1617);
   U715 : OAI22_X1 port map( A1 => n15906, A2 => n14072, B1 => n14164, B2 => 
                           n14071, ZN => n1616);
   U716 : OAI22_X1 port map( A1 => n16401, A2 => n14072, B1 => n14165, B2 => 
                           n14070, ZN => n1615);
   U717 : OAI22_X1 port map( A1 => n16652, A2 => n14072, B1 => n14166, B2 => 
                           n14071, ZN => n1614);
   U718 : OAI22_X1 port map( A1 => n16653, A2 => n14072, B1 => n14167, B2 => 
                           n14070, ZN => n1613);
   U719 : OAI22_X1 port map( A1 => n16654, A2 => n14072, B1 => n14168, B2 => 
                           n14070, ZN => n1612);
   U720 : OAI22_X1 port map( A1 => n16655, A2 => n14072, B1 => n14169, B2 => 
                           n14071, ZN => n1611);
   U721 : OAI22_X1 port map( A1 => n16173, A2 => n14072, B1 => n14170, B2 => 
                           n14070, ZN => n1610);
   U722 : OAI22_X1 port map( A1 => n16174, A2 => n14072, B1 => n14171, B2 => 
                           n14071, ZN => n1609);
   U723 : OAI22_X1 port map( A1 => n16656, A2 => n14072, B1 => n14172, B2 => 
                           n14070, ZN => n1608);
   U724 : OAI22_X1 port map( A1 => n16402, A2 => n14072, B1 => n14173, B2 => 
                           n14071, ZN => n1607);
   U725 : OAI22_X1 port map( A1 => n16403, A2 => n14072, B1 => n14174, B2 => 
                           n14070, ZN => n1606);
   U726 : OAI22_X1 port map( A1 => n15907, A2 => n14072, B1 => n14175, B2 => 
                           n14070, ZN => n1605);
   U727 : OAI22_X1 port map( A1 => n16175, A2 => n14072, B1 => n14176, B2 => 
                           n14070, ZN => n1604);
   U728 : OAI22_X1 port map( A1 => n16404, A2 => n14072, B1 => n14177, B2 => 
                           n14070, ZN => n1603);
   U729 : OAI22_X1 port map( A1 => n16657, A2 => n14072, B1 => n14178, B2 => 
                           n14070, ZN => n1602);
   U730 : OAI22_X1 port map( A1 => n16405, A2 => n14072, B1 => n14179, B2 => 
                           n14070, ZN => n1601);
   U731 : OAI22_X1 port map( A1 => n15908, A2 => n14072, B1 => n14181, B2 => 
                           n14070, ZN => n1600);
   U732 : OAI22_X1 port map( A1 => n15909, A2 => n14072, B1 => n14182, B2 => 
                           n14071, ZN => n1599);
   U733 : OAI22_X1 port map( A1 => n16176, A2 => n14072, B1 => n14183, B2 => 
                           n14071, ZN => n1598);
   U734 : OAI22_X1 port map( A1 => n15910, A2 => n14072, B1 => n14184, B2 => 
                           n14071, ZN => n1597);
   U735 : OAI22_X1 port map( A1 => n15911, A2 => n14072, B1 => n14185, B2 => 
                           n14071, ZN => n1596);
   U736 : OAI22_X1 port map( A1 => n16658, A2 => n14072, B1 => n14186, B2 => 
                           n14071, ZN => n1595);
   U737 : OAI22_X1 port map( A1 => n16177, A2 => n14072, B1 => n14187, B2 => 
                           n14071, ZN => n1594);
   U738 : OAI22_X1 port map( A1 => n16659, A2 => n14072, B1 => n14188, B2 => 
                           n14071, ZN => n1593);
   U739 : OAI22_X1 port map( A1 => n16406, A2 => n14072, B1 => n14189, B2 => 
                           n14071, ZN => n1592);
   U740 : OAI22_X1 port map( A1 => n16407, A2 => n14072, B1 => n14191, B2 => 
                           n14071, ZN => n1591);
   U741 : NAND2_X1 port map( A1 => n14135, A2 => n14120, ZN => n14094);
   U742 : CLKBUF_X1 port map( A => n14094, Z => n14104);
   U743 : OAI22_X1 port map( A1 => n15756, A2 => n14106, B1 => n14121, B2 => 
                           n14104, ZN => n1590);
   U744 : OAI22_X1 port map( A1 => n16178, A2 => n14106, B1 => n14073, B2 => 
                           n14094, ZN => n1589);
   U745 : OAI22_X1 port map( A1 => n15912, A2 => n14106, B1 => n14074, B2 => 
                           n14104, ZN => n1588);
   U746 : OAI22_X1 port map( A1 => n16179, A2 => n14106, B1 => n14075, B2 => 
                           n14094, ZN => n1587);
   U747 : OAI22_X1 port map( A1 => n16180, A2 => n14106, B1 => n14076, B2 => 
                           n14104, ZN => n1586);
   U748 : OAI22_X1 port map( A1 => n16181, A2 => n14106, B1 => n14077, B2 => 
                           n14094, ZN => n1585);
   U749 : OAI22_X1 port map( A1 => n15913, A2 => n14106, B1 => n14078, B2 => 
                           n14104, ZN => n1584);
   U750 : OAI22_X1 port map( A1 => n15914, A2 => n14106, B1 => n14079, B2 => 
                           n14094, ZN => n1583);
   U751 : OAI22_X1 port map( A1 => n15915, A2 => n14106, B1 => n14080, B2 => 
                           n14104, ZN => n1582);
   U752 : OAI22_X1 port map( A1 => n15916, A2 => n14106, B1 => n14081, B2 => 
                           n14094, ZN => n1581);
   U753 : OAI22_X1 port map( A1 => n16182, A2 => n14106, B1 => n14082, B2 => 
                           n14094, ZN => n1580);
   U754 : OAI22_X1 port map( A1 => n16408, A2 => n14106, B1 => n14083, B2 => 
                           n14104, ZN => n1579);
   U755 : OAI22_X1 port map( A1 => n15917, A2 => n14106, B1 => n14084, B2 => 
                           n14094, ZN => n1578);
   U756 : OAI22_X1 port map( A1 => n16183, A2 => n14106, B1 => n14085, B2 => 
                           n14104, ZN => n1577);
   U757 : OAI22_X1 port map( A1 => n16409, A2 => n14106, B1 => n14086, B2 => 
                           n14094, ZN => n1576);
   U758 : OAI22_X1 port map( A1 => n16410, A2 => n14106, B1 => n14087, B2 => 
                           n14104, ZN => n1575);
   U759 : OAI22_X1 port map( A1 => n16184, A2 => n14106, B1 => n14088, B2 => 
                           n14094, ZN => n1574);
   U760 : OAI22_X1 port map( A1 => n16660, A2 => n14106, B1 => n14089, B2 => 
                           n14094, ZN => n1573);
   U761 : OAI22_X1 port map( A1 => n16185, A2 => n14106, B1 => n14090, B2 => 
                           n14094, ZN => n1572);
   U762 : OAI22_X1 port map( A1 => n15918, A2 => n14106, B1 => n14091, B2 => 
                           n14094, ZN => n1571);
   U763 : OAI22_X1 port map( A1 => n16411, A2 => n14106, B1 => n14092, B2 => 
                           n14094, ZN => n1570);
   U764 : OAI22_X1 port map( A1 => n16186, A2 => n14106, B1 => n14093, B2 => 
                           n14094, ZN => n1569);
   U765 : OAI22_X1 port map( A1 => n16661, A2 => n14106, B1 => n14095, B2 => 
                           n14094, ZN => n1568);
   U766 : OAI22_X1 port map( A1 => n15919, A2 => n14106, B1 => n14096, B2 => 
                           n14104, ZN => n1567);
   U767 : OAI22_X1 port map( A1 => n15920, A2 => n14106, B1 => n14097, B2 => 
                           n14104, ZN => n1566);
   U768 : OAI22_X1 port map( A1 => n15921, A2 => n14106, B1 => n14098, B2 => 
                           n14104, ZN => n1565);
   U769 : OAI22_X1 port map( A1 => n16412, A2 => n14106, B1 => n14099, B2 => 
                           n14104, ZN => n1564);
   U770 : OAI22_X1 port map( A1 => n15922, A2 => n14106, B1 => n14100, B2 => 
                           n14104, ZN => n1563);
   U771 : OAI22_X1 port map( A1 => n15923, A2 => n14106, B1 => n14101, B2 => 
                           n14104, ZN => n1562);
   U772 : OAI22_X1 port map( A1 => n15924, A2 => n14106, B1 => n14102, B2 => 
                           n14104, ZN => n1561);
   U773 : OAI22_X1 port map( A1 => n16187, A2 => n14106, B1 => n14103, B2 => 
                           n14104, ZN => n1560);
   U774 : OAI22_X1 port map( A1 => n16188, A2 => n14106, B1 => n14105, B2 => 
                           n14104, ZN => n1559);
   U775 : NAND2_X1 port map( A1 => n14139, A2 => n14120, ZN => n14107);
   U776 : CLKBUF_X1 port map( A => n14110, Z => n14108);
   U777 : CLKBUF_X1 port map( A => n14107, Z => n14109);
   U778 : OAI22_X1 port map( A1 => n16271, A2 => n14108, B1 => n14121, B2 => 
                           n14109, ZN => n1558);
   U779 : OAI22_X1 port map( A1 => n16413, A2 => n14110, B1 => n14159, B2 => 
                           n14107, ZN => n1557);
   U780 : OAI22_X1 port map( A1 => n16662, A2 => n14108, B1 => n14160, B2 => 
                           n14109, ZN => n1556);
   U781 : OAI22_X1 port map( A1 => n16189, A2 => n14110, B1 => n14161, B2 => 
                           n14107, ZN => n1555);
   U782 : OAI22_X1 port map( A1 => n16663, A2 => n14108, B1 => n14162, B2 => 
                           n14109, ZN => n1554);
   U783 : OAI22_X1 port map( A1 => n15925, A2 => n14110, B1 => n14163, B2 => 
                           n14107, ZN => n1553);
   U784 : OAI22_X1 port map( A1 => n16664, A2 => n14108, B1 => n14164, B2 => 
                           n14109, ZN => n1552);
   U785 : OAI22_X1 port map( A1 => n16190, A2 => n14110, B1 => n14165, B2 => 
                           n14107, ZN => n1551);
   U786 : OAI22_X1 port map( A1 => n15926, A2 => n14108, B1 => n14166, B2 => 
                           n14109, ZN => n1550);
   U787 : OAI22_X1 port map( A1 => n16665, A2 => n14110, B1 => n14167, B2 => 
                           n14107, ZN => n1549);
   U788 : OAI22_X1 port map( A1 => n16191, A2 => n14110, B1 => n14168, B2 => 
                           n14107, ZN => n1548);
   U789 : OAI22_X1 port map( A1 => n15927, A2 => n14110, B1 => n14169, B2 => 
                           n14109, ZN => n1547);
   U790 : OAI22_X1 port map( A1 => n16666, A2 => n14108, B1 => n14170, B2 => 
                           n14107, ZN => n1546);
   U791 : OAI22_X1 port map( A1 => n15928, A2 => n14108, B1 => n14171, B2 => 
                           n14109, ZN => n1545);
   U792 : OAI22_X1 port map( A1 => n15929, A2 => n14108, B1 => n14172, B2 => 
                           n14107, ZN => n1544);
   U793 : OAI22_X1 port map( A1 => n16192, A2 => n14108, B1 => n14173, B2 => 
                           n14109, ZN => n1543);
   U794 : OAI22_X1 port map( A1 => n15930, A2 => n14108, B1 => n14174, B2 => 
                           n14107, ZN => n1542);
   U795 : OAI22_X1 port map( A1 => n15931, A2 => n14108, B1 => n14175, B2 => 
                           n14107, ZN => n1541);
   U796 : OAI22_X1 port map( A1 => n16667, A2 => n14108, B1 => n14176, B2 => 
                           n14107, ZN => n1540);
   U797 : OAI22_X1 port map( A1 => n16414, A2 => n14108, B1 => n14177, B2 => 
                           n14107, ZN => n1539);
   U798 : OAI22_X1 port map( A1 => n16415, A2 => n14108, B1 => n14178, B2 => 
                           n14107, ZN => n1538);
   U799 : OAI22_X1 port map( A1 => n16416, A2 => n14108, B1 => n14179, B2 => 
                           n14107, ZN => n1537);
   U800 : OAI22_X1 port map( A1 => n16417, A2 => n14108, B1 => n14181, B2 => 
                           n14107, ZN => n1536);
   U801 : OAI22_X1 port map( A1 => n16193, A2 => n14108, B1 => n14182, B2 => 
                           n14109, ZN => n1535);
   U802 : OAI22_X1 port map( A1 => n16194, A2 => n14110, B1 => n14183, B2 => 
                           n14109, ZN => n1534);
   U803 : OAI22_X1 port map( A1 => n16195, A2 => n14110, B1 => n14184, B2 => 
                           n14109, ZN => n1533);
   U804 : OAI22_X1 port map( A1 => n16196, A2 => n14110, B1 => n14185, B2 => 
                           n14109, ZN => n1532);
   U805 : OAI22_X1 port map( A1 => n16418, A2 => n14110, B1 => n14186, B2 => 
                           n14109, ZN => n1531);
   U806 : OAI22_X1 port map( A1 => n16419, A2 => n14110, B1 => n14187, B2 => 
                           n14109, ZN => n1530);
   U807 : OAI22_X1 port map( A1 => n15932, A2 => n14110, B1 => n14188, B2 => 
                           n14109, ZN => n1529);
   U808 : OAI22_X1 port map( A1 => n16668, A2 => n14110, B1 => n14189, B2 => 
                           n14109, ZN => n1528);
   U809 : OAI22_X1 port map( A1 => n15933, A2 => n14110, B1 => n14191, B2 => 
                           n14109, ZN => n1527);
   U810 : NAND2_X1 port map( A1 => n14143, A2 => n14120, ZN => n14111);
   U811 : CLKBUF_X1 port map( A => n14111, Z => n14112);
   U812 : OAI22_X1 port map( A1 => n16028, A2 => n14113, B1 => n14121, B2 => 
                           n14112, ZN => n1526);
   U813 : OAI22_X1 port map( A1 => n15934, A2 => n14113, B1 => n14159, B2 => 
                           n14111, ZN => n1525);
   U814 : OAI22_X1 port map( A1 => n16197, A2 => n14113, B1 => n14160, B2 => 
                           n14112, ZN => n1524);
   U815 : OAI22_X1 port map( A1 => n15935, A2 => n14113, B1 => n14161, B2 => 
                           n14111, ZN => n1523);
   U816 : OAI22_X1 port map( A1 => n15936, A2 => n14113, B1 => n14162, B2 => 
                           n14112, ZN => n1522);
   U817 : OAI22_X1 port map( A1 => n15937, A2 => n14113, B1 => n14163, B2 => 
                           n14111, ZN => n1521);
   U818 : OAI22_X1 port map( A1 => n15938, A2 => n14113, B1 => n14164, B2 => 
                           n14112, ZN => n1520);
   U819 : OAI22_X1 port map( A1 => n16669, A2 => n14113, B1 => n14165, B2 => 
                           n14111, ZN => n1519);
   U820 : OAI22_X1 port map( A1 => n16198, A2 => n14113, B1 => n14166, B2 => 
                           n14112, ZN => n1518);
   U821 : OAI22_X1 port map( A1 => n16420, A2 => n14113, B1 => n14167, B2 => 
                           n14111, ZN => n1517);
   U822 : OAI22_X1 port map( A1 => n15939, A2 => n14113, B1 => n14168, B2 => 
                           n14111, ZN => n1516);
   U823 : OAI22_X1 port map( A1 => n15940, A2 => n14113, B1 => n14169, B2 => 
                           n14112, ZN => n1515);
   U824 : OAI22_X1 port map( A1 => n16199, A2 => n14113, B1 => n14170, B2 => 
                           n14111, ZN => n1514);
   U825 : OAI22_X1 port map( A1 => n15941, A2 => n14113, B1 => n14171, B2 => 
                           n14112, ZN => n1513);
   U826 : OAI22_X1 port map( A1 => n15942, A2 => n14113, B1 => n14172, B2 => 
                           n14111, ZN => n1512);
   U827 : OAI22_X1 port map( A1 => n16670, A2 => n14113, B1 => n14173, B2 => 
                           n14112, ZN => n1511);
   U828 : OAI22_X1 port map( A1 => n15943, A2 => n14113, B1 => n14174, B2 => 
                           n14111, ZN => n1510);
   U829 : OAI22_X1 port map( A1 => n16200, A2 => n14113, B1 => n14175, B2 => 
                           n14111, ZN => n1509);
   U830 : OAI22_X1 port map( A1 => n15944, A2 => n14113, B1 => n14176, B2 => 
                           n14111, ZN => n1508);
   U831 : OAI22_X1 port map( A1 => n16201, A2 => n14113, B1 => n14177, B2 => 
                           n14111, ZN => n1507);
   U832 : OAI22_X1 port map( A1 => n15945, A2 => n14113, B1 => n14178, B2 => 
                           n14111, ZN => n1506);
   U833 : OAI22_X1 port map( A1 => n16202, A2 => n14113, B1 => n14179, B2 => 
                           n14111, ZN => n1505);
   U834 : OAI22_X1 port map( A1 => n16203, A2 => n14113, B1 => n14181, B2 => 
                           n14111, ZN => n1504);
   U835 : OAI22_X1 port map( A1 => n16421, A2 => n14113, B1 => n14182, B2 => 
                           n14112, ZN => n1503);
   U836 : OAI22_X1 port map( A1 => n16204, A2 => n14113, B1 => n14183, B2 => 
                           n14112, ZN => n1502);
   U837 : OAI22_X1 port map( A1 => n15946, A2 => n14113, B1 => n14184, B2 => 
                           n14112, ZN => n1501);
   U838 : OAI22_X1 port map( A1 => n15947, A2 => n14113, B1 => n14185, B2 => 
                           n14112, ZN => n1500);
   U839 : OAI22_X1 port map( A1 => n15948, A2 => n14113, B1 => n14186, B2 => 
                           n14112, ZN => n1499);
   U840 : OAI22_X1 port map( A1 => n15949, A2 => n14113, B1 => n14187, B2 => 
                           n14112, ZN => n1498);
   U841 : OAI22_X1 port map( A1 => n15950, A2 => n14113, B1 => n14188, B2 => 
                           n14112, ZN => n1497);
   U842 : OAI22_X1 port map( A1 => n16205, A2 => n14113, B1 => n14189, B2 => 
                           n14112, ZN => n1496);
   U843 : OAI22_X1 port map( A1 => n15951, A2 => n14113, B1 => n14191, B2 => 
                           n14112, ZN => n1495);
   U844 : NAND2_X1 port map( A1 => n14147, A2 => n14120, ZN => n14114);
   U845 : CLKBUF_X1 port map( A => n14114, Z => n14115);
   U846 : OAI22_X1 port map( A1 => n15757, A2 => n14116, B1 => n14121, B2 => 
                           n14115, ZN => n1494);
   U847 : OAI22_X1 port map( A1 => n16206, A2 => n14116, B1 => n14159, B2 => 
                           n14114, ZN => n1493);
   U848 : OAI22_X1 port map( A1 => n16207, A2 => n14116, B1 => n14160, B2 => 
                           n14115, ZN => n1492);
   U849 : OAI22_X1 port map( A1 => n15952, A2 => n14116, B1 => n14161, B2 => 
                           n14114, ZN => n1491);
   U850 : OAI22_X1 port map( A1 => n16208, A2 => n14116, B1 => n14162, B2 => 
                           n14115, ZN => n1490);
   U851 : OAI22_X1 port map( A1 => n16671, A2 => n14116, B1 => n14163, B2 => 
                           n14114, ZN => n1489);
   U852 : OAI22_X1 port map( A1 => n16422, A2 => n14116, B1 => n14164, B2 => 
                           n14115, ZN => n1488);
   U853 : OAI22_X1 port map( A1 => n15953, A2 => n14116, B1 => n14165, B2 => 
                           n14114, ZN => n1487);
   U854 : OAI22_X1 port map( A1 => n16423, A2 => n14116, B1 => n14166, B2 => 
                           n14115, ZN => n1486);
   U855 : OAI22_X1 port map( A1 => n15954, A2 => n14116, B1 => n14167, B2 => 
                           n14114, ZN => n1485);
   U856 : OAI22_X1 port map( A1 => n15955, A2 => n14116, B1 => n14168, B2 => 
                           n14114, ZN => n1484);
   U857 : OAI22_X1 port map( A1 => n16672, A2 => n14116, B1 => n14169, B2 => 
                           n14115, ZN => n1483);
   U858 : OAI22_X1 port map( A1 => n15956, A2 => n14116, B1 => n14170, B2 => 
                           n14114, ZN => n1482);
   U859 : OAI22_X1 port map( A1 => n15957, A2 => n14116, B1 => n14171, B2 => 
                           n14115, ZN => n1481);
   U860 : OAI22_X1 port map( A1 => n16209, A2 => n14116, B1 => n14172, B2 => 
                           n14114, ZN => n1480);
   U861 : OAI22_X1 port map( A1 => n15958, A2 => n14116, B1 => n14173, B2 => 
                           n14115, ZN => n1479);
   U862 : OAI22_X1 port map( A1 => n15959, A2 => n14116, B1 => n14174, B2 => 
                           n14114, ZN => n1478);
   U863 : OAI22_X1 port map( A1 => n16424, A2 => n14116, B1 => n14175, B2 => 
                           n14114, ZN => n1477);
   U864 : OAI22_X1 port map( A1 => n16673, A2 => n14116, B1 => n14176, B2 => 
                           n14114, ZN => n1476);
   U865 : OAI22_X1 port map( A1 => n15960, A2 => n14116, B1 => n14177, B2 => 
                           n14114, ZN => n1475);
   U866 : OAI22_X1 port map( A1 => n15961, A2 => n14116, B1 => n14178, B2 => 
                           n14114, ZN => n1474);
   U867 : OAI22_X1 port map( A1 => n15962, A2 => n14116, B1 => n14179, B2 => 
                           n14114, ZN => n1473);
   U868 : OAI22_X1 port map( A1 => n16210, A2 => n14116, B1 => n14181, B2 => 
                           n14114, ZN => n1472);
   U869 : OAI22_X1 port map( A1 => n16211, A2 => n14116, B1 => n14182, B2 => 
                           n14115, ZN => n1471);
   U870 : OAI22_X1 port map( A1 => n16674, A2 => n14116, B1 => n14183, B2 => 
                           n14115, ZN => n1470);
   U871 : OAI22_X1 port map( A1 => n15963, A2 => n14116, B1 => n14184, B2 => 
                           n14115, ZN => n1469);
   U872 : OAI22_X1 port map( A1 => n16675, A2 => n14116, B1 => n14185, B2 => 
                           n14115, ZN => n1468);
   U873 : OAI22_X1 port map( A1 => n16676, A2 => n14116, B1 => n14186, B2 => 
                           n14115, ZN => n1467);
   U874 : OAI22_X1 port map( A1 => n16212, A2 => n14116, B1 => n14187, B2 => 
                           n14115, ZN => n1466);
   U875 : OAI22_X1 port map( A1 => n15964, A2 => n14116, B1 => n14188, B2 => 
                           n14115, ZN => n1465);
   U876 : OAI22_X1 port map( A1 => n16425, A2 => n14116, B1 => n14189, B2 => 
                           n14115, ZN => n1464);
   U877 : OAI22_X1 port map( A1 => n15965, A2 => n14116, B1 => n14191, B2 => 
                           n14115, ZN => n1463);
   U878 : NAND2_X1 port map( A1 => n14151, A2 => n14120, ZN => n14117);
   U879 : CLKBUF_X1 port map( A => n14117, Z => n14118);
   U880 : OAI22_X1 port map( A1 => n16272, A2 => n14119, B1 => n14121, B2 => 
                           n14118, ZN => n1462);
   U881 : OAI22_X1 port map( A1 => n15966, A2 => n14119, B1 => n14159, B2 => 
                           n14117, ZN => n1461);
   U882 : OAI22_X1 port map( A1 => n16426, A2 => n14119, B1 => n14160, B2 => 
                           n14118, ZN => n1460);
   U883 : OAI22_X1 port map( A1 => n16677, A2 => n14119, B1 => n14161, B2 => 
                           n14117, ZN => n1459);
   U884 : OAI22_X1 port map( A1 => n16213, A2 => n14119, B1 => n14162, B2 => 
                           n14118, ZN => n1458);
   U885 : OAI22_X1 port map( A1 => n16427, A2 => n14119, B1 => n14163, B2 => 
                           n14117, ZN => n1457);
   U886 : OAI22_X1 port map( A1 => n16428, A2 => n14119, B1 => n14164, B2 => 
                           n14118, ZN => n1456);
   U887 : OAI22_X1 port map( A1 => n15967, A2 => n14119, B1 => n14165, B2 => 
                           n14117, ZN => n1455);
   U888 : OAI22_X1 port map( A1 => n16678, A2 => n14119, B1 => n14166, B2 => 
                           n14118, ZN => n1454);
   U889 : OAI22_X1 port map( A1 => n16429, A2 => n14119, B1 => n14167, B2 => 
                           n14117, ZN => n1453);
   U890 : OAI22_X1 port map( A1 => n16214, A2 => n14119, B1 => n14168, B2 => 
                           n14117, ZN => n1452);
   U891 : OAI22_X1 port map( A1 => n16215, A2 => n14119, B1 => n14169, B2 => 
                           n14118, ZN => n1451);
   U892 : OAI22_X1 port map( A1 => n16430, A2 => n14119, B1 => n14170, B2 => 
                           n14117, ZN => n1450);
   U893 : OAI22_X1 port map( A1 => n16431, A2 => n14119, B1 => n14171, B2 => 
                           n14118, ZN => n1449);
   U894 : OAI22_X1 port map( A1 => n16432, A2 => n14119, B1 => n14172, B2 => 
                           n14117, ZN => n1448);
   U895 : OAI22_X1 port map( A1 => n16679, A2 => n14119, B1 => n14173, B2 => 
                           n14118, ZN => n1447);
   U896 : OAI22_X1 port map( A1 => n16680, A2 => n14119, B1 => n14174, B2 => 
                           n14117, ZN => n1446);
   U897 : OAI22_X1 port map( A1 => n16681, A2 => n14119, B1 => n14175, B2 => 
                           n14117, ZN => n1445);
   U898 : OAI22_X1 port map( A1 => n16433, A2 => n14119, B1 => n14176, B2 => 
                           n14117, ZN => n1444);
   U899 : OAI22_X1 port map( A1 => n16682, A2 => n14119, B1 => n14177, B2 => 
                           n14117, ZN => n1443);
   U900 : OAI22_X1 port map( A1 => n16216, A2 => n14119, B1 => n14178, B2 => 
                           n14117, ZN => n1442);
   U901 : OAI22_X1 port map( A1 => n15968, A2 => n14119, B1 => n14179, B2 => 
                           n14117, ZN => n1441);
   U902 : OAI22_X1 port map( A1 => n16434, A2 => n14119, B1 => n14181, B2 => 
                           n14117, ZN => n1440);
   U903 : OAI22_X1 port map( A1 => n16683, A2 => n14119, B1 => n14182, B2 => 
                           n14118, ZN => n1439);
   U904 : OAI22_X1 port map( A1 => n16684, A2 => n14119, B1 => n14183, B2 => 
                           n14118, ZN => n1438);
   U905 : OAI22_X1 port map( A1 => n16685, A2 => n14119, B1 => n14184, B2 => 
                           n14118, ZN => n1437);
   U906 : OAI22_X1 port map( A1 => n16435, A2 => n14119, B1 => n14185, B2 => 
                           n14118, ZN => n1436);
   U907 : OAI22_X1 port map( A1 => n16686, A2 => n14119, B1 => n14186, B2 => 
                           n14118, ZN => n1435);
   U908 : OAI22_X1 port map( A1 => n16436, A2 => n14119, B1 => n14187, B2 => 
                           n14118, ZN => n1434);
   U909 : OAI22_X1 port map( A1 => n16437, A2 => n14119, B1 => n14188, B2 => 
                           n14118, ZN => n1433);
   U910 : OAI22_X1 port map( A1 => n16687, A2 => n14119, B1 => n14189, B2 => 
                           n14118, ZN => n1432);
   U911 : OAI22_X1 port map( A1 => n16688, A2 => n14119, B1 => n14191, B2 => 
                           n14118, ZN => n1431);
   U912 : NAND2_X1 port map( A1 => n14157, A2 => n14120, ZN => n14122);
   U913 : OAI22_X1 port map( A1 => n16273, A2 => n14124, B1 => n14121, B2 => 
                           n14123, ZN => n1430);
   U914 : OAI22_X1 port map( A1 => n16438, A2 => n14124, B1 => n14159, B2 => 
                           n14122, ZN => n1429);
   U915 : OAI22_X1 port map( A1 => n16689, A2 => n14124, B1 => n14160, B2 => 
                           n14123, ZN => n1428);
   U916 : OAI22_X1 port map( A1 => n16439, A2 => n14124, B1 => n14161, B2 => 
                           n14122, ZN => n1427);
   U917 : OAI22_X1 port map( A1 => n16440, A2 => n14124, B1 => n14162, B2 => 
                           n14123, ZN => n1426);
   U918 : OAI22_X1 port map( A1 => n16441, A2 => n14124, B1 => n14163, B2 => 
                           n14122, ZN => n1425);
   U919 : OAI22_X1 port map( A1 => n16690, A2 => n14124, B1 => n14164, B2 => 
                           n14123, ZN => n1424);
   U920 : OAI22_X1 port map( A1 => n16691, A2 => n14124, B1 => n14165, B2 => 
                           n14122, ZN => n1423);
   U921 : OAI22_X1 port map( A1 => n16442, A2 => n14124, B1 => n14166, B2 => 
                           n14123, ZN => n1422);
   U922 : OAI22_X1 port map( A1 => n16692, A2 => n14124, B1 => n14167, B2 => 
                           n14122, ZN => n1421);
   U923 : OAI22_X1 port map( A1 => n16443, A2 => n14124, B1 => n14168, B2 => 
                           n14122, ZN => n1420);
   U924 : OAI22_X1 port map( A1 => n16444, A2 => n14124, B1 => n14169, B2 => 
                           n14123, ZN => n1419);
   U925 : OAI22_X1 port map( A1 => n16693, A2 => n14124, B1 => n14170, B2 => 
                           n14122, ZN => n1418);
   U926 : OAI22_X1 port map( A1 => n16445, A2 => n14124, B1 => n14171, B2 => 
                           n14123, ZN => n1417);
   U927 : OAI22_X1 port map( A1 => n16694, A2 => n14124, B1 => n14172, B2 => 
                           n14122, ZN => n1416);
   U928 : OAI22_X1 port map( A1 => n16446, A2 => n14124, B1 => n14173, B2 => 
                           n14123, ZN => n1415);
   U929 : OAI22_X1 port map( A1 => n16695, A2 => n14124, B1 => n14174, B2 => 
                           n14122, ZN => n1414);
   U930 : OAI22_X1 port map( A1 => n16447, A2 => n14124, B1 => n14175, B2 => 
                           n14122, ZN => n1413);
   U931 : OAI22_X1 port map( A1 => n16448, A2 => n14124, B1 => n14176, B2 => 
                           n14122, ZN => n1412);
   U932 : OAI22_X1 port map( A1 => n16449, A2 => n14124, B1 => n14177, B2 => 
                           n14122, ZN => n1411);
   U933 : OAI22_X1 port map( A1 => n16450, A2 => n14124, B1 => n14178, B2 => 
                           n14122, ZN => n1410);
   U934 : OAI22_X1 port map( A1 => n16696, A2 => n14124, B1 => n14179, B2 => 
                           n14122, ZN => n1409);
   U935 : OAI22_X1 port map( A1 => n16451, A2 => n14124, B1 => n14181, B2 => 
                           n14122, ZN => n1408);
   U936 : OAI22_X1 port map( A1 => n16452, A2 => n14124, B1 => n14182, B2 => 
                           n14123, ZN => n1407);
   U937 : OAI22_X1 port map( A1 => n16453, A2 => n14124, B1 => n14183, B2 => 
                           n14123, ZN => n1406);
   U938 : OAI22_X1 port map( A1 => n16454, A2 => n14124, B1 => n14184, B2 => 
                           n14123, ZN => n1405);
   U939 : OAI22_X1 port map( A1 => n16455, A2 => n14124, B1 => n14185, B2 => 
                           n14123, ZN => n1404);
   U940 : OAI22_X1 port map( A1 => n16697, A2 => n14124, B1 => n14186, B2 => 
                           n14123, ZN => n1403);
   U941 : OAI22_X1 port map( A1 => n16698, A2 => n14124, B1 => n14187, B2 => 
                           n14123, ZN => n1402);
   U942 : OAI22_X1 port map( A1 => n16699, A2 => n14124, B1 => n14188, B2 => 
                           n14123, ZN => n1401);
   U943 : OAI22_X1 port map( A1 => n16700, A2 => n14124, B1 => n14189, B2 => 
                           n14123, ZN => n1400);
   U944 : OAI22_X1 port map( A1 => n16701, A2 => n14124, B1 => n14191, B2 => 
                           n14123, ZN => n1399);
   U945 : NOR2_X1 port map( A1 => n14126, A2 => n14125, ZN => n14156);
   U946 : NAND2_X1 port map( A1 => n14127, A2 => n14156, ZN => n14128);
   U947 : CLKBUF_X1 port map( A => n14128, Z => n14129);
   U948 : OAI22_X1 port map( A1 => n16029, A2 => n14130, B1 => n14158, B2 => 
                           n14129, ZN => n1398);
   U949 : OAI22_X1 port map( A1 => n15969, A2 => n14130, B1 => n14159, B2 => 
                           n14128, ZN => n1397);
   U950 : OAI22_X1 port map( A1 => n15970, A2 => n14130, B1 => n14160, B2 => 
                           n14129, ZN => n1396);
   U951 : OAI22_X1 port map( A1 => n15971, A2 => n14130, B1 => n14161, B2 => 
                           n14128, ZN => n1395);
   U952 : OAI22_X1 port map( A1 => n16217, A2 => n14130, B1 => n14162, B2 => 
                           n14129, ZN => n1394);
   U953 : OAI22_X1 port map( A1 => n15972, A2 => n14130, B1 => n14163, B2 => 
                           n14128, ZN => n1393);
   U954 : OAI22_X1 port map( A1 => n16218, A2 => n14130, B1 => n14164, B2 => 
                           n14129, ZN => n1392);
   U955 : OAI22_X1 port map( A1 => n15973, A2 => n14130, B1 => n14165, B2 => 
                           n14128, ZN => n1391);
   U956 : OAI22_X1 port map( A1 => n16219, A2 => n14130, B1 => n14166, B2 => 
                           n14129, ZN => n1390);
   U957 : OAI22_X1 port map( A1 => n16220, A2 => n14130, B1 => n14167, B2 => 
                           n14128, ZN => n1389);
   U958 : OAI22_X1 port map( A1 => n15974, A2 => n14130, B1 => n14168, B2 => 
                           n14128, ZN => n1388);
   U959 : OAI22_X1 port map( A1 => n15975, A2 => n14130, B1 => n14169, B2 => 
                           n14129, ZN => n1387);
   U960 : OAI22_X1 port map( A1 => n16221, A2 => n14130, B1 => n14170, B2 => 
                           n14128, ZN => n1386);
   U961 : OAI22_X1 port map( A1 => n15976, A2 => n14130, B1 => n14171, B2 => 
                           n14129, ZN => n1385);
   U962 : OAI22_X1 port map( A1 => n16222, A2 => n14130, B1 => n14172, B2 => 
                           n14128, ZN => n1384);
   U963 : OAI22_X1 port map( A1 => n15977, A2 => n14130, B1 => n14173, B2 => 
                           n14129, ZN => n1383);
   U964 : OAI22_X1 port map( A1 => n16223, A2 => n14130, B1 => n14174, B2 => 
                           n14128, ZN => n1382);
   U965 : OAI22_X1 port map( A1 => n15978, A2 => n14130, B1 => n14175, B2 => 
                           n14128, ZN => n1381);
   U966 : OAI22_X1 port map( A1 => n15979, A2 => n14130, B1 => n14176, B2 => 
                           n14128, ZN => n1380);
   U967 : OAI22_X1 port map( A1 => n15980, A2 => n14130, B1 => n14177, B2 => 
                           n14128, ZN => n1379);
   U968 : OAI22_X1 port map( A1 => n16224, A2 => n14130, B1 => n14178, B2 => 
                           n14128, ZN => n1378);
   U969 : OAI22_X1 port map( A1 => n15981, A2 => n14130, B1 => n14179, B2 => 
                           n14128, ZN => n1377);
   U970 : OAI22_X1 port map( A1 => n15982, A2 => n14130, B1 => n14181, B2 => 
                           n14128, ZN => n1376);
   U971 : OAI22_X1 port map( A1 => n15983, A2 => n14130, B1 => n14182, B2 => 
                           n14129, ZN => n1375);
   U972 : OAI22_X1 port map( A1 => n15984, A2 => n14130, B1 => n14183, B2 => 
                           n14129, ZN => n1374);
   U973 : OAI22_X1 port map( A1 => n16456, A2 => n14130, B1 => n14184, B2 => 
                           n14129, ZN => n1373);
   U974 : OAI22_X1 port map( A1 => n16225, A2 => n14130, B1 => n14185, B2 => 
                           n14129, ZN => n1372);
   U975 : OAI22_X1 port map( A1 => n16226, A2 => n14130, B1 => n14186, B2 => 
                           n14129, ZN => n1371);
   U976 : OAI22_X1 port map( A1 => n16702, A2 => n14130, B1 => n14187, B2 => 
                           n14129, ZN => n1370);
   U977 : OAI22_X1 port map( A1 => n16227, A2 => n14130, B1 => n14188, B2 => 
                           n14129, ZN => n1369);
   U978 : OAI22_X1 port map( A1 => n15985, A2 => n14130, B1 => n14189, B2 => 
                           n14129, ZN => n1368);
   U979 : OAI22_X1 port map( A1 => n16228, A2 => n14130, B1 => n14191, B2 => 
                           n14129, ZN => n1367);
   U980 : NAND2_X1 port map( A1 => n14131, A2 => n14156, ZN => n14132);
   U981 : CLKBUF_X1 port map( A => n14132, Z => n14133);
   U982 : OAI22_X1 port map( A1 => n16030, A2 => n14134, B1 => n14158, B2 => 
                           n14133, ZN => n1366);
   U983 : OAI22_X1 port map( A1 => n16457, A2 => n14134, B1 => n14159, B2 => 
                           n14132, ZN => n1365);
   U984 : OAI22_X1 port map( A1 => n16703, A2 => n14134, B1 => n14160, B2 => 
                           n14133, ZN => n1364);
   U985 : OAI22_X1 port map( A1 => n16704, A2 => n14134, B1 => n14161, B2 => 
                           n14132, ZN => n1363);
   U986 : OAI22_X1 port map( A1 => n16458, A2 => n14134, B1 => n14162, B2 => 
                           n14133, ZN => n1362);
   U987 : OAI22_X1 port map( A1 => n16229, A2 => n14134, B1 => n14163, B2 => 
                           n14132, ZN => n1361);
   U988 : OAI22_X1 port map( A1 => n16230, A2 => n14134, B1 => n14164, B2 => 
                           n14133, ZN => n1360);
   U989 : OAI22_X1 port map( A1 => n16231, A2 => n14134, B1 => n14165, B2 => 
                           n14132, ZN => n1359);
   U990 : OAI22_X1 port map( A1 => n16232, A2 => n14134, B1 => n14166, B2 => 
                           n14133, ZN => n1358);
   U991 : OAI22_X1 port map( A1 => n16459, A2 => n14134, B1 => n14167, B2 => 
                           n14132, ZN => n1357);
   U992 : OAI22_X1 port map( A1 => n16705, A2 => n14134, B1 => n14168, B2 => 
                           n14132, ZN => n1356);
   U993 : OAI22_X1 port map( A1 => n16233, A2 => n14134, B1 => n14169, B2 => 
                           n14133, ZN => n1355);
   U994 : OAI22_X1 port map( A1 => n16234, A2 => n14134, B1 => n14170, B2 => 
                           n14132, ZN => n1354);
   U995 : OAI22_X1 port map( A1 => n16460, A2 => n14134, B1 => n14171, B2 => 
                           n14133, ZN => n1353);
   U996 : OAI22_X1 port map( A1 => n15986, A2 => n14134, B1 => n14172, B2 => 
                           n14132, ZN => n1352);
   U997 : OAI22_X1 port map( A1 => n15987, A2 => n14134, B1 => n14173, B2 => 
                           n14133, ZN => n1351);
   U998 : OAI22_X1 port map( A1 => n16461, A2 => n14134, B1 => n14174, B2 => 
                           n14132, ZN => n1350);
   U999 : OAI22_X1 port map( A1 => n16235, A2 => n14134, B1 => n14175, B2 => 
                           n14132, ZN => n1349);
   U1000 : OAI22_X1 port map( A1 => n16706, A2 => n14134, B1 => n14176, B2 => 
                           n14132, ZN => n1348);
   U1001 : OAI22_X1 port map( A1 => n15988, A2 => n14134, B1 => n14177, B2 => 
                           n14132, ZN => n1347);
   U1002 : OAI22_X1 port map( A1 => n15989, A2 => n14134, B1 => n14178, B2 => 
                           n14132, ZN => n1346);
   U1003 : OAI22_X1 port map( A1 => n16707, A2 => n14134, B1 => n14179, B2 => 
                           n14132, ZN => n1345);
   U1004 : OAI22_X1 port map( A1 => n16236, A2 => n14134, B1 => n14181, B2 => 
                           n14132, ZN => n1344);
   U1005 : OAI22_X1 port map( A1 => n16462, A2 => n14134, B1 => n14182, B2 => 
                           n14133, ZN => n1343);
   U1006 : OAI22_X1 port map( A1 => n16237, A2 => n14134, B1 => n14183, B2 => 
                           n14133, ZN => n1342);
   U1007 : OAI22_X1 port map( A1 => n16708, A2 => n14134, B1 => n14184, B2 => 
                           n14133, ZN => n1341);
   U1008 : OAI22_X1 port map( A1 => n16238, A2 => n14134, B1 => n14185, B2 => 
                           n14133, ZN => n1340);
   U1009 : OAI22_X1 port map( A1 => n16239, A2 => n14134, B1 => n14186, B2 => 
                           n14133, ZN => n1339);
   U1010 : OAI22_X1 port map( A1 => n16709, A2 => n14134, B1 => n14187, B2 => 
                           n14133, ZN => n1338);
   U1011 : OAI22_X1 port map( A1 => n15990, A2 => n14134, B1 => n14188, B2 => 
                           n14133, ZN => n1337);
   U1012 : OAI22_X1 port map( A1 => n15991, A2 => n14134, B1 => n14189, B2 => 
                           n14133, ZN => n1336);
   U1013 : OAI22_X1 port map( A1 => n16463, A2 => n14134, B1 => n14191, B2 => 
                           n14133, ZN => n1335);
   U1014 : NAND2_X1 port map( A1 => n14135, A2 => n14156, ZN => n14136);
   U1015 : CLKBUF_X1 port map( A => n14136, Z => n14137);
   U1016 : OAI22_X1 port map( A1 => n15758, A2 => n14138, B1 => n14158, B2 => 
                           n14137, ZN => n1334);
   U1017 : OAI22_X1 port map( A1 => n16710, A2 => n14138, B1 => n14159, B2 => 
                           n14136, ZN => n1333);
   U1018 : OAI22_X1 port map( A1 => n16464, A2 => n14138, B1 => n14160, B2 => 
                           n14137, ZN => n1332);
   U1019 : OAI22_X1 port map( A1 => n16711, A2 => n14138, B1 => n14161, B2 => 
                           n14136, ZN => n1331);
   U1020 : OAI22_X1 port map( A1 => n16712, A2 => n14138, B1 => n14162, B2 => 
                           n14137, ZN => n1330);
   U1021 : OAI22_X1 port map( A1 => n16465, A2 => n14138, B1 => n14163, B2 => 
                           n14136, ZN => n1329);
   U1022 : OAI22_X1 port map( A1 => n16466, A2 => n14138, B1 => n14164, B2 => 
                           n14137, ZN => n1328);
   U1023 : OAI22_X1 port map( A1 => n15992, A2 => n14138, B1 => n14165, B2 => 
                           n14136, ZN => n1327);
   U1024 : OAI22_X1 port map( A1 => n16467, A2 => n14138, B1 => n14166, B2 => 
                           n14137, ZN => n1326);
   U1025 : OAI22_X1 port map( A1 => n16240, A2 => n14138, B1 => n14167, B2 => 
                           n14136, ZN => n1325);
   U1026 : OAI22_X1 port map( A1 => n16713, A2 => n14138, B1 => n14168, B2 => 
                           n14136, ZN => n1324);
   U1027 : OAI22_X1 port map( A1 => n16468, A2 => n14138, B1 => n14169, B2 => 
                           n14137, ZN => n1323);
   U1028 : OAI22_X1 port map( A1 => n16469, A2 => n14138, B1 => n14170, B2 => 
                           n14136, ZN => n1322);
   U1029 : OAI22_X1 port map( A1 => n16714, A2 => n14138, B1 => n14171, B2 => 
                           n14137, ZN => n1321);
   U1030 : OAI22_X1 port map( A1 => n16715, A2 => n14138, B1 => n14172, B2 => 
                           n14136, ZN => n1320);
   U1031 : OAI22_X1 port map( A1 => n15993, A2 => n14138, B1 => n14173, B2 => 
                           n14137, ZN => n1319);
   U1032 : OAI22_X1 port map( A1 => n16716, A2 => n14138, B1 => n14174, B2 => 
                           n14136, ZN => n1318);
   U1033 : OAI22_X1 port map( A1 => n16717, A2 => n14138, B1 => n14175, B2 => 
                           n14136, ZN => n1317);
   U1034 : OAI22_X1 port map( A1 => n16241, A2 => n14138, B1 => n14176, B2 => 
                           n14136, ZN => n1316);
   U1035 : OAI22_X1 port map( A1 => n16718, A2 => n14138, B1 => n14177, B2 => 
                           n14136, ZN => n1315);
   U1036 : OAI22_X1 port map( A1 => n16719, A2 => n14138, B1 => n14178, B2 => 
                           n14136, ZN => n1314);
   U1037 : OAI22_X1 port map( A1 => n16720, A2 => n14138, B1 => n14179, B2 => 
                           n14136, ZN => n1313);
   U1038 : OAI22_X1 port map( A1 => n16721, A2 => n14138, B1 => n14181, B2 => 
                           n14136, ZN => n1312);
   U1039 : OAI22_X1 port map( A1 => n16242, A2 => n14138, B1 => n14182, B2 => 
                           n14137, ZN => n1311);
   U1040 : OAI22_X1 port map( A1 => n16470, A2 => n14138, B1 => n14183, B2 => 
                           n14137, ZN => n1310);
   U1041 : OAI22_X1 port map( A1 => n16722, A2 => n14138, B1 => n14184, B2 => 
                           n14137, ZN => n1309);
   U1042 : OAI22_X1 port map( A1 => n16723, A2 => n14138, B1 => n14185, B2 => 
                           n14137, ZN => n1308);
   U1043 : OAI22_X1 port map( A1 => n15994, A2 => n14138, B1 => n14186, B2 => 
                           n14137, ZN => n1307);
   U1044 : OAI22_X1 port map( A1 => n16243, A2 => n14138, B1 => n14187, B2 => 
                           n14137, ZN => n1306);
   U1045 : OAI22_X1 port map( A1 => n16471, A2 => n14138, B1 => n14188, B2 => 
                           n14137, ZN => n1305);
   U1046 : OAI22_X1 port map( A1 => n16244, A2 => n14138, B1 => n14189, B2 => 
                           n14137, ZN => n1304);
   U1047 : OAI22_X1 port map( A1 => n16724, A2 => n14138, B1 => n14191, B2 => 
                           n14137, ZN => n1303);
   U1048 : NAND2_X1 port map( A1 => n14139, A2 => n14156, ZN => n14140);
   U1049 : CLKBUF_X1 port map( A => n14140, Z => n14141);
   U1050 : OAI22_X1 port map( A1 => n15759, A2 => n14142, B1 => n14158, B2 => 
                           n14141, ZN => n1302);
   U1051 : OAI22_X1 port map( A1 => n16725, A2 => n14142, B1 => n14159, B2 => 
                           n14140, ZN => n1301);
   U1052 : OAI22_X1 port map( A1 => n16726, A2 => n14142, B1 => n14160, B2 => 
                           n14141, ZN => n1300);
   U1053 : OAI22_X1 port map( A1 => n16727, A2 => n14142, B1 => n14161, B2 => 
                           n14140, ZN => n1299);
   U1054 : OAI22_X1 port map( A1 => n16472, A2 => n14142, B1 => n14162, B2 => 
                           n14141, ZN => n1298);
   U1055 : OAI22_X1 port map( A1 => n16728, A2 => n14142, B1 => n14163, B2 => 
                           n14140, ZN => n1297);
   U1056 : OAI22_X1 port map( A1 => n16729, A2 => n14142, B1 => n14164, B2 => 
                           n14141, ZN => n1296);
   U1057 : OAI22_X1 port map( A1 => n16730, A2 => n14142, B1 => n14165, B2 => 
                           n14140, ZN => n1295);
   U1058 : OAI22_X1 port map( A1 => n16245, A2 => n14142, B1 => n14166, B2 => 
                           n14141, ZN => n1294);
   U1059 : OAI22_X1 port map( A1 => n16731, A2 => n14142, B1 => n14167, B2 => 
                           n14140, ZN => n1293);
   U1060 : OAI22_X1 port map( A1 => n16473, A2 => n14142, B1 => n14168, B2 => 
                           n14140, ZN => n1292);
   U1061 : OAI22_X1 port map( A1 => n16732, A2 => n14142, B1 => n14169, B2 => 
                           n14141, ZN => n1291);
   U1062 : OAI22_X1 port map( A1 => n16733, A2 => n14142, B1 => n14170, B2 => 
                           n14140, ZN => n1290);
   U1063 : OAI22_X1 port map( A1 => n16246, A2 => n14142, B1 => n14171, B2 => 
                           n14141, ZN => n1289);
   U1064 : OAI22_X1 port map( A1 => n16474, A2 => n14142, B1 => n14172, B2 => 
                           n14140, ZN => n1288);
   U1065 : OAI22_X1 port map( A1 => n16734, A2 => n14142, B1 => n14173, B2 => 
                           n14141, ZN => n1287);
   U1066 : OAI22_X1 port map( A1 => n16475, A2 => n14142, B1 => n14174, B2 => 
                           n14140, ZN => n1286);
   U1067 : OAI22_X1 port map( A1 => n16476, A2 => n14142, B1 => n14175, B2 => 
                           n14140, ZN => n1285);
   U1068 : OAI22_X1 port map( A1 => n16735, A2 => n14142, B1 => n14176, B2 => 
                           n14140, ZN => n1284);
   U1069 : OAI22_X1 port map( A1 => n16736, A2 => n14142, B1 => n14177, B2 => 
                           n14140, ZN => n1283);
   U1070 : OAI22_X1 port map( A1 => n16477, A2 => n14142, B1 => n14178, B2 => 
                           n14140, ZN => n1282);
   U1071 : OAI22_X1 port map( A1 => n16478, A2 => n14142, B1 => n14179, B2 => 
                           n14140, ZN => n1281);
   U1072 : OAI22_X1 port map( A1 => n15995, A2 => n14142, B1 => n14181, B2 => 
                           n14140, ZN => n1280);
   U1073 : OAI22_X1 port map( A1 => n16737, A2 => n14142, B1 => n14182, B2 => 
                           n14141, ZN => n1279);
   U1074 : OAI22_X1 port map( A1 => n15996, A2 => n14142, B1 => n14183, B2 => 
                           n14141, ZN => n1278);
   U1075 : OAI22_X1 port map( A1 => n16479, A2 => n14142, B1 => n14184, B2 => 
                           n14141, ZN => n1277);
   U1076 : OAI22_X1 port map( A1 => n15997, A2 => n14142, B1 => n14185, B2 => 
                           n14141, ZN => n1276);
   U1077 : OAI22_X1 port map( A1 => n16247, A2 => n14142, B1 => n14186, B2 => 
                           n14141, ZN => n1275);
   U1078 : OAI22_X1 port map( A1 => n16480, A2 => n14142, B1 => n14187, B2 => 
                           n14141, ZN => n1274);
   U1079 : OAI22_X1 port map( A1 => n16738, A2 => n14142, B1 => n14188, B2 => 
                           n14141, ZN => n1273);
   U1080 : OAI22_X1 port map( A1 => n16481, A2 => n14142, B1 => n14189, B2 => 
                           n14141, ZN => n1272);
   U1081 : OAI22_X1 port map( A1 => n16739, A2 => n14142, B1 => n14191, B2 => 
                           n14141, ZN => n1271);
   U1082 : NAND2_X1 port map( A1 => n14143, A2 => n14156, ZN => n14144);
   U1083 : CLKBUF_X1 port map( A => n14144, Z => n14145);
   U1084 : OAI22_X1 port map( A1 => n16274, A2 => n14146, B1 => n14158, B2 => 
                           n14145, ZN => n1270);
   U1085 : OAI22_X1 port map( A1 => n16740, A2 => n14146, B1 => n14159, B2 => 
                           n14144, ZN => n1269);
   U1086 : OAI22_X1 port map( A1 => n16482, A2 => n14146, B1 => n14160, B2 => 
                           n14145, ZN => n1268);
   U1087 : OAI22_X1 port map( A1 => n16483, A2 => n14146, B1 => n14161, B2 => 
                           n14144, ZN => n1267);
   U1088 : OAI22_X1 port map( A1 => n16484, A2 => n14146, B1 => n14162, B2 => 
                           n14145, ZN => n1266);
   U1089 : OAI22_X1 port map( A1 => n16741, A2 => n14146, B1 => n14163, B2 => 
                           n14144, ZN => n1265);
   U1090 : OAI22_X1 port map( A1 => n16485, A2 => n14146, B1 => n14164, B2 => 
                           n14145, ZN => n1264);
   U1091 : OAI22_X1 port map( A1 => n16742, A2 => n14146, B1 => n14165, B2 => 
                           n14144, ZN => n1263);
   U1092 : OAI22_X1 port map( A1 => n16743, A2 => n14146, B1 => n14166, B2 => 
                           n14145, ZN => n1262);
   U1093 : OAI22_X1 port map( A1 => n15998, A2 => n14146, B1 => n14167, B2 => 
                           n14144, ZN => n1261);
   U1094 : OAI22_X1 port map( A1 => n16486, A2 => n14146, B1 => n14168, B2 => 
                           n14144, ZN => n1260);
   U1095 : OAI22_X1 port map( A1 => n16744, A2 => n14146, B1 => n14169, B2 => 
                           n14145, ZN => n1259);
   U1096 : OAI22_X1 port map( A1 => n16487, A2 => n14146, B1 => n14170, B2 => 
                           n14144, ZN => n1258);
   U1097 : OAI22_X1 port map( A1 => n16745, A2 => n14146, B1 => n14171, B2 => 
                           n14145, ZN => n1257);
   U1098 : OAI22_X1 port map( A1 => n16746, A2 => n14146, B1 => n14172, B2 => 
                           n14144, ZN => n1256);
   U1099 : OAI22_X1 port map( A1 => n16747, A2 => n14146, B1 => n14173, B2 => 
                           n14145, ZN => n1255);
   U1100 : OAI22_X1 port map( A1 => n15999, A2 => n14146, B1 => n14174, B2 => 
                           n14144, ZN => n1254);
   U1101 : OAI22_X1 port map( A1 => n16748, A2 => n14146, B1 => n14175, B2 => 
                           n14144, ZN => n1253);
   U1102 : OAI22_X1 port map( A1 => n16488, A2 => n14146, B1 => n14176, B2 => 
                           n14144, ZN => n1252);
   U1103 : OAI22_X1 port map( A1 => n16749, A2 => n14146, B1 => n14177, B2 => 
                           n14144, ZN => n1251);
   U1104 : OAI22_X1 port map( A1 => n16750, A2 => n14146, B1 => n14178, B2 => 
                           n14144, ZN => n1250);
   U1105 : OAI22_X1 port map( A1 => n16751, A2 => n14146, B1 => n14179, B2 => 
                           n14144, ZN => n1249);
   U1106 : OAI22_X1 port map( A1 => n16752, A2 => n14146, B1 => n14181, B2 => 
                           n14144, ZN => n1248);
   U1107 : OAI22_X1 port map( A1 => n16753, A2 => n14146, B1 => n14182, B2 => 
                           n14145, ZN => n1247);
   U1108 : OAI22_X1 port map( A1 => n16489, A2 => n14146, B1 => n14183, B2 => 
                           n14145, ZN => n1246);
   U1109 : OAI22_X1 port map( A1 => n16754, A2 => n14146, B1 => n14184, B2 => 
                           n14145, ZN => n1245);
   U1110 : OAI22_X1 port map( A1 => n16755, A2 => n14146, B1 => n14185, B2 => 
                           n14145, ZN => n1244);
   U1111 : OAI22_X1 port map( A1 => n16490, A2 => n14146, B1 => n14186, B2 => 
                           n14145, ZN => n1243);
   U1112 : OAI22_X1 port map( A1 => n16000, A2 => n14146, B1 => n14187, B2 => 
                           n14145, ZN => n1242);
   U1113 : OAI22_X1 port map( A1 => n16756, A2 => n14146, B1 => n14188, B2 => 
                           n14145, ZN => n1241);
   U1114 : OAI22_X1 port map( A1 => n16757, A2 => n14146, B1 => n14189, B2 => 
                           n14145, ZN => n1240);
   U1115 : OAI22_X1 port map( A1 => n16758, A2 => n14146, B1 => n14191, B2 => 
                           n14145, ZN => n1239);
   U1116 : NAND2_X1 port map( A1 => n14147, A2 => n14156, ZN => n14148);
   U1117 : CLKBUF_X1 port map( A => n14148, Z => n14149);
   U1118 : OAI22_X1 port map( A1 => n16031, A2 => n14150, B1 => n14158, B2 => 
                           n14149, ZN => n1238);
   U1119 : OAI22_X1 port map( A1 => n16491, A2 => n14150, B1 => n14159, B2 => 
                           n14148, ZN => n1237);
   U1120 : OAI22_X1 port map( A1 => n16759, A2 => n14150, B1 => n14160, B2 => 
                           n14149, ZN => n1236);
   U1121 : OAI22_X1 port map( A1 => n16492, A2 => n14150, B1 => n14161, B2 => 
                           n14148, ZN => n1235);
   U1122 : OAI22_X1 port map( A1 => n16493, A2 => n14150, B1 => n14162, B2 => 
                           n14149, ZN => n1234);
   U1123 : OAI22_X1 port map( A1 => n16760, A2 => n14150, B1 => n14163, B2 => 
                           n14148, ZN => n1233);
   U1124 : OAI22_X1 port map( A1 => n16001, A2 => n14150, B1 => n14164, B2 => 
                           n14149, ZN => n1232);
   U1125 : OAI22_X1 port map( A1 => n16494, A2 => n14150, B1 => n14165, B2 => 
                           n14148, ZN => n1231);
   U1126 : OAI22_X1 port map( A1 => n16761, A2 => n14150, B1 => n14166, B2 => 
                           n14149, ZN => n1230);
   U1127 : OAI22_X1 port map( A1 => n16762, A2 => n14150, B1 => n14167, B2 => 
                           n14148, ZN => n1229);
   U1128 : OAI22_X1 port map( A1 => n16495, A2 => n14150, B1 => n14168, B2 => 
                           n14148, ZN => n1228);
   U1129 : OAI22_X1 port map( A1 => n16763, A2 => n14150, B1 => n14169, B2 => 
                           n14149, ZN => n1227);
   U1130 : OAI22_X1 port map( A1 => n16496, A2 => n14150, B1 => n14170, B2 => 
                           n14148, ZN => n1226);
   U1131 : OAI22_X1 port map( A1 => n16497, A2 => n14150, B1 => n14171, B2 => 
                           n14149, ZN => n1225);
   U1132 : OAI22_X1 port map( A1 => n16498, A2 => n14150, B1 => n14172, B2 => 
                           n14148, ZN => n1224);
   U1133 : OAI22_X1 port map( A1 => n16764, A2 => n14150, B1 => n14173, B2 => 
                           n14149, ZN => n1223);
   U1134 : OAI22_X1 port map( A1 => n16765, A2 => n14150, B1 => n14174, B2 => 
                           n14148, ZN => n1222);
   U1135 : OAI22_X1 port map( A1 => n16002, A2 => n14150, B1 => n14175, B2 => 
                           n14148, ZN => n1221);
   U1136 : OAI22_X1 port map( A1 => n16499, A2 => n14150, B1 => n14176, B2 => 
                           n14148, ZN => n1220);
   U1137 : OAI22_X1 port map( A1 => n16766, A2 => n14150, B1 => n14177, B2 => 
                           n14148, ZN => n1219);
   U1138 : OAI22_X1 port map( A1 => n16767, A2 => n14150, B1 => n14178, B2 => 
                           n14148, ZN => n1218);
   U1139 : OAI22_X1 port map( A1 => n16500, A2 => n14150, B1 => n14179, B2 => 
                           n14148, ZN => n1217);
   U1140 : OAI22_X1 port map( A1 => n16501, A2 => n14150, B1 => n14181, B2 => 
                           n14148, ZN => n1216);
   U1141 : OAI22_X1 port map( A1 => n16768, A2 => n14150, B1 => n14182, B2 => 
                           n14149, ZN => n1215);
   U1142 : OAI22_X1 port map( A1 => n16502, A2 => n14150, B1 => n14183, B2 => 
                           n14149, ZN => n1214);
   U1143 : OAI22_X1 port map( A1 => n16769, A2 => n14150, B1 => n14184, B2 => 
                           n14149, ZN => n1213);
   U1144 : OAI22_X1 port map( A1 => n16503, A2 => n14150, B1 => n14185, B2 => 
                           n14149, ZN => n1212);
   U1145 : OAI22_X1 port map( A1 => n16770, A2 => n14150, B1 => n14186, B2 => 
                           n14149, ZN => n1211);
   U1146 : OAI22_X1 port map( A1 => n16504, A2 => n14150, B1 => n14187, B2 => 
                           n14149, ZN => n1210);
   U1147 : OAI22_X1 port map( A1 => n16505, A2 => n14150, B1 => n14188, B2 => 
                           n14149, ZN => n1209);
   U1148 : OAI22_X1 port map( A1 => n16506, A2 => n14150, B1 => n14189, B2 => 
                           n14149, ZN => n1208);
   U1149 : OAI22_X1 port map( A1 => n16248, A2 => n14150, B1 => n14191, B2 => 
                           n14149, ZN => n1207);
   U1150 : NAND2_X1 port map( A1 => n14151, A2 => n14156, ZN => n14152);
   U1151 : CLKBUF_X1 port map( A => n14155, Z => n14153);
   U1152 : CLKBUF_X1 port map( A => n14152, Z => n14154);
   U1153 : OAI22_X1 port map( A1 => n15760, A2 => n14153, B1 => n14158, B2 => 
                           n14154, ZN => n1206);
   U1154 : OAI22_X1 port map( A1 => n16249, A2 => n14155, B1 => n14159, B2 => 
                           n14152, ZN => n1205);
   U1155 : OAI22_X1 port map( A1 => n16003, A2 => n14153, B1 => n14160, B2 => 
                           n14154, ZN => n1204);
   U1156 : OAI22_X1 port map( A1 => n16250, A2 => n14155, B1 => n14161, B2 => 
                           n14152, ZN => n1203);
   U1157 : OAI22_X1 port map( A1 => n16251, A2 => n14153, B1 => n14162, B2 => 
                           n14154, ZN => n1202);
   U1158 : OAI22_X1 port map( A1 => n16252, A2 => n14155, B1 => n14163, B2 => 
                           n14152, ZN => n1201);
   U1159 : OAI22_X1 port map( A1 => n16253, A2 => n14153, B1 => n14164, B2 => 
                           n14154, ZN => n1200);
   U1160 : OAI22_X1 port map( A1 => n16004, A2 => n14155, B1 => n14165, B2 => 
                           n14152, ZN => n1199);
   U1161 : OAI22_X1 port map( A1 => n16005, A2 => n14153, B1 => n14166, B2 => 
                           n14154, ZN => n1198);
   U1162 : OAI22_X1 port map( A1 => n16006, A2 => n14155, B1 => n14167, B2 => 
                           n14152, ZN => n1197);
   U1163 : OAI22_X1 port map( A1 => n16254, A2 => n14155, B1 => n14168, B2 => 
                           n14152, ZN => n1196);
   U1164 : OAI22_X1 port map( A1 => n16007, A2 => n14155, B1 => n14169, B2 => 
                           n14154, ZN => n1195);
   U1165 : OAI22_X1 port map( A1 => n16008, A2 => n14153, B1 => n14170, B2 => 
                           n14152, ZN => n1194);
   U1166 : OAI22_X1 port map( A1 => n16255, A2 => n14153, B1 => n14171, B2 => 
                           n14154, ZN => n1193);
   U1167 : OAI22_X1 port map( A1 => n16009, A2 => n14153, B1 => n14172, B2 => 
                           n14152, ZN => n1192);
   U1168 : OAI22_X1 port map( A1 => n16256, A2 => n14153, B1 => n14173, B2 => 
                           n14154, ZN => n1191);
   U1169 : OAI22_X1 port map( A1 => n16010, A2 => n14153, B1 => n14174, B2 => 
                           n14152, ZN => n1190);
   U1170 : OAI22_X1 port map( A1 => n16257, A2 => n14153, B1 => n14175, B2 => 
                           n14152, ZN => n1189);
   U1171 : OAI22_X1 port map( A1 => n16011, A2 => n14153, B1 => n14176, B2 => 
                           n14152, ZN => n1188);
   U1172 : OAI22_X1 port map( A1 => n16012, A2 => n14153, B1 => n14177, B2 => 
                           n14152, ZN => n1187);
   U1173 : OAI22_X1 port map( A1 => n16013, A2 => n14153, B1 => n14178, B2 => 
                           n14152, ZN => n1186);
   U1174 : OAI22_X1 port map( A1 => n16258, A2 => n14153, B1 => n14179, B2 => 
                           n14152, ZN => n1185);
   U1175 : OAI22_X1 port map( A1 => n16014, A2 => n14153, B1 => n14181, B2 => 
                           n14152, ZN => n1184);
   U1176 : OAI22_X1 port map( A1 => n16015, A2 => n14153, B1 => n14182, B2 => 
                           n14154, ZN => n1183);
   U1177 : OAI22_X1 port map( A1 => n16259, A2 => n14155, B1 => n14183, B2 => 
                           n14154, ZN => n1182);
   U1178 : OAI22_X1 port map( A1 => n16260, A2 => n14155, B1 => n14184, B2 => 
                           n14154, ZN => n1181);
   U1179 : OAI22_X1 port map( A1 => n16016, A2 => n14155, B1 => n14185, B2 => 
                           n14154, ZN => n1180);
   U1180 : OAI22_X1 port map( A1 => n16017, A2 => n14155, B1 => n14186, B2 => 
                           n14154, ZN => n1179);
   U1181 : OAI22_X1 port map( A1 => n16018, A2 => n14155, B1 => n14187, B2 => 
                           n14154, ZN => n1178);
   U1182 : OAI22_X1 port map( A1 => n16261, A2 => n14155, B1 => n14188, B2 => 
                           n14154, ZN => n1177);
   U1183 : OAI22_X1 port map( A1 => n16262, A2 => n14155, B1 => n14189, B2 => 
                           n14154, ZN => n1176);
   U1184 : OAI22_X1 port map( A1 => n16019, A2 => n14155, B1 => n14191, B2 => 
                           n14154, ZN => n1175);
   U1185 : NAND2_X1 port map( A1 => n14157, A2 => n14156, ZN => n14180);
   U1186 : CLKBUF_X1 port map( A => n14180, Z => n14190);
   U1187 : OAI22_X1 port map( A1 => n16275, A2 => n14192, B1 => n14158, B2 => 
                           n14190, ZN => n1174);
   U1188 : OAI22_X1 port map( A1 => n16771, A2 => n14192, B1 => n14159, B2 => 
                           n14180, ZN => n1173);
   U1189 : OAI22_X1 port map( A1 => n16263, A2 => n14192, B1 => n14160, B2 => 
                           n14190, ZN => n1172);
   U1190 : OAI22_X1 port map( A1 => n16020, A2 => n14192, B1 => n14161, B2 => 
                           n14180, ZN => n1171);
   U1191 : OAI22_X1 port map( A1 => n16507, A2 => n14192, B1 => n14162, B2 => 
                           n14190, ZN => n1170);
   U1192 : OAI22_X1 port map( A1 => n16508, A2 => n14192, B1 => n14163, B2 => 
                           n14180, ZN => n1169);
   U1193 : OAI22_X1 port map( A1 => n16772, A2 => n14192, B1 => n14164, B2 => 
                           n14190, ZN => n1168);
   U1194 : OAI22_X1 port map( A1 => n16773, A2 => n14192, B1 => n14165, B2 => 
                           n14180, ZN => n1167);
   U1195 : OAI22_X1 port map( A1 => n16509, A2 => n14192, B1 => n14166, B2 => 
                           n14190, ZN => n1166);
   U1196 : OAI22_X1 port map( A1 => n16264, A2 => n14192, B1 => n14167, B2 => 
                           n14180, ZN => n1165);
   U1197 : OAI22_X1 port map( A1 => n16021, A2 => n14192, B1 => n14168, B2 => 
                           n14180, ZN => n1164);
   U1198 : OAI22_X1 port map( A1 => n16022, A2 => n14192, B1 => n14169, B2 => 
                           n14190, ZN => n1163);
   U1199 : OAI22_X1 port map( A1 => n16510, A2 => n14192, B1 => n14170, B2 => 
                           n14180, ZN => n1162);
   U1200 : OAI22_X1 port map( A1 => n16774, A2 => n14192, B1 => n14171, B2 => 
                           n14190, ZN => n1161);
   U1201 : OAI22_X1 port map( A1 => n16265, A2 => n14192, B1 => n14172, B2 => 
                           n14180, ZN => n1160);
   U1202 : OAI22_X1 port map( A1 => n16023, A2 => n14192, B1 => n14173, B2 => 
                           n14190, ZN => n1159);
   U1203 : OAI22_X1 port map( A1 => n16775, A2 => n14192, B1 => n14174, B2 => 
                           n14180, ZN => n1158);
   U1204 : OAI22_X1 port map( A1 => n16776, A2 => n14192, B1 => n14175, B2 => 
                           n14180, ZN => n1157);
   U1205 : OAI22_X1 port map( A1 => n16024, A2 => n14192, B1 => n14176, B2 => 
                           n14180, ZN => n1156);
   U1206 : OAI22_X1 port map( A1 => n16266, A2 => n14192, B1 => n14177, B2 => 
                           n14180, ZN => n1155);
   U1207 : OAI22_X1 port map( A1 => n16267, A2 => n14192, B1 => n14178, B2 => 
                           n14180, ZN => n1154);
   U1208 : OAI22_X1 port map( A1 => n16268, A2 => n14192, B1 => n14179, B2 => 
                           n14180, ZN => n1153);
   U1209 : OAI22_X1 port map( A1 => n16269, A2 => n14192, B1 => n14181, B2 => 
                           n14180, ZN => n1152);
   U1210 : OAI22_X1 port map( A1 => n16511, A2 => n14192, B1 => n14182, B2 => 
                           n14190, ZN => n1151);
   U1211 : OAI22_X1 port map( A1 => n16512, A2 => n14192, B1 => n14183, B2 => 
                           n14190, ZN => n1150);
   U1212 : OAI22_X1 port map( A1 => n16270, A2 => n14192, B1 => n14184, B2 => 
                           n14190, ZN => n1149);
   U1213 : OAI22_X1 port map( A1 => n16777, A2 => n14192, B1 => n14185, B2 => 
                           n14190, ZN => n1148);
   U1214 : OAI22_X1 port map( A1 => n16513, A2 => n14192, B1 => n14186, B2 => 
                           n14190, ZN => n1147);
   U1215 : OAI22_X1 port map( A1 => n16778, A2 => n14192, B1 => n14187, B2 => 
                           n14190, ZN => n1146);
   U1216 : OAI22_X1 port map( A1 => n16779, A2 => n14192, B1 => n14188, B2 => 
                           n14190, ZN => n1145);
   U1217 : OAI22_X1 port map( A1 => n16025, A2 => n14192, B1 => n14189, B2 => 
                           n14190, ZN => n1144);
   U1218 : OAI22_X1 port map( A1 => n16514, A2 => n14192, B1 => n14191, B2 => 
                           n14190, ZN => n1143);
   U1219 : NAND3_X1 port map( A1 => n14003, A2 => ENABLE, A3 => RD2, ZN => 
                           n14973);
   U1220 : INV_X1 port map( A => ADD_RD2(3), ZN => n14218);
   U1221 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n14218, ZN => n14201);
   U1222 : INV_X1 port map( A => ADD_RD2(2), ZN => n14194);
   U1223 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n14194,
                           ZN => n14210);
   U1224 : NOR2_X1 port map( A1 => n14201, A2 => n14210, ZN => n14697);
   U1225 : INV_X1 port map( A => ADD_RD2(1), ZN => n14193);
   U1226 : OR3_X1 port map( A1 => n14193, A2 => ADD_RD2(2), A3 => ADD_RD2(0), 
                           ZN => n14237);
   U1227 : NOR2_X1 port map( A1 => n14201, A2 => n14237, ZN => n14653);
   U1228 : CLKBUF_X1 port map( A => n14653, Z => n14935);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n14697, B1 => 
                           REGISTERS_18_31_port, B2 => n14935, ZN => n14199);
   U1230 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n14200)
                           ;
   U1231 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n14194, A3 => n14193, ZN 
                           => n14211);
   U1232 : NOR2_X1 port map( A1 => n14200, A2 => n14211, ZN => n14928);
   U1233 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n14193,
                           ZN => n14212);
   U1234 : NOR2_X1 port map( A1 => n14201, A2 => n14212, ZN => n14608);
   U1235 : CLKBUF_X1 port map( A => n14608, Z => n14923);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n14928, B1 => 
                           REGISTERS_21_31_port, B2 => n14923, ZN => n14198);
   U1237 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), ZN => n14195);
   U1238 : NAND2_X1 port map( A1 => ADD_RD2(2), A2 => n14195, ZN => n14213);
   U1239 : NOR2_X1 port map( A1 => n14201, A2 => n14213, ZN => n14541);
   U1240 : OR3_X1 port map( A1 => n14194, A2 => n14193, A3 => ADD_RD2(0), ZN =>
                           n14242);
   U1241 : NOR2_X1 port map( A1 => n14200, A2 => n14242, ZN => n14921);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n14541, B1 => 
                           REGISTERS_30_31_port, B2 => n14921, ZN => n14197);
   U1243 : NAND2_X1 port map( A1 => n14195, A2 => n14194, ZN => n14209);
   U1244 : NOR2_X1 port map( A1 => n14201, A2 => n14209, ZN => n14702);
   U1245 : NOR2_X1 port map( A1 => n14200, A2 => n14209, ZN => n14839);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n14702, B1 => 
                           REGISTERS_24_31_port, B2 => n14839, ZN => n14196);
   U1247 : NAND4_X1 port map( A1 => n14199, A2 => n14198, A3 => n14197, A4 => 
                           n14196, ZN => n14207);
   U1248 : NOR2_X1 port map( A1 => n14201, A2 => n14242, ZN => n14678);
   U1249 : NOR2_X1 port map( A1 => n14200, A2 => n14210, ZN => n14820);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n14678, B1 => 
                           REGISTERS_27_31_port, B2 => n14820, ZN => n14205);
   U1251 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => 
                           ADD_RD2(1), ZN => n14208);
   U1252 : NOR2_X1 port map( A1 => n14201, A2 => n14208, ZN => n14940);
   U1253 : NOR2_X1 port map( A1 => n14200, A2 => n14212, ZN => n14939);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n14940, B1 => 
                           REGISTERS_29_31_port, B2 => n14939, ZN => n14204);
   U1255 : NOR2_X1 port map( A1 => n14208, A2 => n14200, ZN => n14893);
   U1256 : NOR2_X1 port map( A1 => n14200, A2 => n14237, ZN => n14891);
   U1257 : CLKBUF_X1 port map( A => n14891, Z => n14922);
   U1258 : AOI22_X1 port map( A1 => REGISTERS_31_31_port, A2 => n14893, B1 => 
                           REGISTERS_26_31_port, B2 => n14922, ZN => n14203);
   U1259 : NOR2_X1 port map( A1 => n14200, A2 => n14213, ZN => n14840);
   U1260 : NOR2_X1 port map( A1 => n14201, A2 => n14211, ZN => n14846);
   U1261 : CLKBUF_X1 port map( A => n14846, Z => n14924);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n14840, B1 => 
                           REGISTERS_17_31_port, B2 => n14924, ZN => n14202);
   U1263 : NAND4_X1 port map( A1 => n14205, A2 => n14204, A3 => n14203, A4 => 
                           n14202, ZN => n14206);
   U1264 : NOR2_X1 port map( A1 => n14207, A2 => n14206, ZN => n14226);
   U1265 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n14920, 
                           ZN => n14970);
   U1266 : CLKBUF_X1 port map( A => n14970, Z => n14788);
   U1267 : INV_X1 port map( A => n14242, ZN => n14882);
   U1268 : INV_X1 port map( A => n14237, ZN => n14958);
   U1269 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_6_31_port, B1 => 
                           n14958, B2 => REGISTERS_2_31_port, ZN => n14217);
   U1270 : INV_X1 port map( A => n14208, ZN => n14877);
   U1271 : CLKBUF_X1 port map( A => n14877, Z => n14664);
   U1272 : INV_X1 port map( A => n14209, ZN => n14876);
   U1273 : CLKBUF_X1 port map( A => n14876, Z => n14665);
   U1274 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_31_port, B1 => 
                           n14665, B2 => REGISTERS_0_31_port, ZN => n14216);
   U1275 : INV_X1 port map( A => n14210, ZN => n14801);
   U1276 : CLKBUF_X1 port map( A => n14801, Z => n14911);
   U1277 : INV_X1 port map( A => n14211, ZN => n14909);
   U1278 : CLKBUF_X1 port map( A => n14909, Z => n14948);
   U1279 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_31_port, B1 => 
                           n14948, B2 => REGISTERS_1_31_port, ZN => n14215);
   U1280 : INV_X1 port map( A => n14212, ZN => n14733);
   U1281 : INV_X1 port map( A => n14213, ZN => n14910);
   U1282 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_31_port, B1 => 
                           n14910, B2 => REGISTERS_4_31_port, ZN => n14214);
   U1283 : NAND4_X1 port map( A1 => n14217, A2 => n14216, A3 => n14215, A4 => 
                           n14214, ZN => n14224);
   U1284 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n14218, A3 => n14920, ZN 
                           => n14968);
   U1285 : CLKBUF_X1 port map( A => n14968, Z => n14811);
   U1286 : CLKBUF_X1 port map( A => n14910, Z => n14853);
   U1287 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_11_31_port, B1 => 
                           n14853, B2 => REGISTERS_12_31_port, ZN => n14222);
   U1288 : INV_X1 port map( A => n14237, ZN => n14904);
   U1289 : AOI22_X1 port map( A1 => n14904, A2 => REGISTERS_10_31_port, B1 => 
                           n14665, B2 => REGISTERS_8_31_port, ZN => n14221);
   U1290 : CLKBUF_X1 port map( A => n14733, Z => n14961);
   U1291 : INV_X1 port map( A => n14242, ZN => n14949);
   U1292 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_13_31_port, B1 => 
                           n14949, B2 => REGISTERS_14_31_port, ZN => n14220);
   U1293 : CLKBUF_X1 port map( A => n14909, Z => n14959);
   U1294 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_31_port, B1 => 
                           n14959, B2 => REGISTERS_9_31_port, ZN => n14219);
   U1295 : NAND4_X1 port map( A1 => n14222, A2 => n14221, A3 => n14220, A4 => 
                           n14219, ZN => n14223);
   U1296 : AOI22_X1 port map( A1 => n14788, A2 => n14224, B1 => n14811, B2 => 
                           n14223, ZN => n14225);
   U1297 : OAI21_X1 port map( B1 => n14920, B2 => n14226, A => n14225, ZN => 
                           N448);
   U1298 : CLKBUF_X1 port map( A => n14940, Z => n14721);
   U1299 : CLKBUF_X1 port map( A => n14541, Z => n14933);
   U1300 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_30_port, B1 => 
                           n14933, B2 => REGISTERS_20_30_port, ZN => n14230);
   U1301 : CLKBUF_X1 port map( A => n14928, Z => n14845);
   U1302 : CLKBUF_X1 port map( A => n14839, Z => n14937);
   U1303 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_30_port, B1 => 
                           n14937, B2 => REGISTERS_24_30_port, ZN => n14229);
   U1304 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_30_port, B1 => 
                           n14678, B2 => REGISTERS_22_30_port, ZN => n14228);
   U1305 : CLKBUF_X1 port map( A => n14702, Z => n14927);
   U1306 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_30_port, B1 => 
                           n14927, B2 => REGISTERS_16_30_port, ZN => n14227);
   U1307 : NAND4_X1 port map( A1 => n14230, A2 => n14229, A3 => n14228, A4 => 
                           n14227, ZN => n14236);
   U1308 : CLKBUF_X1 port map( A => n14840, Z => n14934);
   U1309 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_30_port, B1 => 
                           n14923, B2 => REGISTERS_21_30_port, ZN => n14234);
   U1310 : CLKBUF_X1 port map( A => n14893, Z => n14926);
   U1311 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_30_port, B1 => 
                           n14935, B2 => REGISTERS_18_30_port, ZN => n14233);
   U1312 : CLKBUF_X1 port map( A => n14697, Z => n14925);
   U1313 : CLKBUF_X1 port map( A => n14921, Z => n14726);
   U1314 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_30_port, B1 => 
                           n14726, B2 => REGISTERS_30_30_port, ZN => n14232);
   U1315 : AOI22_X1 port map( A1 => n14820, A2 => REGISTERS_27_30_port, B1 => 
                           n14846, B2 => REGISTERS_17_30_port, ZN => n14231);
   U1316 : NAND4_X1 port map( A1 => n14234, A2 => n14233, A3 => n14232, A4 => 
                           n14231, ZN => n14235);
   U1317 : NOR2_X1 port map( A1 => n14236, A2 => n14235, ZN => n14250);
   U1318 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_3_30_port, B1 => 
                           n14959, B2 => REGISTERS_1_30_port, ZN => n14241);
   U1319 : CLKBUF_X1 port map( A => n14910, Z => n14955);
   U1320 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_30_port, B1 => 
                           n14665, B2 => REGISTERS_0_30_port, ZN => n14240);
   U1321 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_30_port, B1 => 
                           n14949, B2 => REGISTERS_6_30_port, ZN => n14239);
   U1322 : INV_X1 port map( A => n14237, ZN => n14947);
   U1323 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_30_port, B1 => 
                           n14947, B2 => REGISTERS_2_30_port, ZN => n14238);
   U1324 : NAND4_X1 port map( A1 => n14241, A2 => n14240, A3 => n14239, A4 => 
                           n14238, ZN => n14248);
   U1325 : INV_X1 port map( A => n14242, ZN => n14960);
   U1326 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_30_port, B1 => 
                           n14959, B2 => REGISTERS_9_30_port, ZN => n14246);
   U1327 : CLKBUF_X1 port map( A => n14801, Z => n14956);
   U1328 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_30_port, B1 => 
                           n14956, B2 => REGISTERS_11_30_port, ZN => n14245);
   U1329 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_30_port, B1 => 
                           n14665, B2 => REGISTERS_8_30_port, ZN => n14244);
   U1330 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_30_port, B1 => 
                           n14947, B2 => REGISTERS_10_30_port, ZN => n14243);
   U1331 : NAND4_X1 port map( A1 => n14246, A2 => n14245, A3 => n14244, A4 => 
                           n14243, ZN => n14247);
   U1332 : AOI22_X1 port map( A1 => n14788, A2 => n14248, B1 => n14811, B2 => 
                           n14247, ZN => n14249);
   U1333 : OAI21_X1 port map( B1 => n14920, B2 => n14250, A => n14249, ZN => 
                           N447);
   U1334 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_29_port, B1 => 
                           n14726, B2 => REGISTERS_30_29_port, ZN => n14254);
   U1335 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_29_port, B1 => 
                           n14608, B2 => REGISTERS_21_29_port, ZN => n14253);
   U1336 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_29_port, B1 => 
                           n14839, B2 => REGISTERS_24_29_port, ZN => n14252);
   U1337 : AOI22_X1 port map( A1 => n14678, A2 => REGISTERS_22_29_port, B1 => 
                           n14893, B2 => REGISTERS_31_29_port, ZN => n14251);
   U1338 : NAND4_X1 port map( A1 => n14254, A2 => n14253, A3 => n14252, A4 => 
                           n14251, ZN => n14260);
   U1339 : AOI22_X1 port map( A1 => n14820, A2 => REGISTERS_27_29_port, B1 => 
                           n14846, B2 => REGISTERS_17_29_port, ZN => n14258);
   U1340 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_29_port, B1 => 
                           n14541, B2 => REGISTERS_20_29_port, ZN => n14257);
   U1341 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_29_port, B1 => 
                           n14702, B2 => REGISTERS_16_29_port, ZN => n14256);
   U1342 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_29_port, B1 => 
                           n14653, B2 => REGISTERS_18_29_port, ZN => n14255);
   U1343 : NAND4_X1 port map( A1 => n14258, A2 => n14257, A3 => n14256, A4 => 
                           n14255, ZN => n14259);
   U1344 : NOR2_X1 port map( A1 => n14260, A2 => n14259, ZN => n14272);
   U1345 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_29_port, B1 => 
                           n14947, B2 => REGISTERS_2_29_port, ZN => n14264);
   U1346 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_29_port, B1 => 
                           n14665, B2 => REGISTERS_0_29_port, ZN => n14263);
   U1347 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_29_port, B1 => 
                           n14853, B2 => REGISTERS_4_29_port, ZN => n14262);
   U1348 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_3_29_port, B1 => 
                           n14959, B2 => REGISTERS_1_29_port, ZN => n14261);
   U1349 : NAND4_X1 port map( A1 => n14264, A2 => n14263, A3 => n14262, A4 => 
                           n14261, ZN => n14270);
   U1350 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_29_port, B1 => 
                           n14665, B2 => REGISTERS_8_29_port, ZN => n14268);
   U1351 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_29_port, B1 => 
                           n14947, B2 => REGISTERS_10_29_port, ZN => n14267);
   U1352 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_11_29_port, B1 => 
                           n14853, B2 => REGISTERS_12_29_port, ZN => n14266);
   U1353 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_29_port, B1 => 
                           n14959, B2 => REGISTERS_9_29_port, ZN => n14265);
   U1354 : NAND4_X1 port map( A1 => n14268, A2 => n14267, A3 => n14266, A4 => 
                           n14265, ZN => n14269);
   U1355 : AOI22_X1 port map( A1 => n14788, A2 => n14270, B1 => n14811, B2 => 
                           n14269, ZN => n14271);
   U1356 : OAI21_X1 port map( B1 => n14920, B2 => n14272, A => n14271, ZN => 
                           N446);
   U1357 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_28_port, B1 => 
                           n14839, B2 => REGISTERS_24_28_port, ZN => n14276);
   U1358 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_28_port, B1 => 
                           n14608, B2 => REGISTERS_21_28_port, ZN => n14275);
   U1359 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_28_port, B1 => 
                           n14702, B2 => REGISTERS_16_28_port, ZN => n14274);
   U1360 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_28_port, B1 => 
                           n14893, B2 => REGISTERS_31_28_port, ZN => n14273);
   U1361 : NAND4_X1 port map( A1 => n14276, A2 => n14275, A3 => n14274, A4 => 
                           n14273, ZN => n14282);
   U1362 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_28_port, B1 => 
                           n14726, B2 => REGISTERS_30_28_port, ZN => n14280);
   U1363 : CLKBUF_X1 port map( A => n14678, Z => n14936);
   U1364 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_28_port, B1 => 
                           n14925, B2 => REGISTERS_19_28_port, ZN => n14279);
   U1365 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_28_port, B1 => 
                           n14653, B2 => REGISTERS_18_28_port, ZN => n14278);
   U1366 : AOI22_X1 port map( A1 => n14820, A2 => REGISTERS_27_28_port, B1 => 
                           n14541, B2 => REGISTERS_20_28_port, ZN => n14277);
   U1367 : NAND4_X1 port map( A1 => n14280, A2 => n14279, A3 => n14278, A4 => 
                           n14277, ZN => n14281);
   U1368 : NOR2_X1 port map( A1 => n14282, A2 => n14281, ZN => n14294);
   U1369 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_28_port, B1 => 
                           n14853, B2 => REGISTERS_4_28_port, ZN => n14286);
   U1370 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_28_port, B1 => 
                           n14909, B2 => REGISTERS_1_28_port, ZN => n14285);
   U1371 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_28_port, B1 => 
                           n14801, B2 => REGISTERS_3_28_port, ZN => n14284);
   U1372 : AOI22_X1 port map( A1 => n14958, A2 => REGISTERS_2_28_port, B1 => 
                           n14665, B2 => REGISTERS_0_28_port, ZN => n14283);
   U1373 : NAND4_X1 port map( A1 => n14286, A2 => n14285, A3 => n14284, A4 => 
                           n14283, ZN => n14292);
   U1374 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_28_port, B1 => 
                           n14801, B2 => REGISTERS_11_28_port, ZN => n14290);
   U1375 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_28_port, B1 => 
                           n14949, B2 => REGISTERS_14_28_port, ZN => n14289);
   U1376 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_28_port, B1 => 
                           n14959, B2 => REGISTERS_9_28_port, ZN => n14288);
   U1377 : AOI22_X1 port map( A1 => n14958, A2 => REGISTERS_10_28_port, B1 => 
                           n14665, B2 => REGISTERS_8_28_port, ZN => n14287);
   U1378 : NAND4_X1 port map( A1 => n14290, A2 => n14289, A3 => n14288, A4 => 
                           n14287, ZN => n14291);
   U1379 : AOI22_X1 port map( A1 => n14788, A2 => n14292, B1 => n14811, B2 => 
                           n14291, ZN => n14293);
   U1380 : OAI21_X1 port map( B1 => n14920, B2 => n14294, A => n14293, ZN => 
                           N445);
   U1381 : CLKBUF_X1 port map( A => n14820, Z => n14938);
   U1382 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_27_port, B1 => 
                           n14924, B2 => REGISTERS_17_27_port, ZN => n14298);
   U1383 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_27_port, B1 => 
                           n14608, B2 => REGISTERS_21_27_port, ZN => n14297);
   U1384 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_27_port, B1 => 
                           n14678, B2 => REGISTERS_22_27_port, ZN => n14296);
   U1385 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_27_port, B1 => 
                           n14541, B2 => REGISTERS_20_27_port, ZN => n14295);
   U1386 : NAND4_X1 port map( A1 => n14298, A2 => n14297, A3 => n14296, A4 => 
                           n14295, ZN => n14304);
   U1387 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_27_port, B1 => 
                           n14726, B2 => REGISTERS_30_27_port, ZN => n14302);
   U1388 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_27_port, B1 => 
                           n14839, B2 => REGISTERS_24_27_port, ZN => n14301);
   U1389 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_27_port, B1 => 
                           n14702, B2 => REGISTERS_16_27_port, ZN => n14300);
   U1390 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_27_port, B1 => 
                           n14653, B2 => REGISTERS_18_27_port, ZN => n14299);
   U1391 : NAND4_X1 port map( A1 => n14302, A2 => n14301, A3 => n14300, A4 => 
                           n14299, ZN => n14303);
   U1392 : NOR2_X1 port map( A1 => n14304, A2 => n14303, ZN => n14316);
   U1393 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_27_port, B1 => 
                           n14958, B2 => REGISTERS_2_27_port, ZN => n14308);
   U1394 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_27_port, B1 => 
                           n14665, B2 => REGISTERS_0_27_port, ZN => n14307);
   U1395 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_27_port, B1 => 
                           n14882, B2 => REGISTERS_6_27_port, ZN => n14306);
   U1396 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_3_27_port, B1 => 
                           n14853, B2 => REGISTERS_4_27_port, ZN => n14305);
   U1397 : NAND4_X1 port map( A1 => n14308, A2 => n14307, A3 => n14306, A4 => 
                           n14305, ZN => n14314);
   U1398 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_27_port, B1 => 
                           n14958, B2 => REGISTERS_10_27_port, ZN => n14312);
   U1399 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_27_port, B1 => 
                           n14882, B2 => REGISTERS_14_27_port, ZN => n14311);
   U1400 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_11_27_port, B1 => 
                           n14665, B2 => REGISTERS_8_27_port, ZN => n14310);
   U1401 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_27_port, B1 => 
                           n14909, B2 => REGISTERS_9_27_port, ZN => n14309);
   U1402 : NAND4_X1 port map( A1 => n14312, A2 => n14311, A3 => n14310, A4 => 
                           n14309, ZN => n14313);
   U1403 : AOI22_X1 port map( A1 => n14788, A2 => n14314, B1 => n14811, B2 => 
                           n14313, ZN => n14315);
   U1404 : OAI21_X1 port map( B1 => n14920, B2 => n14316, A => n14315, ZN => 
                           N444);
   U1405 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_26_port, B1 => 
                           n14924, B2 => REGISTERS_17_26_port, ZN => n14320);
   U1406 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_26_port, B1 => 
                           n14839, B2 => REGISTERS_24_26_port, ZN => n14319);
   U1407 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_26_port, B1 => 
                           n14541, B2 => REGISTERS_20_26_port, ZN => n14318);
   U1408 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_26_port, B1 => 
                           n14697, B2 => REGISTERS_19_26_port, ZN => n14317);
   U1409 : NAND4_X1 port map( A1 => n14320, A2 => n14319, A3 => n14318, A4 => 
                           n14317, ZN => n14326);
   U1410 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_26_port, B1 => 
                           n14928, B2 => REGISTERS_25_26_port, ZN => n14324);
   U1411 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_26_port, B1 => 
                           n14702, B2 => REGISTERS_16_26_port, ZN => n14323);
   U1412 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_26_port, B1 => 
                           n14653, B2 => REGISTERS_18_26_port, ZN => n14322);
   U1413 : AOI22_X1 port map( A1 => n14820, A2 => REGISTERS_27_26_port, B1 => 
                           n14726, B2 => REGISTERS_30_26_port, ZN => n14321);
   U1414 : NAND4_X1 port map( A1 => n14324, A2 => n14323, A3 => n14322, A4 => 
                           n14321, ZN => n14325);
   U1415 : NOR2_X1 port map( A1 => n14326, A2 => n14325, ZN => n14338);
   U1416 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_26_port, B1 => 
                           n14882, B2 => REGISTERS_6_26_port, ZN => n14330);
   U1417 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_26_port, B1 => 
                           n14958, B2 => REGISTERS_2_26_port, ZN => n14329);
   U1418 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_26_port, B1 => 
                           n14910, B2 => REGISTERS_4_26_port, ZN => n14328);
   U1419 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_26_port, B1 => 
                           n14665, B2 => REGISTERS_0_26_port, ZN => n14327);
   U1420 : NAND4_X1 port map( A1 => n14330, A2 => n14329, A3 => n14328, A4 => 
                           n14327, ZN => n14336);
   U1421 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_26_port, B1 => 
                           n14665, B2 => REGISTERS_8_26_port, ZN => n14334);
   U1422 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_26_port, B1 => 
                           n14882, B2 => REGISTERS_14_26_port, ZN => n14333);
   U1423 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_13_26_port, B1 => 
                           n14853, B2 => REGISTERS_12_26_port, ZN => n14332);
   U1424 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_9_26_port, B1 => 
                           n14958, B2 => REGISTERS_10_26_port, ZN => n14331);
   U1425 : NAND4_X1 port map( A1 => n14334, A2 => n14333, A3 => n14332, A4 => 
                           n14331, ZN => n14335);
   U1426 : AOI22_X1 port map( A1 => n14788, A2 => n14336, B1 => n14811, B2 => 
                           n14335, ZN => n14337);
   U1427 : OAI21_X1 port map( B1 => n14920, B2 => n14338, A => n14337, ZN => 
                           N443);
   U1428 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_25_port, B1 => 
                           n14839, B2 => REGISTERS_24_25_port, ZN => n14342);
   U1429 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_25_port, B1 => 
                           n14653, B2 => REGISTERS_18_25_port, ZN => n14341);
   U1430 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_25_port, B1 => 
                           n14924, B2 => REGISTERS_17_25_port, ZN => n14340);
   U1431 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_25_port, B1 => 
                           n14541, B2 => REGISTERS_20_25_port, ZN => n14339);
   U1432 : NAND4_X1 port map( A1 => n14342, A2 => n14341, A3 => n14340, A4 => 
                           n14339, ZN => n14348);
   U1433 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_25_port, B1 => 
                           n14726, B2 => REGISTERS_30_25_port, ZN => n14346);
   U1434 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_25_port, B1 => 
                           n14702, B2 => REGISTERS_16_25_port, ZN => n14345);
   U1435 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_25_port, B1 => 
                           n14939, B2 => REGISTERS_29_25_port, ZN => n14344);
   U1436 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_25_port, B1 => 
                           n14928, B2 => REGISTERS_25_25_port, ZN => n14343);
   U1437 : NAND4_X1 port map( A1 => n14346, A2 => n14345, A3 => n14344, A4 => 
                           n14343, ZN => n14347);
   U1438 : NOR2_X1 port map( A1 => n14348, A2 => n14347, ZN => n14360);
   U1439 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_25_port, B1 => 
                           n14956, B2 => REGISTERS_3_25_port, ZN => n14352);
   U1440 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_25_port, B1 => 
                           n14959, B2 => REGISTERS_1_25_port, ZN => n14351);
   U1441 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_25_port, B1 => 
                           n14910, B2 => REGISTERS_4_25_port, ZN => n14350);
   U1442 : AOI22_X1 port map( A1 => n14947, A2 => REGISTERS_2_25_port, B1 => 
                           n14665, B2 => REGISTERS_0_25_port, ZN => n14349);
   U1443 : NAND4_X1 port map( A1 => n14352, A2 => n14351, A3 => n14350, A4 => 
                           n14349, ZN => n14358);
   U1444 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_25_port, B1 => 
                           n14909, B2 => REGISTERS_9_25_port, ZN => n14356);
   U1445 : CLKBUF_X1 port map( A => n14877, Z => n14962);
   U1446 : CLKBUF_X1 port map( A => n14876, Z => n14957);
   U1447 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_25_port, B1 => 
                           n14957, B2 => REGISTERS_8_25_port, ZN => n14355);
   U1448 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_25_port, B1 => 
                           n14958, B2 => REGISTERS_10_25_port, ZN => n14354);
   U1449 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_11_25_port, B1 => 
                           n14853, B2 => REGISTERS_12_25_port, ZN => n14353);
   U1450 : NAND4_X1 port map( A1 => n14356, A2 => n14355, A3 => n14354, A4 => 
                           n14353, ZN => n14357);
   U1451 : AOI22_X1 port map( A1 => n14788, A2 => n14358, B1 => n14811, B2 => 
                           n14357, ZN => n14359);
   U1452 : OAI21_X1 port map( B1 => n14920, B2 => n14360, A => n14359, ZN => 
                           N442);
   U1453 : CLKBUF_X1 port map( A => n14939, Z => n14892);
   U1454 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_24_port, B1 => 
                           n14678, B2 => REGISTERS_22_24_port, ZN => n14364);
   U1455 : AOI22_X1 port map( A1 => n14933, A2 => REGISTERS_20_24_port, B1 => 
                           n14726, B2 => REGISTERS_30_24_port, ZN => n14363);
   U1456 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_24_port, B1 => 
                           n14891, B2 => REGISTERS_26_24_port, ZN => n14362);
   U1457 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_24_port, B1 => 
                           n14608, B2 => REGISTERS_21_24_port, ZN => n14361);
   U1458 : NAND4_X1 port map( A1 => n14364, A2 => n14363, A3 => n14362, A4 => 
                           n14361, ZN => n14370);
   U1459 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_24_port, B1 => 
                           n14697, B2 => REGISTERS_19_24_port, ZN => n14368);
   U1460 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_24_port, B1 => 
                           n14845, B2 => REGISTERS_25_24_port, ZN => n14367);
   U1461 : AOI22_X1 port map( A1 => n14927, A2 => REGISTERS_16_24_port, B1 => 
                           n14839, B2 => REGISTERS_24_24_port, ZN => n14366);
   U1462 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_24_port, B1 => 
                           n14653, B2 => REGISTERS_18_24_port, ZN => n14365);
   U1463 : NAND4_X1 port map( A1 => n14368, A2 => n14367, A3 => n14366, A4 => 
                           n14365, ZN => n14369);
   U1464 : NOR2_X1 port map( A1 => n14370, A2 => n14369, ZN => n14382);
   U1465 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_24_port, B1 => 
                           n14956, B2 => REGISTERS_3_24_port, ZN => n14374);
   U1466 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_24_port, B1 => 
                           n14876, B2 => REGISTERS_0_24_port, ZN => n14373);
   U1467 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_24_port, B1 => 
                           n14958, B2 => REGISTERS_2_24_port, ZN => n14372);
   U1468 : CLKBUF_X1 port map( A => n14733, Z => n14950);
   U1469 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_24_port, B1 => 
                           n14959, B2 => REGISTERS_1_24_port, ZN => n14371);
   U1470 : NAND4_X1 port map( A1 => n14374, A2 => n14373, A3 => n14372, A4 => 
                           n14371, ZN => n14380);
   U1471 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_13_24_port, B1 => 
                           n14956, B2 => REGISTERS_11_24_port, ZN => n14378);
   U1472 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_24_port, B1 => 
                           n14958, B2 => REGISTERS_10_24_port, ZN => n14377);
   U1473 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_9_24_port, B1 => 
                           n14665, B2 => REGISTERS_8_24_port, ZN => n14376);
   U1474 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_24_port, B1 => 
                           n14910, B2 => REGISTERS_12_24_port, ZN => n14375);
   U1475 : NAND4_X1 port map( A1 => n14378, A2 => n14377, A3 => n14376, A4 => 
                           n14375, ZN => n14379);
   U1476 : AOI22_X1 port map( A1 => n14788, A2 => n14380, B1 => n14811, B2 => 
                           n14379, ZN => n14381);
   U1477 : OAI21_X1 port map( B1 => n14920, B2 => n14382, A => n14381, ZN => 
                           N441);
   U1478 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_23_port, B1 => 
                           n14653, B2 => REGISTERS_18_23_port, ZN => n14386);
   U1479 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_23_port, B1 => 
                           n14845, B2 => REGISTERS_25_23_port, ZN => n14385);
   U1480 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_23_port, B1 => 
                           n14726, B2 => REGISTERS_30_23_port, ZN => n14384);
   U1481 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_23_port, B1 => 
                           n14697, B2 => REGISTERS_19_23_port, ZN => n14383);
   U1482 : NAND4_X1 port map( A1 => n14386, A2 => n14385, A3 => n14384, A4 => 
                           n14383, ZN => n14392);
   U1483 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_23_port, B1 => 
                           n14541, B2 => REGISTERS_20_23_port, ZN => n14390);
   U1484 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_23_port, B1 => 
                           n14839, B2 => REGISTERS_24_23_port, ZN => n14389);
   U1485 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_23_port, B1 => 
                           n14702, B2 => REGISTERS_16_23_port, ZN => n14388);
   U1486 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_23_port, B1 => 
                           n14820, B2 => REGISTERS_27_23_port, ZN => n14387);
   U1487 : NAND4_X1 port map( A1 => n14390, A2 => n14389, A3 => n14388, A4 => 
                           n14387, ZN => n14391);
   U1488 : NOR2_X1 port map( A1 => n14392, A2 => n14391, ZN => n14404);
   U1489 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_23_port, B1 => 
                           n14853, B2 => REGISTERS_4_23_port, ZN => n14396);
   U1490 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_23_port, B1 => 
                           n14958, B2 => REGISTERS_2_23_port, ZN => n14395);
   U1491 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_23_port, B1 => 
                           n14956, B2 => REGISTERS_3_23_port, ZN => n14394);
   U1492 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_23_port, B1 => 
                           n14957, B2 => REGISTERS_0_23_port, ZN => n14393);
   U1493 : NAND4_X1 port map( A1 => n14396, A2 => n14395, A3 => n14394, A4 => 
                           n14393, ZN => n14402);
   U1494 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_23_port, B1 => 
                           n14911, B2 => REGISTERS_11_23_port, ZN => n14400);
   U1495 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_13_23_port, B1 => 
                           n14876, B2 => REGISTERS_8_23_port, ZN => n14399);
   U1496 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_23_port, B1 => 
                           n14958, B2 => REGISTERS_10_23_port, ZN => n14398);
   U1497 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_23_port, B1 => 
                           n14909, B2 => REGISTERS_9_23_port, ZN => n14397);
   U1498 : NAND4_X1 port map( A1 => n14400, A2 => n14399, A3 => n14398, A4 => 
                           n14397, ZN => n14401);
   U1499 : AOI22_X1 port map( A1 => n14788, A2 => n14402, B1 => n14811, B2 => 
                           n14401, ZN => n14403);
   U1500 : OAI21_X1 port map( B1 => n14973, B2 => n14404, A => n14403, ZN => 
                           N440);
   U1501 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_22_port, B1 => 
                           n14653, B2 => REGISTERS_18_22_port, ZN => n14408);
   U1502 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_22_port, B1 => 
                           n14702, B2 => REGISTERS_16_22_port, ZN => n14407);
   U1503 : AOI22_X1 port map( A1 => n14541, A2 => REGISTERS_20_22_port, B1 => 
                           n14726, B2 => REGISTERS_30_22_port, ZN => n14406);
   U1504 : AOI22_X1 port map( A1 => n14928, A2 => REGISTERS_25_22_port, B1 => 
                           n14608, B2 => REGISTERS_21_22_port, ZN => n14405);
   U1505 : NAND4_X1 port map( A1 => n14408, A2 => n14407, A3 => n14406, A4 => 
                           n14405, ZN => n14414);
   U1506 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_22_port, B1 => 
                           n14839, B2 => REGISTERS_24_22_port, ZN => n14412);
   U1507 : AOI22_X1 port map( A1 => n14939, A2 => REGISTERS_29_22_port, B1 => 
                           n14891, B2 => REGISTERS_26_22_port, ZN => n14411);
   U1508 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_22_port, B1 => 
                           n14840, B2 => REGISTERS_28_22_port, ZN => n14410);
   U1509 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_22_port, B1 => 
                           n14926, B2 => REGISTERS_31_22_port, ZN => n14409);
   U1510 : NAND4_X1 port map( A1 => n14412, A2 => n14411, A3 => n14410, A4 => 
                           n14409, ZN => n14413);
   U1511 : NOR2_X1 port map( A1 => n14414, A2 => n14413, ZN => n14426);
   U1512 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_22_port, B1 => 
                           n14665, B2 => REGISTERS_0_22_port, ZN => n14418);
   U1513 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_22_port, B1 => 
                           n14958, B2 => REGISTERS_2_22_port, ZN => n14417);
   U1514 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_22_port, B1 => 
                           n14956, B2 => REGISTERS_3_22_port, ZN => n14416);
   U1515 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_22_port, B1 => 
                           n14910, B2 => REGISTERS_4_22_port, ZN => n14415);
   U1516 : NAND4_X1 port map( A1 => n14418, A2 => n14417, A3 => n14416, A4 => 
                           n14415, ZN => n14424);
   U1517 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_11_22_port, B1 => 
                           n14959, B2 => REGISTERS_9_22_port, ZN => n14422);
   U1518 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_22_port, B1 => 
                           n14958, B2 => REGISTERS_10_22_port, ZN => n14421);
   U1519 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_22_port, B1 => 
                           n14960, B2 => REGISTERS_14_22_port, ZN => n14420);
   U1520 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_22_port, B1 => 
                           n14957, B2 => REGISTERS_8_22_port, ZN => n14419);
   U1521 : NAND4_X1 port map( A1 => n14422, A2 => n14421, A3 => n14420, A4 => 
                           n14419, ZN => n14423);
   U1522 : AOI22_X1 port map( A1 => n14788, A2 => n14424, B1 => n14811, B2 => 
                           n14423, ZN => n14425);
   U1523 : OAI21_X1 port map( B1 => n14973, B2 => n14426, A => n14425, ZN => 
                           N439);
   U1524 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_21_port, B1 => 
                           n14926, B2 => REGISTERS_31_21_port, ZN => n14430);
   U1525 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_21_port, B1 => 
                           n14608, B2 => REGISTERS_21_21_port, ZN => n14429);
   U1526 : AOI22_X1 port map( A1 => n14927, A2 => REGISTERS_16_21_port, B1 => 
                           n14541, B2 => REGISTERS_20_21_port, ZN => n14428);
   U1527 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_21_port, B1 => 
                           n14937, B2 => REGISTERS_24_21_port, ZN => n14427);
   U1528 : NAND4_X1 port map( A1 => n14430, A2 => n14429, A3 => n14428, A4 => 
                           n14427, ZN => n14436);
   U1529 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_21_port, B1 => 
                           n14935, B2 => REGISTERS_18_21_port, ZN => n14434);
   U1530 : AOI22_X1 port map( A1 => n14846, A2 => REGISTERS_17_21_port, B1 => 
                           n14921, B2 => REGISTERS_30_21_port, ZN => n14433);
   U1531 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_21_port, B1 => 
                           n14697, B2 => REGISTERS_19_21_port, ZN => n14432);
   U1532 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_21_port, B1 => 
                           n14678, B2 => REGISTERS_22_21_port, ZN => n14431);
   U1533 : NAND4_X1 port map( A1 => n14434, A2 => n14433, A3 => n14432, A4 => 
                           n14431, ZN => n14435);
   U1534 : NOR2_X1 port map( A1 => n14436, A2 => n14435, ZN => n14448);
   U1535 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_21_port, B1 => 
                           n14853, B2 => REGISTERS_4_21_port, ZN => n14440);
   U1536 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_21_port, B1 => 
                           n14958, B2 => REGISTERS_2_21_port, ZN => n14439);
   U1537 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_21_port, B1 => 
                           n14801, B2 => REGISTERS_3_21_port, ZN => n14438);
   U1538 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_21_port, B1 => 
                           n14876, B2 => REGISTERS_0_21_port, ZN => n14437);
   U1539 : NAND4_X1 port map( A1 => n14440, A2 => n14439, A3 => n14438, A4 => 
                           n14437, ZN => n14446);
   U1540 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_21_port, B1 => 
                           n14909, B2 => REGISTERS_9_21_port, ZN => n14444);
   U1541 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_21_port, B1 => 
                           n14904, B2 => REGISTERS_10_21_port, ZN => n14443);
   U1542 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_21_port, B1 => 
                           n14882, B2 => REGISTERS_14_21_port, ZN => n14442);
   U1543 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_11_21_port, B1 => 
                           n14665, B2 => REGISTERS_8_21_port, ZN => n14441);
   U1544 : NAND4_X1 port map( A1 => n14444, A2 => n14443, A3 => n14442, A4 => 
                           n14441, ZN => n14445);
   U1545 : AOI22_X1 port map( A1 => n14788, A2 => n14446, B1 => n14811, B2 => 
                           n14445, ZN => n14447);
   U1546 : OAI21_X1 port map( B1 => n14973, B2 => n14448, A => n14447, ZN => 
                           N438);
   U1547 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_20_port, B1 => 
                           n14697, B2 => REGISTERS_19_20_port, ZN => n14452);
   U1548 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_20_port, B1 => 
                           n14845, B2 => REGISTERS_25_20_port, ZN => n14451);
   U1549 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_20_port, B1 => 
                           n14541, B2 => REGISTERS_20_20_port, ZN => n14450);
   U1550 : AOI22_X1 port map( A1 => n14935, A2 => REGISTERS_18_20_port, B1 => 
                           n14937, B2 => REGISTERS_24_20_port, ZN => n14449);
   U1551 : NAND4_X1 port map( A1 => n14452, A2 => n14451, A3 => n14450, A4 => 
                           n14449, ZN => n14458);
   U1552 : AOI22_X1 port map( A1 => n14608, A2 => REGISTERS_21_20_port, B1 => 
                           n14702, B2 => REGISTERS_16_20_port, ZN => n14456);
   U1553 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_20_port, B1 => 
                           n14678, B2 => REGISTERS_22_20_port, ZN => n14455);
   U1554 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_20_port, B1 => 
                           n14921, B2 => REGISTERS_30_20_port, ZN => n14454);
   U1555 : AOI22_X1 port map( A1 => n14846, A2 => REGISTERS_17_20_port, B1 => 
                           n14926, B2 => REGISTERS_31_20_port, ZN => n14453);
   U1556 : NAND4_X1 port map( A1 => n14456, A2 => n14455, A3 => n14454, A4 => 
                           n14453, ZN => n14457);
   U1557 : NOR2_X1 port map( A1 => n14458, A2 => n14457, ZN => n14470);
   U1558 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_20_port, B1 => 
                           n14960, B2 => REGISTERS_6_20_port, ZN => n14462);
   U1559 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_20_port, B1 => 
                           n14910, B2 => REGISTERS_4_20_port, ZN => n14461);
   U1560 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_20_port, B1 => 
                           n14957, B2 => REGISTERS_0_20_port, ZN => n14460);
   U1561 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_20_port, B1 => 
                           n14904, B2 => REGISTERS_2_20_port, ZN => n14459);
   U1562 : NAND4_X1 port map( A1 => n14462, A2 => n14461, A3 => n14460, A4 => 
                           n14459, ZN => n14468);
   U1563 : AOI22_X1 port map( A1 => n14904, A2 => REGISTERS_10_20_port, B1 => 
                           n14876, B2 => REGISTERS_8_20_port, ZN => n14466);
   U1564 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_20_port, B1 => 
                           n14959, B2 => REGISTERS_9_20_port, ZN => n14465);
   U1565 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_20_port, B1 => 
                           n14853, B2 => REGISTERS_12_20_port, ZN => n14464);
   U1566 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_20_port, B1 => 
                           n14801, B2 => REGISTERS_11_20_port, ZN => n14463);
   U1567 : NAND4_X1 port map( A1 => n14466, A2 => n14465, A3 => n14464, A4 => 
                           n14463, ZN => n14467);
   U1568 : AOI22_X1 port map( A1 => n14788, A2 => n14468, B1 => n14968, B2 => 
                           n14467, ZN => n14469);
   U1569 : OAI21_X1 port map( B1 => n14973, B2 => n14470, A => n14469, ZN => 
                           N437);
   U1570 : AOI22_X1 port map( A1 => n14893, A2 => REGISTERS_31_19_port, B1 => 
                           n14927, B2 => REGISTERS_16_19_port, ZN => n14474);
   U1571 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_19_port, B1 => 
                           n14726, B2 => REGISTERS_30_19_port, ZN => n14473);
   U1572 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_19_port, B1 => 
                           n14935, B2 => REGISTERS_18_19_port, ZN => n14472);
   U1573 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_19_port, B1 => 
                           n14608, B2 => REGISTERS_21_19_port, ZN => n14471);
   U1574 : NAND4_X1 port map( A1 => n14474, A2 => n14473, A3 => n14472, A4 => 
                           n14471, ZN => n14480);
   U1575 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_19_port, B1 => 
                           n14937, B2 => REGISTERS_24_19_port, ZN => n14478);
   U1576 : AOI22_X1 port map( A1 => n14697, A2 => REGISTERS_19_19_port, B1 => 
                           n14933, B2 => REGISTERS_20_19_port, ZN => n14477);
   U1577 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_19_port, B1 => 
                           n14924, B2 => REGISTERS_17_19_port, ZN => n14476);
   U1578 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_19_port, B1 => 
                           n14845, B2 => REGISTERS_25_19_port, ZN => n14475);
   U1579 : NAND4_X1 port map( A1 => n14478, A2 => n14477, A3 => n14476, A4 => 
                           n14475, ZN => n14479);
   U1580 : NOR2_X1 port map( A1 => n14480, A2 => n14479, ZN => n14492);
   U1581 : CLKBUF_X1 port map( A => n14970, Z => n14813);
   U1582 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_19_port, B1 => 
                           n14911, B2 => REGISTERS_3_19_port, ZN => n14484);
   U1583 : AOI22_X1 port map( A1 => n14853, A2 => REGISTERS_4_19_port, B1 => 
                           n14909, B2 => REGISTERS_1_19_port, ZN => n14483);
   U1584 : AOI22_X1 port map( A1 => n14947, A2 => REGISTERS_2_19_port, B1 => 
                           n14665, B2 => REGISTERS_0_19_port, ZN => n14482);
   U1585 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_19_port, B1 => 
                           n14882, B2 => REGISTERS_6_19_port, ZN => n14481);
   U1586 : NAND4_X1 port map( A1 => n14484, A2 => n14483, A3 => n14482, A4 => 
                           n14481, ZN => n14490);
   U1587 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_19_port, B1 => 
                           n14960, B2 => REGISTERS_14_19_port, ZN => n14488);
   U1588 : AOI22_X1 port map( A1 => n14910, A2 => REGISTERS_12_19_port, B1 => 
                           n14957, B2 => REGISTERS_8_19_port, ZN => n14487);
   U1589 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_19_port, B1 => 
                           n14909, B2 => REGISTERS_9_19_port, ZN => n14486);
   U1590 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_19_port, B1 => 
                           n14904, B2 => REGISTERS_10_19_port, ZN => n14485);
   U1591 : NAND4_X1 port map( A1 => n14488, A2 => n14487, A3 => n14486, A4 => 
                           n14485, ZN => n14489);
   U1592 : AOI22_X1 port map( A1 => n14813, A2 => n14490, B1 => n14811, B2 => 
                           n14489, ZN => n14491);
   U1593 : OAI21_X1 port map( B1 => n14973, B2 => n14492, A => n14491, ZN => 
                           N436);
   U1594 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_18_port, B1 => 
                           n14697, B2 => REGISTERS_19_18_port, ZN => n14496);
   U1595 : AOI22_X1 port map( A1 => n14891, A2 => REGISTERS_26_18_port, B1 => 
                           n14937, B2 => REGISTERS_24_18_port, ZN => n14495);
   U1596 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_18_port, B1 => 
                           n14608, B2 => REGISTERS_21_18_port, ZN => n14494);
   U1597 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_18_port, B1 => 
                           n14924, B2 => REGISTERS_17_18_port, ZN => n14493);
   U1598 : NAND4_X1 port map( A1 => n14496, A2 => n14495, A3 => n14494, A4 => 
                           n14493, ZN => n14502);
   U1599 : AOI22_X1 port map( A1 => n14702, A2 => REGISTERS_16_18_port, B1 => 
                           n14933, B2 => REGISTERS_20_18_port, ZN => n14500);
   U1600 : AOI22_X1 port map( A1 => n14893, A2 => REGISTERS_31_18_port, B1 => 
                           n14935, B2 => REGISTERS_18_18_port, ZN => n14499);
   U1601 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_18_port, B1 => 
                           n14820, B2 => REGISTERS_27_18_port, ZN => n14498);
   U1602 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_18_port, B1 => 
                           n14726, B2 => REGISTERS_30_18_port, ZN => n14497);
   U1603 : NAND4_X1 port map( A1 => n14500, A2 => n14499, A3 => n14498, A4 => 
                           n14497, ZN => n14501);
   U1604 : NOR2_X1 port map( A1 => n14502, A2 => n14501, ZN => n14514);
   U1605 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_18_port, B1 => 
                           n14956, B2 => REGISTERS_3_18_port, ZN => n14506);
   U1606 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_18_port, B1 => 
                           n14876, B2 => REGISTERS_0_18_port, ZN => n14505);
   U1607 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_6_18_port, B1 => 
                           n14910, B2 => REGISTERS_4_18_port, ZN => n14504);
   U1608 : AOI22_X1 port map( A1 => n14959, A2 => REGISTERS_1_18_port, B1 => 
                           n14904, B2 => REGISTERS_2_18_port, ZN => n14503);
   U1609 : NAND4_X1 port map( A1 => n14506, A2 => n14505, A3 => n14504, A4 => 
                           n14503, ZN => n14512);
   U1610 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_18_port, B1 => 
                           n14665, B2 => REGISTERS_8_18_port, ZN => n14510);
   U1611 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_11_18_port, B1 => 
                           n14904, B2 => REGISTERS_10_18_port, ZN => n14509);
   U1612 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_18_port, B1 => 
                           n14961, B2 => REGISTERS_13_18_port, ZN => n14508);
   U1613 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_18_port, B1 => 
                           n14959, B2 => REGISTERS_9_18_port, ZN => n14507);
   U1614 : NAND4_X1 port map( A1 => n14510, A2 => n14509, A3 => n14508, A4 => 
                           n14507, ZN => n14511);
   U1615 : AOI22_X1 port map( A1 => n14813, A2 => n14512, B1 => n14811, B2 => 
                           n14511, ZN => n14513);
   U1616 : OAI21_X1 port map( B1 => n14973, B2 => n14514, A => n14513, ZN => 
                           N435);
   U1617 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_17_port, B1 => 
                           n14923, B2 => REGISTERS_21_17_port, ZN => n14518);
   U1618 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_17_port, B1 => 
                           n14927, B2 => REGISTERS_16_17_port, ZN => n14517);
   U1619 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_17_port, B1 => 
                           n14697, B2 => REGISTERS_19_17_port, ZN => n14516);
   U1620 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_17_port, B1 => 
                           n14726, B2 => REGISTERS_30_17_port, ZN => n14515);
   U1621 : NAND4_X1 port map( A1 => n14518, A2 => n14517, A3 => n14516, A4 => 
                           n14515, ZN => n14524);
   U1622 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_17_port, B1 => 
                           n14845, B2 => REGISTERS_25_17_port, ZN => n14522);
   U1623 : AOI22_X1 port map( A1 => n14891, A2 => REGISTERS_26_17_port, B1 => 
                           n14937, B2 => REGISTERS_24_17_port, ZN => n14521);
   U1624 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_17_port, B1 => 
                           n14926, B2 => REGISTERS_31_17_port, ZN => n14520);
   U1625 : AOI22_X1 port map( A1 => n14935, A2 => REGISTERS_18_17_port, B1 => 
                           n14933, B2 => REGISTERS_20_17_port, ZN => n14519);
   U1626 : NAND4_X1 port map( A1 => n14522, A2 => n14521, A3 => n14520, A4 => 
                           n14519, ZN => n14523);
   U1627 : NOR2_X1 port map( A1 => n14524, A2 => n14523, ZN => n14536);
   U1628 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_17_port, B1 => 
                           n14665, B2 => REGISTERS_0_17_port, ZN => n14528);
   U1629 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_3_17_port, B1 => 
                           n14910, B2 => REGISTERS_4_17_port, ZN => n14527);
   U1630 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_17_port, B1 => 
                           n14733, B2 => REGISTERS_5_17_port, ZN => n14526);
   U1631 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_6_17_port, B1 => 
                           n14904, B2 => REGISTERS_2_17_port, ZN => n14525);
   U1632 : NAND4_X1 port map( A1 => n14528, A2 => n14527, A3 => n14526, A4 => 
                           n14525, ZN => n14534);
   U1633 : AOI22_X1 port map( A1 => n14910, A2 => REGISTERS_12_17_port, B1 => 
                           n14904, B2 => REGISTERS_10_17_port, ZN => n14532);
   U1634 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_17_port, B1 => 
                           n14960, B2 => REGISTERS_14_17_port, ZN => n14531);
   U1635 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_13_17_port, B1 => 
                           n14801, B2 => REGISTERS_11_17_port, ZN => n14530);
   U1636 : AOI22_X1 port map( A1 => n14909, A2 => REGISTERS_9_17_port, B1 => 
                           n14957, B2 => REGISTERS_8_17_port, ZN => n14529);
   U1637 : NAND4_X1 port map( A1 => n14532, A2 => n14531, A3 => n14530, A4 => 
                           n14529, ZN => n14533);
   U1638 : AOI22_X1 port map( A1 => n14813, A2 => n14534, B1 => n14811, B2 => 
                           n14533, ZN => n14535);
   U1639 : OAI21_X1 port map( B1 => n14973, B2 => n14536, A => n14535, ZN => 
                           N434);
   U1640 : AOI22_X1 port map( A1 => n14653, A2 => REGISTERS_18_16_port, B1 => 
                           n14937, B2 => REGISTERS_24_16_port, ZN => n14540);
   U1641 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_16_port, B1 => 
                           n14891, B2 => REGISTERS_26_16_port, ZN => n14539);
   U1642 : AOI22_X1 port map( A1 => n14846, A2 => REGISTERS_17_16_port, B1 => 
                           n14893, B2 => REGISTERS_31_16_port, ZN => n14538);
   U1643 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_16_port, B1 => 
                           n14845, B2 => REGISTERS_25_16_port, ZN => n14537);
   U1644 : NAND4_X1 port map( A1 => n14540, A2 => n14539, A3 => n14538, A4 => 
                           n14537, ZN => n14547);
   U1645 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_16_port, B1 => 
                           n14697, B2 => REGISTERS_19_16_port, ZN => n14545);
   U1646 : AOI22_X1 port map( A1 => n14541, A2 => REGISTERS_20_16_port, B1 => 
                           n14726, B2 => REGISTERS_30_16_port, ZN => n14544);
   U1647 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_16_port, B1 => 
                           n14923, B2 => REGISTERS_21_16_port, ZN => n14543);
   U1648 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_16_port, B1 => 
                           n14927, B2 => REGISTERS_16_16_port, ZN => n14542);
   U1649 : NAND4_X1 port map( A1 => n14545, A2 => n14544, A3 => n14543, A4 => 
                           n14542, ZN => n14546);
   U1650 : NOR2_X1 port map( A1 => n14547, A2 => n14546, ZN => n14559);
   U1651 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_16_port, B1 => 
                           n14876, B2 => REGISTERS_0_16_port, ZN => n14551);
   U1652 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_16_port, B1 => 
                           n14904, B2 => REGISTERS_2_16_port, ZN => n14550);
   U1653 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_16_port, B1 => 
                           n14882, B2 => REGISTERS_6_16_port, ZN => n14549);
   U1654 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_16_port, B1 => 
                           n14909, B2 => REGISTERS_1_16_port, ZN => n14548);
   U1655 : NAND4_X1 port map( A1 => n14551, A2 => n14550, A3 => n14549, A4 => 
                           n14548, ZN => n14557);
   U1656 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_11_16_port, B1 => 
                           n14904, B2 => REGISTERS_10_16_port, ZN => n14555);
   U1657 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_16_port, B1 => 
                           n14853, B2 => REGISTERS_12_16_port, ZN => n14554);
   U1658 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_16_port, B1 => 
                           n14959, B2 => REGISTERS_9_16_port, ZN => n14553);
   U1659 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_14_16_port, B1 => 
                           n14957, B2 => REGISTERS_8_16_port, ZN => n14552);
   U1660 : NAND4_X1 port map( A1 => n14555, A2 => n14554, A3 => n14553, A4 => 
                           n14552, ZN => n14556);
   U1661 : AOI22_X1 port map( A1 => n14813, A2 => n14557, B1 => n14811, B2 => 
                           n14556, ZN => n14558);
   U1662 : OAI21_X1 port map( B1 => n14973, B2 => n14559, A => n14558, ZN => 
                           N433);
   U1663 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_15_port, B1 => 
                           n14933, B2 => REGISTERS_20_15_port, ZN => n14563);
   U1664 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_15_port, B1 => 
                           n14923, B2 => REGISTERS_21_15_port, ZN => n14562);
   U1665 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_15_port, B1 => 
                           n14726, B2 => REGISTERS_30_15_port, ZN => n14561);
   U1666 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_15_port, B1 => 
                           n14925, B2 => REGISTERS_19_15_port, ZN => n14560);
   U1667 : NAND4_X1 port map( A1 => n14563, A2 => n14562, A3 => n14561, A4 => 
                           n14560, ZN => n14569);
   U1668 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_15_port, B1 => 
                           n14927, B2 => REGISTERS_16_15_port, ZN => n14567);
   U1669 : AOI22_X1 port map( A1 => n14891, A2 => REGISTERS_26_15_port, B1 => 
                           n14935, B2 => REGISTERS_18_15_port, ZN => n14566);
   U1670 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_15_port, B1 => 
                           n14937, B2 => REGISTERS_24_15_port, ZN => n14565);
   U1671 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_15_port, B1 => 
                           n14840, B2 => REGISTERS_28_15_port, ZN => n14564);
   U1672 : NAND4_X1 port map( A1 => n14567, A2 => n14566, A3 => n14565, A4 => 
                           n14564, ZN => n14568);
   U1673 : NOR2_X1 port map( A1 => n14569, A2 => n14568, ZN => n14581);
   U1674 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_15_port, B1 => 
                           n14665, B2 => REGISTERS_0_15_port, ZN => n14573);
   U1675 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_15_port, B1 => 
                           n14801, B2 => REGISTERS_3_15_port, ZN => n14572);
   U1676 : AOI22_X1 port map( A1 => n14909, A2 => REGISTERS_1_15_port, B1 => 
                           n14904, B2 => REGISTERS_2_15_port, ZN => n14571);
   U1677 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_15_port, B1 => 
                           n14960, B2 => REGISTERS_6_15_port, ZN => n14570);
   U1678 : NAND4_X1 port map( A1 => n14573, A2 => n14572, A3 => n14571, A4 => 
                           n14570, ZN => n14579);
   U1679 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_15_port, B1 => 
                           n14910, B2 => REGISTERS_12_15_port, ZN => n14577);
   U1680 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_15_port, B1 => 
                           n14957, B2 => REGISTERS_8_15_port, ZN => n14576);
   U1681 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_15_port, B1 => 
                           n14909, B2 => REGISTERS_9_15_port, ZN => n14575);
   U1682 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_11_15_port, B1 => 
                           n14904, B2 => REGISTERS_10_15_port, ZN => n14574);
   U1683 : NAND4_X1 port map( A1 => n14577, A2 => n14576, A3 => n14575, A4 => 
                           n14574, ZN => n14578);
   U1684 : AOI22_X1 port map( A1 => n14813, A2 => n14579, B1 => n14811, B2 => 
                           n14578, ZN => n14580);
   U1685 : OAI21_X1 port map( B1 => n14920, B2 => n14581, A => n14580, ZN => 
                           N432);
   U1686 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_14_port, B1 => 
                           n14927, B2 => REGISTERS_16_14_port, ZN => n14585);
   U1687 : AOI22_X1 port map( A1 => n14608, A2 => REGISTERS_21_14_port, B1 => 
                           n14925, B2 => REGISTERS_19_14_port, ZN => n14584);
   U1688 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_14_port, B1 => 
                           n14939, B2 => REGISTERS_29_14_port, ZN => n14583);
   U1689 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_14_port, B1 => 
                           n14924, B2 => REGISTERS_17_14_port, ZN => n14582);
   U1690 : NAND4_X1 port map( A1 => n14585, A2 => n14584, A3 => n14583, A4 => 
                           n14582, ZN => n14591);
   U1691 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_14_port, B1 => 
                           n14845, B2 => REGISTERS_25_14_port, ZN => n14589);
   U1692 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_14_port, B1 => 
                           n14726, B2 => REGISTERS_30_14_port, ZN => n14588);
   U1693 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_14_port, B1 => 
                           n14933, B2 => REGISTERS_20_14_port, ZN => n14587);
   U1694 : AOI22_X1 port map( A1 => n14653, A2 => REGISTERS_18_14_port, B1 => 
                           n14937, B2 => REGISTERS_24_14_port, ZN => n14586);
   U1695 : NAND4_X1 port map( A1 => n14589, A2 => n14588, A3 => n14587, A4 => 
                           n14586, ZN => n14590);
   U1696 : NOR2_X1 port map( A1 => n14591, A2 => n14590, ZN => n14603);
   U1697 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_14_port, B1 => 
                           n14911, B2 => REGISTERS_3_14_port, ZN => n14595);
   U1698 : AOI22_X1 port map( A1 => n14959, A2 => REGISTERS_1_14_port, B1 => 
                           n14904, B2 => REGISTERS_2_14_port, ZN => n14594);
   U1699 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_14_port, B1 => 
                           n14876, B2 => REGISTERS_0_14_port, ZN => n14593);
   U1700 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_14_port, B1 => 
                           n14853, B2 => REGISTERS_4_14_port, ZN => n14592);
   U1701 : NAND4_X1 port map( A1 => n14595, A2 => n14594, A3 => n14593, A4 => 
                           n14592, ZN => n14601);
   U1702 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_9_14_port, B1 => 
                           n14876, B2 => REGISTERS_8_14_port, ZN => n14599);
   U1703 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_14_port, B1 => 
                           n14801, B2 => REGISTERS_11_14_port, ZN => n14598);
   U1704 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_14_port, B1 => 
                           n14910, B2 => REGISTERS_12_14_port, ZN => n14597);
   U1705 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_14_port, B1 => 
                           n14947, B2 => REGISTERS_10_14_port, ZN => n14596);
   U1706 : NAND4_X1 port map( A1 => n14599, A2 => n14598, A3 => n14597, A4 => 
                           n14596, ZN => n14600);
   U1707 : AOI22_X1 port map( A1 => n14813, A2 => n14601, B1 => n14811, B2 => 
                           n14600, ZN => n14602);
   U1708 : OAI21_X1 port map( B1 => n14973, B2 => n14603, A => n14602, ZN => 
                           N431);
   U1709 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_13_port, B1 => 
                           n14891, B2 => REGISTERS_26_13_port, ZN => n14607);
   U1710 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_13_port, B1 => 
                           n14933, B2 => REGISTERS_20_13_port, ZN => n14606);
   U1711 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_13_port, B1 => 
                           n14926, B2 => REGISTERS_31_13_port, ZN => n14605);
   U1712 : AOI22_X1 port map( A1 => n14678, A2 => REGISTERS_22_13_port, B1 => 
                           n14937, B2 => REGISTERS_24_13_port, ZN => n14604);
   U1713 : NAND4_X1 port map( A1 => n14607, A2 => n14606, A3 => n14605, A4 => 
                           n14604, ZN => n14614);
   U1714 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_13_port, B1 => 
                           n14924, B2 => REGISTERS_17_13_port, ZN => n14612);
   U1715 : AOI22_X1 port map( A1 => n14608, A2 => REGISTERS_21_13_port, B1 => 
                           n14935, B2 => REGISTERS_18_13_port, ZN => n14611);
   U1716 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_13_port, B1 => 
                           n14927, B2 => REGISTERS_16_13_port, ZN => n14610);
   U1717 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_13_port, B1 => 
                           n14726, B2 => REGISTERS_30_13_port, ZN => n14609);
   U1718 : NAND4_X1 port map( A1 => n14612, A2 => n14611, A3 => n14610, A4 => 
                           n14609, ZN => n14613);
   U1719 : NOR2_X1 port map( A1 => n14614, A2 => n14613, ZN => n14626);
   U1720 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_13_port, B1 => 
                           n14947, B2 => REGISTERS_2_13_port, ZN => n14618);
   U1721 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_13_port, B1 => 
                           n14665, B2 => REGISTERS_0_13_port, ZN => n14617);
   U1722 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_6_13_port, B1 => 
                           n14853, B2 => REGISTERS_4_13_port, ZN => n14616);
   U1723 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_7_13_port, B1 => 
                           n14961, B2 => REGISTERS_5_13_port, ZN => n14615);
   U1724 : NAND4_X1 port map( A1 => n14618, A2 => n14617, A3 => n14616, A4 => 
                           n14615, ZN => n14624);
   U1725 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_13_port, B1 => 
                           n14959, B2 => REGISTERS_9_13_port, ZN => n14622);
   U1726 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_11_13_port, B1 => 
                           n14957, B2 => REGISTERS_8_13_port, ZN => n14621);
   U1727 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_13_port, B1 => 
                           n14910, B2 => REGISTERS_12_13_port, ZN => n14620);
   U1728 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_13_port, B1 => 
                           n14947, B2 => REGISTERS_10_13_port, ZN => n14619);
   U1729 : NAND4_X1 port map( A1 => n14622, A2 => n14621, A3 => n14620, A4 => 
                           n14619, ZN => n14623);
   U1730 : AOI22_X1 port map( A1 => n14813, A2 => n14624, B1 => n14811, B2 => 
                           n14623, ZN => n14625);
   U1731 : OAI21_X1 port map( B1 => n14920, B2 => n14626, A => n14625, ZN => 
                           N430);
   U1732 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_12_port, B1 => 
                           n14935, B2 => REGISTERS_18_12_port, ZN => n14630);
   U1733 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_12_port, B1 => 
                           n14893, B2 => REGISTERS_31_12_port, ZN => n14629);
   U1734 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_12_port, B1 => 
                           n14726, B2 => REGISTERS_30_12_port, ZN => n14628);
   U1735 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_12_port, B1 => 
                           n14845, B2 => REGISTERS_25_12_port, ZN => n14627);
   U1736 : NAND4_X1 port map( A1 => n14630, A2 => n14629, A3 => n14628, A4 => 
                           n14627, ZN => n14636);
   U1737 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_12_port, B1 => 
                           n14927, B2 => REGISTERS_16_12_port, ZN => n14634);
   U1738 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_12_port, B1 => 
                           n14933, B2 => REGISTERS_20_12_port, ZN => n14633);
   U1739 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_12_port, B1 => 
                           n14923, B2 => REGISTERS_21_12_port, ZN => n14632);
   U1740 : AOI22_X1 port map( A1 => n14678, A2 => REGISTERS_22_12_port, B1 => 
                           n14937, B2 => REGISTERS_24_12_port, ZN => n14631);
   U1741 : NAND4_X1 port map( A1 => n14634, A2 => n14633, A3 => n14632, A4 => 
                           n14631, ZN => n14635);
   U1742 : NOR2_X1 port map( A1 => n14636, A2 => n14635, ZN => n14648);
   U1743 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_3_12_port, B1 => 
                           n14909, B2 => REGISTERS_1_12_port, ZN => n14640);
   U1744 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_12_port, B1 => 
                           n14955, B2 => REGISTERS_4_12_port, ZN => n14639);
   U1745 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_12_port, B1 => 
                           n14947, B2 => REGISTERS_2_12_port, ZN => n14638);
   U1746 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_12_port, B1 => 
                           n14876, B2 => REGISTERS_0_12_port, ZN => n14637);
   U1747 : NAND4_X1 port map( A1 => n14640, A2 => n14639, A3 => n14638, A4 => 
                           n14637, ZN => n14646);
   U1748 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_9_12_port, B1 => 
                           n14876, B2 => REGISTERS_8_12_port, ZN => n14644);
   U1749 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_12_port, B1 => 
                           n14910, B2 => REGISTERS_12_12_port, ZN => n14643);
   U1750 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_12_port, B1 => 
                           n14947, B2 => REGISTERS_10_12_port, ZN => n14642);
   U1751 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_12_port, B1 => 
                           n14956, B2 => REGISTERS_11_12_port, ZN => n14641);
   U1752 : NAND4_X1 port map( A1 => n14644, A2 => n14643, A3 => n14642, A4 => 
                           n14641, ZN => n14645);
   U1753 : AOI22_X1 port map( A1 => n14813, A2 => n14646, B1 => n14811, B2 => 
                           n14645, ZN => n14647);
   U1754 : OAI21_X1 port map( B1 => n14973, B2 => n14648, A => n14647, ZN => 
                           N429);
   U1755 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_11_port, B1 => 
                           n14926, B2 => REGISTERS_31_11_port, ZN => n14652);
   U1756 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_11_port, B1 => 
                           n14923, B2 => REGISTERS_21_11_port, ZN => n14651);
   U1757 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_11_port, B1 => 
                           n14845, B2 => REGISTERS_25_11_port, ZN => n14650);
   U1758 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_11_port, B1 => 
                           n14933, B2 => REGISTERS_20_11_port, ZN => n14649);
   U1759 : NAND4_X1 port map( A1 => n14652, A2 => n14651, A3 => n14650, A4 => 
                           n14649, ZN => n14659);
   U1760 : AOI22_X1 port map( A1 => n14653, A2 => REGISTERS_18_11_port, B1 => 
                           n14927, B2 => REGISTERS_16_11_port, ZN => n14657);
   U1761 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_11_port, B1 => 
                           n14678, B2 => REGISTERS_22_11_port, ZN => n14656);
   U1762 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_11_port, B1 => 
                           n14726, B2 => REGISTERS_30_11_port, ZN => n14655);
   U1763 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_11_port, B1 => 
                           n14937, B2 => REGISTERS_24_11_port, ZN => n14654);
   U1764 : NAND4_X1 port map( A1 => n14657, A2 => n14656, A3 => n14655, A4 => 
                           n14654, ZN => n14658);
   U1765 : NOR2_X1 port map( A1 => n14659, A2 => n14658, ZN => n14673);
   U1766 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_11_port, B1 => 
                           n14960, B2 => REGISTERS_6_11_port, ZN => n14663);
   U1767 : AOI22_X1 port map( A1 => n14947, A2 => REGISTERS_2_11_port, B1 => 
                           n14876, B2 => REGISTERS_0_11_port, ZN => n14662);
   U1768 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_11_port, B1 => 
                           n14909, B2 => REGISTERS_1_11_port, ZN => n14661);
   U1769 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_11_port, B1 => 
                           n14853, B2 => REGISTERS_4_11_port, ZN => n14660);
   U1770 : NAND4_X1 port map( A1 => n14663, A2 => n14662, A3 => n14661, A4 => 
                           n14660, ZN => n14671);
   U1771 : AOI22_X1 port map( A1 => n14910, A2 => REGISTERS_12_11_port, B1 => 
                           n14947, B2 => REGISTERS_10_11_port, ZN => n14669);
   U1772 : AOI22_X1 port map( A1 => n14664, A2 => REGISTERS_15_11_port, B1 => 
                           n14801, B2 => REGISTERS_11_11_port, ZN => n14668);
   U1773 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_13_11_port, B1 => 
                           n14960, B2 => REGISTERS_14_11_port, ZN => n14667);
   U1774 : AOI22_X1 port map( A1 => n14909, A2 => REGISTERS_9_11_port, B1 => 
                           n14665, B2 => REGISTERS_8_11_port, ZN => n14666);
   U1775 : NAND4_X1 port map( A1 => n14669, A2 => n14668, A3 => n14667, A4 => 
                           n14666, ZN => n14670);
   U1776 : AOI22_X1 port map( A1 => n14813, A2 => n14671, B1 => n14811, B2 => 
                           n14670, ZN => n14672);
   U1777 : OAI21_X1 port map( B1 => n14973, B2 => n14673, A => n14672, ZN => 
                           N428);
   U1778 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_10_port, B1 => 
                           n14937, B2 => REGISTERS_24_10_port, ZN => n14677);
   U1779 : AOI22_X1 port map( A1 => n14840, A2 => REGISTERS_28_10_port, B1 => 
                           n14893, B2 => REGISTERS_31_10_port, ZN => n14676);
   U1780 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_10_port, B1 => 
                           n14923, B2 => REGISTERS_21_10_port, ZN => n14675);
   U1781 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_10_port, B1 => 
                           n14927, B2 => REGISTERS_16_10_port, ZN => n14674);
   U1782 : NAND4_X1 port map( A1 => n14677, A2 => n14676, A3 => n14675, A4 => 
                           n14674, ZN => n14684);
   U1783 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_10_port, B1 => 
                           n14678, B2 => REGISTERS_22_10_port, ZN => n14682);
   U1784 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_10_port, B1 => 
                           n14933, B2 => REGISTERS_20_10_port, ZN => n14681);
   U1785 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_10_port, B1 => 
                           n14726, B2 => REGISTERS_30_10_port, ZN => n14680);
   U1786 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_10_port, B1 => 
                           n14935, B2 => REGISTERS_18_10_port, ZN => n14679);
   U1787 : NAND4_X1 port map( A1 => n14682, A2 => n14681, A3 => n14680, A4 => 
                           n14679, ZN => n14683);
   U1788 : NOR2_X1 port map( A1 => n14684, A2 => n14683, ZN => n14696);
   U1789 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_10_port, B1 => 
                           n14957, B2 => REGISTERS_0_10_port, ZN => n14688);
   U1790 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_10_port, B1 => 
                           n14882, B2 => REGISTERS_6_10_port, ZN => n14687);
   U1791 : AOI22_X1 port map( A1 => n14801, A2 => REGISTERS_3_10_port, B1 => 
                           n14947, B2 => REGISTERS_2_10_port, ZN => n14686);
   U1792 : AOI22_X1 port map( A1 => n14853, A2 => REGISTERS_4_10_port, B1 => 
                           n14959, B2 => REGISTERS_1_10_port, ZN => n14685);
   U1793 : NAND4_X1 port map( A1 => n14688, A2 => n14687, A3 => n14686, A4 => 
                           n14685, ZN => n14694);
   U1794 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_14_10_port, B1 => 
                           n14801, B2 => REGISTERS_11_10_port, ZN => n14692);
   U1795 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_10_port, B1 => 
                           n14947, B2 => REGISTERS_10_10_port, ZN => n14691);
   U1796 : AOI22_X1 port map( A1 => n14910, A2 => REGISTERS_12_10_port, B1 => 
                           n14876, B2 => REGISTERS_8_10_port, ZN => n14690);
   U1797 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_13_10_port, B1 => 
                           n14948, B2 => REGISTERS_9_10_port, ZN => n14689);
   U1798 : NAND4_X1 port map( A1 => n14692, A2 => n14691, A3 => n14690, A4 => 
                           n14689, ZN => n14693);
   U1799 : AOI22_X1 port map( A1 => n14813, A2 => n14694, B1 => n14811, B2 => 
                           n14693, ZN => n14695);
   U1800 : OAI21_X1 port map( B1 => n14973, B2 => n14696, A => n14695, ZN => 
                           N427);
   U1801 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_9_port, B1 => 
                           n14893, B2 => REGISTERS_31_9_port, ZN => n14701);
   U1802 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_9_port, B1 => 
                           n14846, B2 => REGISTERS_17_9_port, ZN => n14700);
   U1803 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_9_port, B1 => 
                           n14820, B2 => REGISTERS_27_9_port, ZN => n14699);
   U1804 : AOI22_X1 port map( A1 => n14697, A2 => REGISTERS_19_9_port, B1 => 
                           n14726, B2 => REGISTERS_30_9_port, ZN => n14698);
   U1805 : NAND4_X1 port map( A1 => n14701, A2 => n14700, A3 => n14699, A4 => 
                           n14698, ZN => n14708);
   U1806 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_9_port, B1 => 
                           n14928, B2 => REGISTERS_25_9_port, ZN => n14706);
   U1807 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_9_port, B1 => 
                           n14923, B2 => REGISTERS_21_9_port, ZN => n14705);
   U1808 : AOI22_X1 port map( A1 => n14702, A2 => REGISTERS_16_9_port, B1 => 
                           n14937, B2 => REGISTERS_24_9_port, ZN => n14704);
   U1809 : AOI22_X1 port map( A1 => n14935, A2 => REGISTERS_18_9_port, B1 => 
                           n14933, B2 => REGISTERS_20_9_port, ZN => n14703);
   U1810 : NAND4_X1 port map( A1 => n14706, A2 => n14705, A3 => n14704, A4 => 
                           n14703, ZN => n14707);
   U1811 : NOR2_X1 port map( A1 => n14708, A2 => n14707, ZN => n14720);
   U1812 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_9_port, B1 => 
                           n14910, B2 => REGISTERS_4_9_port, ZN => n14712);
   U1813 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_3_9_port, B1 => 
                           n14957, B2 => REGISTERS_0_9_port, ZN => n14711);
   U1814 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_9_port, B1 => 
                           n14909, B2 => REGISTERS_1_9_port, ZN => n14710);
   U1815 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_9_port, B1 => 
                           n14904, B2 => REGISTERS_2_9_port, ZN => n14709);
   U1816 : NAND4_X1 port map( A1 => n14712, A2 => n14711, A3 => n14710, A4 => 
                           n14709, ZN => n14718);
   U1817 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_9_port, B1 => 
                           n14959, B2 => REGISTERS_9_9_port, ZN => n14716);
   U1818 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_9_port, B1 => 
                           n14958, B2 => REGISTERS_10_9_port, ZN => n14715);
   U1819 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_9_port, B1 => 
                           n14876, B2 => REGISTERS_8_9_port, ZN => n14714);
   U1820 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_9_port, B1 => 
                           n14955, B2 => REGISTERS_12_9_port, ZN => n14713);
   U1821 : NAND4_X1 port map( A1 => n14716, A2 => n14715, A3 => n14714, A4 => 
                           n14713, ZN => n14717);
   U1822 : AOI22_X1 port map( A1 => n14813, A2 => n14718, B1 => n14811, B2 => 
                           n14717, ZN => n14719);
   U1823 : OAI21_X1 port map( B1 => n14920, B2 => n14720, A => n14719, ZN => 
                           N426);
   U1824 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_8_port, B1 => 
                           n14925, B2 => REGISTERS_19_8_port, ZN => n14725);
   U1825 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_8_port, B1 => 
                           n14846, B2 => REGISTERS_17_8_port, ZN => n14724);
   U1826 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_8_port, B1 => 
                           n14935, B2 => REGISTERS_18_8_port, ZN => n14723);
   U1827 : AOI22_X1 port map( A1 => n14721, A2 => REGISTERS_23_8_port, B1 => 
                           n14927, B2 => REGISTERS_16_8_port, ZN => n14722);
   U1828 : NAND4_X1 port map( A1 => n14725, A2 => n14724, A3 => n14723, A4 => 
                           n14722, ZN => n14732);
   U1829 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_8_port, B1 => 
                           n14891, B2 => REGISTERS_26_8_port, ZN => n14730);
   U1830 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_8_port, B1 => 
                           n14923, B2 => REGISTERS_21_8_port, ZN => n14729);
   U1831 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_8_port, B1 => 
                           n14937, B2 => REGISTERS_24_8_port, ZN => n14728);
   U1832 : AOI22_X1 port map( A1 => n14933, A2 => REGISTERS_20_8_port, B1 => 
                           n14726, B2 => REGISTERS_30_8_port, ZN => n14727);
   U1833 : NAND4_X1 port map( A1 => n14730, A2 => n14729, A3 => n14728, A4 => 
                           n14727, ZN => n14731);
   U1834 : NOR2_X1 port map( A1 => n14732, A2 => n14731, ZN => n14745);
   U1835 : AOI22_X1 port map( A1 => n14733, A2 => REGISTERS_5_8_port, B1 => 
                           n14882, B2 => REGISTERS_6_8_port, ZN => n14737);
   U1836 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_8_port, B1 => 
                           n14947, B2 => REGISTERS_2_8_port, ZN => n14736);
   U1837 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_8_port, B1 => 
                           n14956, B2 => REGISTERS_3_8_port, ZN => n14735);
   U1838 : AOI22_X1 port map( A1 => n14910, A2 => REGISTERS_4_8_port, B1 => 
                           n14957, B2 => REGISTERS_0_8_port, ZN => n14734);
   U1839 : NAND4_X1 port map( A1 => n14737, A2 => n14736, A3 => n14735, A4 => 
                           n14734, ZN => n14743);
   U1840 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_15_8_port, B1 => 
                           n14961, B2 => REGISTERS_13_8_port, ZN => n14741);
   U1841 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_9_8_port, B1 => 
                           n14947, B2 => REGISTERS_10_8_port, ZN => n14740);
   U1842 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_14_8_port, B1 => 
                           n14853, B2 => REGISTERS_12_8_port, ZN => n14739);
   U1843 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_8_port, B1 => 
                           n14876, B2 => REGISTERS_8_8_port, ZN => n14738);
   U1844 : NAND4_X1 port map( A1 => n14741, A2 => n14740, A3 => n14739, A4 => 
                           n14738, ZN => n14742);
   U1845 : AOI22_X1 port map( A1 => n14813, A2 => n14743, B1 => n14811, B2 => 
                           n14742, ZN => n14744);
   U1846 : OAI21_X1 port map( B1 => n14973, B2 => n14745, A => n14744, ZN => 
                           N425);
   U1847 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_7_port, B1 => 
                           n14846, B2 => REGISTERS_17_7_port, ZN => n14749);
   U1848 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_7_port, B1 => 
                           n14937, B2 => REGISTERS_24_7_port, ZN => n14748);
   U1849 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_7_port, B1 => 
                           n14935, B2 => REGISTERS_18_7_port, ZN => n14747);
   U1850 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_7_port, B1 => 
                           n14820, B2 => REGISTERS_27_7_port, ZN => n14746);
   U1851 : NAND4_X1 port map( A1 => n14749, A2 => n14748, A3 => n14747, A4 => 
                           n14746, ZN => n14755);
   U1852 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_7_port, B1 => 
                           n14925, B2 => REGISTERS_19_7_port, ZN => n14753);
   U1853 : AOI22_X1 port map( A1 => n14927, A2 => REGISTERS_16_7_port, B1 => 
                           n14921, B2 => REGISTERS_30_7_port, ZN => n14752);
   U1854 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_7_port, B1 => 
                           n14928, B2 => REGISTERS_25_7_port, ZN => n14751);
   U1855 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_7_port, B1 => 
                           n14933, B2 => REGISTERS_20_7_port, ZN => n14750);
   U1856 : NAND4_X1 port map( A1 => n14753, A2 => n14752, A3 => n14751, A4 => 
                           n14750, ZN => n14754);
   U1857 : NOR2_X1 port map( A1 => n14755, A2 => n14754, ZN => n14767);
   U1858 : AOI22_X1 port map( A1 => n14910, A2 => REGISTERS_4_7_port, B1 => 
                           n14958, B2 => REGISTERS_2_7_port, ZN => n14759);
   U1859 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_7_port, B1 => 
                           n14876, B2 => REGISTERS_0_7_port, ZN => n14758);
   U1860 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_7_port, B1 => 
                           n14948, B2 => REGISTERS_1_7_port, ZN => n14757);
   U1861 : AOI22_X1 port map( A1 => n14961, A2 => REGISTERS_5_7_port, B1 => 
                           n14956, B2 => REGISTERS_3_7_port, ZN => n14756);
   U1862 : NAND4_X1 port map( A1 => n14759, A2 => n14758, A3 => n14757, A4 => 
                           n14756, ZN => n14765);
   U1863 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_7_port, B1 => 
                           n14957, B2 => REGISTERS_8_7_port, ZN => n14763);
   U1864 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_7_port, B1 => 
                           n14947, B2 => REGISTERS_10_7_port, ZN => n14762);
   U1865 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_7_port, B1 => 
                           n14882, B2 => REGISTERS_14_7_port, ZN => n14761);
   U1866 : AOI22_X1 port map( A1 => n14853, A2 => REGISTERS_12_7_port, B1 => 
                           n14909, B2 => REGISTERS_9_7_port, ZN => n14760);
   U1867 : NAND4_X1 port map( A1 => n14763, A2 => n14762, A3 => n14761, A4 => 
                           n14760, ZN => n14764);
   U1868 : AOI22_X1 port map( A1 => n14813, A2 => n14765, B1 => n14811, B2 => 
                           n14764, ZN => n14766);
   U1869 : OAI21_X1 port map( B1 => n14920, B2 => n14767, A => n14766, ZN => 
                           N424);
   U1870 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_6_port, B1 => 
                           n14935, B2 => REGISTERS_18_6_port, ZN => n14771);
   U1871 : AOI22_X1 port map( A1 => n14839, A2 => REGISTERS_24_6_port, B1 => 
                           n14933, B2 => REGISTERS_20_6_port, ZN => n14770);
   U1872 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_6_port, B1 => 
                           n14846, B2 => REGISTERS_17_6_port, ZN => n14769);
   U1873 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_6_port, B1 => 
                           n14927, B2 => REGISTERS_16_6_port, ZN => n14768);
   U1874 : NAND4_X1 port map( A1 => n14771, A2 => n14770, A3 => n14769, A4 => 
                           n14768, ZN => n14777);
   U1875 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_6_port, B1 => 
                           n14921, B2 => REGISTERS_30_6_port, ZN => n14775);
   U1876 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_6_port, B1 => 
                           n14925, B2 => REGISTERS_19_6_port, ZN => n14774);
   U1877 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_6_port, B1 => 
                           n14923, B2 => REGISTERS_21_6_port, ZN => n14773);
   U1878 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_6_port, B1 => 
                           n14893, B2 => REGISTERS_31_6_port, ZN => n14772);
   U1879 : NAND4_X1 port map( A1 => n14775, A2 => n14774, A3 => n14773, A4 => 
                           n14772, ZN => n14776);
   U1880 : NOR2_X1 port map( A1 => n14777, A2 => n14776, ZN => n14790);
   U1881 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_6_port, B1 => 
                           n14876, B2 => REGISTERS_0_6_port, ZN => n14781);
   U1882 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_6_port, B1 => 
                           n14853, B2 => REGISTERS_4_6_port, ZN => n14780);
   U1883 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_6_6_port, B1 => 
                           n14909, B2 => REGISTERS_1_6_port, ZN => n14779);
   U1884 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_6_port, B1 => 
                           n14947, B2 => REGISTERS_2_6_port, ZN => n14778);
   U1885 : NAND4_X1 port map( A1 => n14781, A2 => n14780, A3 => n14779, A4 => 
                           n14778, ZN => n14787);
   U1886 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_14_6_port, B1 => 
                           n14957, B2 => REGISTERS_8_6_port, ZN => n14785);
   U1887 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_6_port, B1 => 
                           n14948, B2 => REGISTERS_9_6_port, ZN => n14784);
   U1888 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_6_port, B1 => 
                           n14956, B2 => REGISTERS_11_6_port, ZN => n14783);
   U1889 : AOI22_X1 port map( A1 => n14853, A2 => REGISTERS_12_6_port, B1 => 
                           n14904, B2 => REGISTERS_10_6_port, ZN => n14782);
   U1890 : NAND4_X1 port map( A1 => n14785, A2 => n14784, A3 => n14783, A4 => 
                           n14782, ZN => n14786);
   U1891 : AOI22_X1 port map( A1 => n14788, A2 => n14787, B1 => n14811, B2 => 
                           n14786, ZN => n14789);
   U1892 : OAI21_X1 port map( B1 => n14973, B2 => n14790, A => n14789, ZN => 
                           N423);
   U1893 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_5_port, B1 => 
                           n14921, B2 => REGISTERS_30_5_port, ZN => n14794);
   U1894 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_5_port, B1 => 
                           n14846, B2 => REGISTERS_17_5_port, ZN => n14793);
   U1895 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_5_port, B1 => 
                           n14820, B2 => REGISTERS_27_5_port, ZN => n14792);
   U1896 : AOI22_X1 port map( A1 => n14935, A2 => REGISTERS_18_5_port, B1 => 
                           n14933, B2 => REGISTERS_20_5_port, ZN => n14791);
   U1897 : NAND4_X1 port map( A1 => n14794, A2 => n14793, A3 => n14792, A4 => 
                           n14791, ZN => n14800);
   U1898 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_5_port, B1 => 
                           n14937, B2 => REGISTERS_24_5_port, ZN => n14798);
   U1899 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_5_port, B1 => 
                           n14928, B2 => REGISTERS_25_5_port, ZN => n14797);
   U1900 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_5_port, B1 => 
                           n14925, B2 => REGISTERS_19_5_port, ZN => n14796);
   U1901 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_5_port, B1 => 
                           n14927, B2 => REGISTERS_16_5_port, ZN => n14795);
   U1902 : NAND4_X1 port map( A1 => n14798, A2 => n14797, A3 => n14796, A4 => 
                           n14795, ZN => n14799);
   U1903 : NOR2_X1 port map( A1 => n14800, A2 => n14799, ZN => n14815);
   U1904 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_5_port, B1 => 
                           n14909, B2 => REGISTERS_1_5_port, ZN => n14805);
   U1905 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_5_port, B1 => 
                           n14876, B2 => REGISTERS_0_5_port, ZN => n14804);
   U1906 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_5_port, B1 => 
                           n14958, B2 => REGISTERS_2_5_port, ZN => n14803);
   U1907 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_5_port, B1 => 
                           n14801, B2 => REGISTERS_3_5_port, ZN => n14802);
   U1908 : NAND4_X1 port map( A1 => n14805, A2 => n14804, A3 => n14803, A4 => 
                           n14802, ZN => n14812);
   U1909 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_5_port, B1 => 
                           n14904, B2 => REGISTERS_10_5_port, ZN => n14809);
   U1910 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_5_port, B1 => 
                           n14909, B2 => REGISTERS_9_5_port, ZN => n14808);
   U1911 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_5_port, B1 => 
                           n14957, B2 => REGISTERS_8_5_port, ZN => n14807);
   U1912 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_5_port, B1 => 
                           n14955, B2 => REGISTERS_12_5_port, ZN => n14806);
   U1913 : NAND4_X1 port map( A1 => n14809, A2 => n14808, A3 => n14807, A4 => 
                           n14806, ZN => n14810);
   U1914 : AOI22_X1 port map( A1 => n14813, A2 => n14812, B1 => n14811, B2 => 
                           n14810, ZN => n14814);
   U1915 : OAI21_X1 port map( B1 => n14920, B2 => n14815, A => n14814, ZN => 
                           N422);
   U1916 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_4_port, B1 => 
                           n14921, B2 => REGISTERS_30_4_port, ZN => n14819);
   U1917 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_4_port, B1 => 
                           n14933, B2 => REGISTERS_20_4_port, ZN => n14818);
   U1918 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_4_port, B1 => 
                           n14927, B2 => REGISTERS_16_4_port, ZN => n14817);
   U1919 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_4_port, B1 => 
                           n14935, B2 => REGISTERS_18_4_port, ZN => n14816);
   U1920 : NAND4_X1 port map( A1 => n14819, A2 => n14818, A3 => n14817, A4 => 
                           n14816, ZN => n14826);
   U1921 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_4_port, B1 => 
                           n14937, B2 => REGISTERS_24_4_port, ZN => n14824);
   U1922 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_4_port, B1 => 
                           n14820, B2 => REGISTERS_27_4_port, ZN => n14823);
   U1923 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_4_port, B1 => 
                           n14891, B2 => REGISTERS_26_4_port, ZN => n14822);
   U1924 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_4_port, B1 => 
                           n14928, B2 => REGISTERS_25_4_port, ZN => n14821);
   U1925 : NAND4_X1 port map( A1 => n14824, A2 => n14823, A3 => n14822, A4 => 
                           n14821, ZN => n14825);
   U1926 : NOR2_X1 port map( A1 => n14826, A2 => n14825, ZN => n14838);
   U1927 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_4_port, B1 => 
                           n14853, B2 => REGISTERS_4_4_port, ZN => n14830);
   U1928 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_4_port, B1 => 
                           n14876, B2 => REGISTERS_0_4_port, ZN => n14829);
   U1929 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_4_port, B1 => 
                           n14948, B2 => REGISTERS_1_4_port, ZN => n14828);
   U1930 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_6_4_port, B1 => 
                           n14947, B2 => REGISTERS_2_4_port, ZN => n14827);
   U1931 : NAND4_X1 port map( A1 => n14830, A2 => n14829, A3 => n14828, A4 => 
                           n14827, ZN => n14836);
   U1932 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_4_port, B1 => 
                           n14959, B2 => REGISTERS_9_4_port, ZN => n14834);
   U1933 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_4_port, B1 => 
                           n14957, B2 => REGISTERS_8_4_port, ZN => n14833);
   U1934 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_4_port, B1 => 
                           n14958, B2 => REGISTERS_10_4_port, ZN => n14832);
   U1935 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_4_port, B1 => 
                           n14882, B2 => REGISTERS_14_4_port, ZN => n14831);
   U1936 : NAND4_X1 port map( A1 => n14834, A2 => n14833, A3 => n14832, A4 => 
                           n14831, ZN => n14835);
   U1937 : AOI22_X1 port map( A1 => n14970, A2 => n14836, B1 => n14968, B2 => 
                           n14835, ZN => n14837);
   U1938 : OAI21_X1 port map( B1 => n14973, B2 => n14838, A => n14837, ZN => 
                           N421);
   U1939 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_3_port, B1 => 
                           n14927, B2 => REGISTERS_16_3_port, ZN => n14844);
   U1940 : AOI22_X1 port map( A1 => n14839, A2 => REGISTERS_24_3_port, B1 => 
                           n14921, B2 => REGISTERS_30_3_port, ZN => n14843);
   U1941 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_3_port, B1 => 
                           n14933, B2 => REGISTERS_20_3_port, ZN => n14842);
   U1942 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_3_port, B1 => 
                           n14840, B2 => REGISTERS_28_3_port, ZN => n14841);
   U1943 : NAND4_X1 port map( A1 => n14844, A2 => n14843, A3 => n14842, A4 => 
                           n14841, ZN => n14852);
   U1944 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_3_port, B1 => 
                           n14891, B2 => REGISTERS_26_3_port, ZN => n14850);
   U1945 : AOI22_X1 port map( A1 => n14845, A2 => REGISTERS_25_3_port, B1 => 
                           n14923, B2 => REGISTERS_21_3_port, ZN => n14849);
   U1946 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_3_port, B1 => 
                           n14935, B2 => REGISTERS_18_3_port, ZN => n14848);
   U1947 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_3_port, B1 => 
                           n14846, B2 => REGISTERS_17_3_port, ZN => n14847);
   U1948 : NAND4_X1 port map( A1 => n14850, A2 => n14849, A3 => n14848, A4 => 
                           n14847, ZN => n14851);
   U1949 : NOR2_X1 port map( A1 => n14852, A2 => n14851, ZN => n14865);
   U1950 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_3_port, B1 => 
                           n14904, B2 => REGISTERS_2_3_port, ZN => n14857);
   U1951 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_3_port, B1 => 
                           n14853, B2 => REGISTERS_4_3_port, ZN => n14856);
   U1952 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_3_port, B1 => 
                           n14959, B2 => REGISTERS_1_3_port, ZN => n14855);
   U1953 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_3_port, B1 => 
                           n14876, B2 => REGISTERS_0_3_port, ZN => n14854);
   U1954 : NAND4_X1 port map( A1 => n14857, A2 => n14856, A3 => n14855, A4 => 
                           n14854, ZN => n14863);
   U1955 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_3_port, B1 => 
                           n14904, B2 => REGISTERS_10_3_port, ZN => n14861);
   U1956 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_3_port, B1 => 
                           n14959, B2 => REGISTERS_9_3_port, ZN => n14860);
   U1957 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_3_port, B1 => 
                           n14910, B2 => REGISTERS_12_3_port, ZN => n14859);
   U1958 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_3_port, B1 => 
                           n14957, B2 => REGISTERS_8_3_port, ZN => n14858);
   U1959 : NAND4_X1 port map( A1 => n14861, A2 => n14860, A3 => n14859, A4 => 
                           n14858, ZN => n14862);
   U1960 : AOI22_X1 port map( A1 => n14970, A2 => n14863, B1 => n14968, B2 => 
                           n14862, ZN => n14864);
   U1961 : OAI21_X1 port map( B1 => n14920, B2 => n14865, A => n14864, ZN => 
                           N420);
   U1962 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_2_port, B1 => 
                           n14923, B2 => REGISTERS_21_2_port, ZN => n14869);
   U1963 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_2_port, B1 => 
                           n14933, B2 => REGISTERS_20_2_port, ZN => n14868);
   U1964 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_2_port, B1 => 
                           n14928, B2 => REGISTERS_25_2_port, ZN => n14867);
   U1965 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_2_port, B1 => 
                           n14925, B2 => REGISTERS_19_2_port, ZN => n14866);
   U1966 : NAND4_X1 port map( A1 => n14869, A2 => n14868, A3 => n14867, A4 => 
                           n14866, ZN => n14875);
   U1967 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_2_port, B1 => 
                           n14935, B2 => REGISTERS_18_2_port, ZN => n14873);
   U1968 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_2_port, B1 => 
                           n14921, B2 => REGISTERS_30_2_port, ZN => n14872);
   U1969 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_2_port, B1 => 
                           n14937, B2 => REGISTERS_24_2_port, ZN => n14871);
   U1970 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_2_port, B1 => 
                           n14927, B2 => REGISTERS_16_2_port, ZN => n14870);
   U1971 : NAND4_X1 port map( A1 => n14873, A2 => n14872, A3 => n14871, A4 => 
                           n14870, ZN => n14874);
   U1972 : NOR2_X1 port map( A1 => n14875, A2 => n14874, ZN => n14890);
   U1973 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_2_port, B1 => 
                           n14876, B2 => REGISTERS_0_2_port, ZN => n14881);
   U1974 : AOI22_X1 port map( A1 => n14882, A2 => REGISTERS_6_2_port, B1 => 
                           n14956, B2 => REGISTERS_3_2_port, ZN => n14880);
   U1975 : AOI22_X1 port map( A1 => n14877, A2 => REGISTERS_7_2_port, B1 => 
                           n14948, B2 => REGISTERS_1_2_port, ZN => n14879);
   U1976 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_2_port, B1 => 
                           n14958, B2 => REGISTERS_2_2_port, ZN => n14878);
   U1977 : NAND4_X1 port map( A1 => n14881, A2 => n14880, A3 => n14879, A4 => 
                           n14878, ZN => n14888);
   U1978 : AOI22_X1 port map( A1 => n14904, A2 => REGISTERS_10_2_port, B1 => 
                           n14957, B2 => REGISTERS_8_2_port, ZN => n14886);
   U1979 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_2_port, B1 => 
                           n14956, B2 => REGISTERS_11_2_port, ZN => n14885);
   U1980 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_12_2_port, B1 => 
                           n14909, B2 => REGISTERS_9_2_port, ZN => n14884);
   U1981 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_2_port, B1 => 
                           n14882, B2 => REGISTERS_14_2_port, ZN => n14883);
   U1982 : NAND4_X1 port map( A1 => n14886, A2 => n14885, A3 => n14884, A4 => 
                           n14883, ZN => n14887);
   U1983 : AOI22_X1 port map( A1 => n14970, A2 => n14888, B1 => n14968, B2 => 
                           n14887, ZN => n14889);
   U1984 : OAI21_X1 port map( B1 => n14973, B2 => n14890, A => n14889, ZN => 
                           N419);
   U1985 : AOI22_X1 port map( A1 => n14923, A2 => REGISTERS_21_1_port, B1 => 
                           n14927, B2 => REGISTERS_16_1_port, ZN => n14897);
   U1986 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_1_port, B1 => 
                           n14891, B2 => REGISTERS_26_1_port, ZN => n14896);
   U1987 : AOI22_X1 port map( A1 => n14892, A2 => REGISTERS_29_1_port, B1 => 
                           n14928, B2 => REGISTERS_25_1_port, ZN => n14895);
   U1988 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_1_port, B1 => 
                           n14893, B2 => REGISTERS_31_1_port, ZN => n14894);
   U1989 : NAND4_X1 port map( A1 => n14897, A2 => n14896, A3 => n14895, A4 => 
                           n14894, ZN => n14903);
   U1990 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_1_port, B1 => 
                           n14921, B2 => REGISTERS_30_1_port, ZN => n14901);
   U1991 : AOI22_X1 port map( A1 => n14925, A2 => REGISTERS_19_1_port, B1 => 
                           n14935, B2 => REGISTERS_18_1_port, ZN => n14900);
   U1992 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_1_port, B1 => 
                           n14937, B2 => REGISTERS_24_1_port, ZN => n14899);
   U1993 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_1_port, B1 => 
                           n14933, B2 => REGISTERS_20_1_port, ZN => n14898);
   U1994 : NAND4_X1 port map( A1 => n14901, A2 => n14900, A3 => n14899, A4 => 
                           n14898, ZN => n14902);
   U1995 : NOR2_X1 port map( A1 => n14903, A2 => n14902, ZN => n14919);
   U1996 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_3_1_port, B1 => 
                           n14959, B2 => REGISTERS_1_1_port, ZN => n14908);
   U1997 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_1_port, B1 => 
                           n14961, B2 => REGISTERS_5_1_port, ZN => n14907);
   U1998 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_1_port, B1 => 
                           n14957, B2 => REGISTERS_0_1_port, ZN => n14906);
   U1999 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_6_1_port, B1 => 
                           n14904, B2 => REGISTERS_2_1_port, ZN => n14905);
   U2000 : NAND4_X1 port map( A1 => n14908, A2 => n14907, A3 => n14906, A4 => 
                           n14905, ZN => n14917);
   U2001 : AOI22_X1 port map( A1 => n14949, A2 => REGISTERS_14_1_port, B1 => 
                           n14909, B2 => REGISTERS_9_1_port, ZN => n14915);
   U2002 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_1_port, B1 => 
                           n14947, B2 => REGISTERS_10_1_port, ZN => n14914);
   U2003 : AOI22_X1 port map( A1 => n14911, A2 => REGISTERS_11_1_port, B1 => 
                           n14910, B2 => REGISTERS_12_1_port, ZN => n14913);
   U2004 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_13_1_port, B1 => 
                           n14957, B2 => REGISTERS_8_1_port, ZN => n14912);
   U2005 : NAND4_X1 port map( A1 => n14915, A2 => n14914, A3 => n14913, A4 => 
                           n14912, ZN => n14916);
   U2006 : AOI22_X1 port map( A1 => n14970, A2 => n14917, B1 => n14968, B2 => 
                           n14916, ZN => n14918);
   U2007 : OAI21_X1 port map( B1 => n14920, B2 => n14919, A => n14918, ZN => 
                           N418);
   U2008 : AOI22_X1 port map( A1 => n14922, A2 => REGISTERS_26_0_port, B1 => 
                           n14921, B2 => REGISTERS_30_0_port, ZN => n14932);
   U2009 : AOI22_X1 port map( A1 => n14924, A2 => REGISTERS_17_0_port, B1 => 
                           n14923, B2 => REGISTERS_21_0_port, ZN => n14931);
   U2010 : AOI22_X1 port map( A1 => n14926, A2 => REGISTERS_31_0_port, B1 => 
                           n14925, B2 => REGISTERS_19_0_port, ZN => n14930);
   U2011 : AOI22_X1 port map( A1 => n14928, A2 => REGISTERS_25_0_port, B1 => 
                           n14927, B2 => REGISTERS_16_0_port, ZN => n14929);
   U2012 : NAND4_X1 port map( A1 => n14932, A2 => n14931, A3 => n14930, A4 => 
                           n14929, ZN => n14946);
   U2013 : AOI22_X1 port map( A1 => n14934, A2 => REGISTERS_28_0_port, B1 => 
                           n14933, B2 => REGISTERS_20_0_port, ZN => n14944);
   U2014 : AOI22_X1 port map( A1 => n14936, A2 => REGISTERS_22_0_port, B1 => 
                           n14935, B2 => REGISTERS_18_0_port, ZN => n14943);
   U2015 : AOI22_X1 port map( A1 => n14938, A2 => REGISTERS_27_0_port, B1 => 
                           n14937, B2 => REGISTERS_24_0_port, ZN => n14942);
   U2016 : AOI22_X1 port map( A1 => n14940, A2 => REGISTERS_23_0_port, B1 => 
                           n14939, B2 => REGISTERS_29_0_port, ZN => n14941);
   U2017 : NAND4_X1 port map( A1 => n14944, A2 => n14943, A3 => n14942, A4 => 
                           n14941, ZN => n14945);
   U2018 : NOR2_X1 port map( A1 => n14946, A2 => n14945, ZN => n14972);
   U2019 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_7_0_port, B1 => 
                           n14956, B2 => REGISTERS_3_0_port, ZN => n14954);
   U2020 : AOI22_X1 port map( A1 => n14955, A2 => REGISTERS_4_0_port, B1 => 
                           n14957, B2 => REGISTERS_0_0_port, ZN => n14953);
   U2021 : AOI22_X1 port map( A1 => n14948, A2 => REGISTERS_1_0_port, B1 => 
                           n14947, B2 => REGISTERS_2_0_port, ZN => n14952);
   U2022 : AOI22_X1 port map( A1 => n14950, A2 => REGISTERS_5_0_port, B1 => 
                           n14949, B2 => REGISTERS_6_0_port, ZN => n14951);
   U2023 : NAND4_X1 port map( A1 => n14954, A2 => n14953, A3 => n14952, A4 => 
                           n14951, ZN => n14969);
   U2024 : AOI22_X1 port map( A1 => n14956, A2 => REGISTERS_11_0_port, B1 => 
                           n14955, B2 => REGISTERS_12_0_port, ZN => n14966);
   U2025 : AOI22_X1 port map( A1 => n14958, A2 => REGISTERS_10_0_port, B1 => 
                           n14957, B2 => REGISTERS_8_0_port, ZN => n14965);
   U2026 : AOI22_X1 port map( A1 => n14960, A2 => REGISTERS_14_0_port, B1 => 
                           n14959, B2 => REGISTERS_9_0_port, ZN => n14964);
   U2027 : AOI22_X1 port map( A1 => n14962, A2 => REGISTERS_15_0_port, B1 => 
                           n14961, B2 => REGISTERS_13_0_port, ZN => n14963);
   U2028 : NAND4_X1 port map( A1 => n14966, A2 => n14965, A3 => n14964, A4 => 
                           n14963, ZN => n14967);
   U2029 : AOI22_X1 port map( A1 => n14970, A2 => n14969, B1 => n14968, B2 => 
                           n14967, ZN => n14971);
   U2030 : OAI21_X1 port map( B1 => n14973, B2 => n14972, A => n14971, ZN => 
                           N417);
   U2031 : NAND3_X1 port map( A1 => n14005, A2 => ENABLE, A3 => RD1, ZN => 
                           n15755);
   U2032 : INV_X1 port map( A => ADD_RD1(2), ZN => n14974);
   U2033 : OR3_X1 port map( A1 => n14974, A2 => ADD_RD1(0), A3 => ADD_RD1(1), 
                           ZN => n15061);
   U2034 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n14983)
                           ;
   U2035 : NOR2_X1 port map( A1 => n15061, A2 => n14983, ZN => n15619);
   U2036 : CLKBUF_X1 port map( A => n15619, Z => n15702);
   U2037 : INV_X1 port map( A => ADD_RD1(3), ZN => n14996);
   U2038 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n14996, ZN => n14982);
   U2039 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), ZN => n14981);
   U2040 : INV_X1 port map( A => ADD_RD1(0), ZN => n14976);
   U2041 : NAND2_X1 port map( A1 => n14981, A2 => n14976, ZN => n14990);
   U2042 : NOR2_X1 port map( A1 => n14982, A2 => n14990, ZN => n15703);
   U2043 : CLKBUF_X1 port map( A => n15703, Z => n15669);
   U2044 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n15702, B1 => 
                           REGISTERS_16_31_port, B2 => n15669, ZN => n14980);
   U2045 : OR3_X1 port map( A1 => n14974, A2 => n14976, A3 => ADD_RD1(1), ZN =>
                           n15085);
   U2046 : NOR2_X1 port map( A1 => n14983, A2 => n15085, ZN => n15718);
   U2047 : CLKBUF_X1 port map( A => n15718, Z => n15596);
   U2048 : INV_X1 port map( A => ADD_RD1(1), ZN => n14975);
   U2049 : OR3_X1 port map( A1 => n14975, A2 => ADD_RD1(0), A3 => ADD_RD1(2), 
                           ZN => n15134);
   U2050 : NOR2_X1 port map( A1 => n14983, A2 => n15134, ZN => n15549);
   U2051 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n15596, B1 => 
                           REGISTERS_26_31_port, B2 => n15549, ZN => n14979);
   U2052 : OR3_X1 port map( A1 => n14976, A2 => n14974, A3 => n14975, ZN => 
                           n15019);
   U2053 : NOR2_X1 port map( A1 => n14982, A2 => n15019, ZN => n15453);
   U2054 : CLKBUF_X1 port map( A => n15453, Z => n15708);
   U2055 : NOR2_X1 port map( A1 => n14982, A2 => n15085, ZN => n15499);
   U2056 : CLKBUF_X1 port map( A => n15499, Z => n15719);
   U2057 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n15708, B1 => 
                           REGISTERS_21_31_port, B2 => n15719, ZN => n14978);
   U2058 : OR3_X1 port map( A1 => n14974, A2 => n14975, A3 => ADD_RD1(0), ZN =>
                           n15038);
   U2059 : NOR2_X1 port map( A1 => n14982, A2 => n15038, ZN => n15706);
   U2060 : CLKBUF_X1 port map( A => n15706, Z => n15676);
   U2061 : OR3_X1 port map( A1 => n14976, A2 => n14975, A3 => ADD_RD1(2), ZN =>
                           n15066);
   U2062 : NOR2_X1 port map( A1 => n14983, A2 => n15066, ZN => n15675);
   U2063 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n15676, B1 => 
                           REGISTERS_27_31_port, B2 => n15675, ZN => n14977);
   U2064 : NAND4_X1 port map( A1 => n14980, A2 => n14979, A3 => n14978, A4 => 
                           n14977, ZN => n14989);
   U2065 : NOR2_X1 port map( A1 => n14983, A2 => n15019, ZN => n15575);
   U2066 : CLKBUF_X1 port map( A => n15575, Z => n15707);
   U2067 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n14981, ZN => n14991);
   U2068 : NOR2_X1 port map( A1 => n14983, A2 => n14991, ZN => n15412);
   U2069 : CLKBUF_X1 port map( A => n15412, Z => n15701);
   U2070 : AOI22_X1 port map( A1 => REGISTERS_31_31_port, A2 => n15707, B1 => 
                           REGISTERS_25_31_port, B2 => n15701, ZN => n14987);
   U2071 : NOR2_X1 port map( A1 => n14983, A2 => n14990, ZN => n15670);
   U2072 : CLKBUF_X1 port map( A => n15670, Z => n15720);
   U2073 : NOR2_X1 port map( A1 => n14982, A2 => n15061, ZN => n15476);
   U2074 : CLKBUF_X1 port map( A => n15476, Z => n15705);
   U2075 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n15720, B1 => 
                           REGISTERS_20_31_port, B2 => n15705, ZN => n14986);
   U2076 : NOR2_X1 port map( A1 => n14982, A2 => n14991, ZN => n15407);
   U2077 : CLKBUF_X1 port map( A => n15407, Z => n15717);
   U2078 : NOR2_X1 port map( A1 => n14982, A2 => n15134, ZN => n15704);
   U2079 : CLKBUF_X1 port map( A => n15704, Z => n15677);
   U2080 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n15717, B1 => 
                           REGISTERS_18_31_port, B2 => n15677, ZN => n14985);
   U2081 : NOR2_X1 port map( A1 => n14982, A2 => n15066, ZN => n15574);
   U2082 : CLKBUF_X1 port map( A => n15574, Z => n15715);
   U2083 : NOR2_X1 port map( A1 => n14983, A2 => n15038, ZN => n15548);
   U2084 : CLKBUF_X1 port map( A => n15548, Z => n15713);
   U2085 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n15715, B1 => 
                           REGISTERS_30_31_port, B2 => n15713, ZN => n14984);
   U2086 : NAND4_X1 port map( A1 => n14987, A2 => n14986, A3 => n14985, A4 => 
                           n14984, ZN => n14988);
   U2087 : NOR2_X1 port map( A1 => n14989, A2 => n14988, ZN => n15004);
   U2088 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n15700, 
                           ZN => n15752);
   U2089 : CLKBUF_X1 port map( A => n15752, Z => n15567);
   U2090 : INV_X1 port map( A => n14990, ZN => n15637);
   U2091 : CLKBUF_X1 port map( A => n15637, Z => n15738);
   U2092 : INV_X1 port map( A => n15066, ZN => n15684);
   U2093 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n15738, B1 => 
                           REGISTERS_3_31_port, B2 => n15684, ZN => n14995);
   U2094 : INV_X1 port map( A => n15038, ZN => n15690);
   U2095 : INV_X1 port map( A => n15085, ZN => n15743);
   U2096 : AOI22_X1 port map( A1 => REGISTERS_6_31_port, A2 => n15690, B1 => 
                           REGISTERS_5_31_port, B2 => n15743, ZN => n14994);
   U2097 : INV_X1 port map( A => n15134, ZN => n15685);
   U2098 : INV_X1 port map( A => n15061, ZN => n15744);
   U2099 : AOI22_X1 port map( A1 => REGISTERS_2_31_port, A2 => n15685, B1 => 
                           REGISTERS_4_31_port, B2 => n15744, ZN => n14993);
   U2100 : INV_X1 port map( A => n15019, ZN => n15636);
   U2101 : INV_X1 port map( A => n14991, ZN => n15728);
   U2102 : CLKBUF_X1 port map( A => n15728, Z => n15660);
   U2103 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n15636, B1 => 
                           REGISTERS_1_31_port, B2 => n15660, ZN => n14992);
   U2104 : NAND4_X1 port map( A1 => n14995, A2 => n14994, A3 => n14993, A4 => 
                           n14992, ZN => n15002);
   U2105 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n14996, A3 => n15700, ZN 
                           => n15750);
   U2106 : CLKBUF_X1 port map( A => n15750, Z => n15591);
   U2107 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n15744, B1 => 
                           REGISTERS_10_31_port, B2 => n15685, ZN => n15000);
   U2108 : CLKBUF_X1 port map( A => n15637, Z => n15730);
   U2109 : INV_X1 port map( A => n15019, ZN => n15727);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n15730, B1 => 
                           REGISTERS_15_31_port, B2 => n15727, ZN => n14999);
   U2111 : INV_X1 port map( A => n15066, ZN => n15691);
   U2112 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n15691, B1 => 
                           REGISTERS_14_31_port, B2 => n15690, ZN => n14998);
   U2113 : INV_X1 port map( A => n15085, ZN => n15630);
   U2114 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n15630, B1 => 
                           REGISTERS_9_31_port, B2 => n15660, ZN => n14997);
   U2115 : NAND4_X1 port map( A1 => n15000, A2 => n14999, A3 => n14998, A4 => 
                           n14997, ZN => n15001);
   U2116 : AOI22_X1 port map( A1 => n15567, A2 => n15002, B1 => n15591, B2 => 
                           n15001, ZN => n15003);
   U2117 : OAI21_X1 port map( B1 => n15700, B2 => n15004, A => n15003, ZN => 
                           N416);
   U2118 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n15702, B1 => 
                           REGISTERS_19_30_port, B2 => n15715, ZN => n15008);
   U2119 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n15717, B1 => 
                           REGISTERS_20_30_port, B2 => n15476, ZN => n15007);
   U2120 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n15719, B1 => 
                           REGISTERS_24_30_port, B2 => n15670, ZN => n15006);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_30_30_port, A2 => n15713, B1 => 
                           REGISTERS_25_30_port, B2 => n15412, ZN => n15005);
   U2122 : NAND4_X1 port map( A1 => n15008, A2 => n15007, A3 => n15006, A4 => 
                           n15005, ZN => n15014);
   U2123 : AOI22_X1 port map( A1 => REGISTERS_31_30_port, A2 => n15707, B1 => 
                           REGISTERS_22_30_port, B2 => n15706, ZN => n15012);
   U2124 : CLKBUF_X1 port map( A => n15549, Z => n15716);
   U2125 : AOI22_X1 port map( A1 => REGISTERS_26_30_port, A2 => n15716, B1 => 
                           REGISTERS_16_30_port, B2 => n15703, ZN => n15011);
   U2126 : AOI22_X1 port map( A1 => REGISTERS_18_30_port, A2 => n15677, B1 => 
                           REGISTERS_23_30_port, B2 => n15708, ZN => n15010);
   U2127 : CLKBUF_X1 port map( A => n15675, Z => n15714);
   U2128 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n15714, B1 => 
                           REGISTERS_29_30_port, B2 => n15718, ZN => n15009);
   U2129 : NAND4_X1 port map( A1 => n15012, A2 => n15011, A3 => n15010, A4 => 
                           n15009, ZN => n15013);
   U2130 : NOR2_X1 port map( A1 => n15014, A2 => n15013, ZN => n15027);
   U2131 : AOI22_X1 port map( A1 => REGISTERS_3_30_port, A2 => n15684, B1 => 
                           REGISTERS_0_30_port, B2 => n15730, ZN => n15018);
   U2132 : INV_X1 port map( A => n15038, ZN => n15737);
   U2133 : AOI22_X1 port map( A1 => REGISTERS_6_30_port, A2 => n15737, B1 => 
                           REGISTERS_5_30_port, B2 => n15630, ZN => n15017);
   U2134 : CLKBUF_X1 port map( A => n15728, Z => n15741);
   U2135 : INV_X1 port map( A => n15061, ZN => n15732);
   U2136 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n15741, B1 => 
                           REGISTERS_4_30_port, B2 => n15732, ZN => n15016);
   U2137 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n15727, B1 => 
                           REGISTERS_2_30_port, B2 => n15685, ZN => n15015);
   U2138 : NAND4_X1 port map( A1 => n15018, A2 => n15017, A3 => n15016, A4 => 
                           n15015, ZN => n15025);
   U2139 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n15743, B1 => 
                           REGISTERS_10_30_port, B2 => n15685, ZN => n15023);
   U2140 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n15637, B1 => 
                           REGISTERS_12_30_port, B2 => n15732, ZN => n15022);
   U2141 : INV_X1 port map( A => n15019, ZN => n15739);
   U2142 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n15741, B1 => 
                           REGISTERS_15_30_port, B2 => n15739, ZN => n15021);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_14_30_port, A2 => n15690, B1 => 
                           REGISTERS_11_30_port, B2 => n15684, ZN => n15020);
   U2144 : NAND4_X1 port map( A1 => n15023, A2 => n15022, A3 => n15021, A4 => 
                           n15020, ZN => n15024);
   U2145 : AOI22_X1 port map( A1 => n15567, A2 => n15025, B1 => n15591, B2 => 
                           n15024, ZN => n15026);
   U2146 : OAI21_X1 port map( B1 => n15700, B2 => n15027, A => n15026, ZN => 
                           N415);
   U2147 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n15701, B1 => 
                           REGISTERS_18_29_port, B2 => n15704, ZN => n15031);
   U2148 : AOI22_X1 port map( A1 => REGISTERS_31_29_port, A2 => n15707, B1 => 
                           REGISTERS_24_29_port, B2 => n15670, ZN => n15030);
   U2149 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n15705, B1 => 
                           REGISTERS_17_29_port, B2 => n15717, ZN => n15029);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n15719, B1 => 
                           REGISTERS_30_29_port, B2 => n15548, ZN => n15028);
   U2151 : NAND4_X1 port map( A1 => n15031, A2 => n15030, A3 => n15029, A4 => 
                           n15028, ZN => n15037);
   U2152 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n15715, B1 => 
                           REGISTERS_16_29_port, B2 => n15703, ZN => n15035);
   U2153 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n15708, B1 => 
                           REGISTERS_26_29_port, B2 => n15716, ZN => n15034);
   U2154 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n15714, B1 => 
                           REGISTERS_22_29_port, B2 => n15706, ZN => n15033);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n15596, B1 => 
                           REGISTERS_28_29_port, B2 => n15619, ZN => n15032);
   U2156 : NAND4_X1 port map( A1 => n15035, A2 => n15034, A3 => n15033, A4 => 
                           n15032, ZN => n15036);
   U2157 : NOR2_X1 port map( A1 => n15037, A2 => n15036, ZN => n15050);
   U2158 : INV_X1 port map( A => n15038, ZN => n15631);
   U2159 : AOI22_X1 port map( A1 => REGISTERS_6_29_port, A2 => n15631, B1 => 
                           REGISTERS_1_29_port, B2 => n15660, ZN => n15042);
   U2160 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n15630, B1 => 
                           REGISTERS_3_29_port, B2 => n15691, ZN => n15041);
   U2161 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n15738, B1 => 
                           REGISTERS_4_29_port, B2 => n15732, ZN => n15040);
   U2162 : AOI22_X1 port map( A1 => REGISTERS_2_29_port, A2 => n15685, B1 => 
                           REGISTERS_7_29_port, B2 => n15739, ZN => n15039);
   U2163 : NAND4_X1 port map( A1 => n15042, A2 => n15041, A3 => n15040, A4 => 
                           n15039, ZN => n15048);
   U2164 : INV_X1 port map( A => n15134, ZN => n15742);
   U2165 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n15637, B1 => 
                           REGISTERS_10_29_port, B2 => n15742, ZN => n15046);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n15691, B1 => 
                           REGISTERS_13_29_port, B2 => n15630, ZN => n15045);
   U2167 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n15732, B1 => 
                           REGISTERS_9_29_port, B2 => n15660, ZN => n15044);
   U2168 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n15727, B1 => 
                           REGISTERS_14_29_port, B2 => n15690, ZN => n15043);
   U2169 : NAND4_X1 port map( A1 => n15046, A2 => n15045, A3 => n15044, A4 => 
                           n15043, ZN => n15047);
   U2170 : AOI22_X1 port map( A1 => n15567, A2 => n15048, B1 => n15591, B2 => 
                           n15047, ZN => n15049);
   U2171 : OAI21_X1 port map( B1 => n15700, B2 => n15050, A => n15049, ZN => 
                           N414);
   U2172 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n15717, B1 => 
                           REGISTERS_16_28_port, B2 => n15703, ZN => n15054);
   U2173 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n15701, B1 => 
                           REGISTERS_29_28_port, B2 => n15718, ZN => n15053);
   U2174 : AOI22_X1 port map( A1 => REGISTERS_22_28_port, A2 => n15676, B1 => 
                           REGISTERS_20_28_port, B2 => n15476, ZN => n15052);
   U2175 : AOI22_X1 port map( A1 => REGISTERS_30_28_port, A2 => n15713, B1 => 
                           REGISTERS_23_28_port, B2 => n15453, ZN => n15051);
   U2176 : NAND4_X1 port map( A1 => n15054, A2 => n15053, A3 => n15052, A4 => 
                           n15051, ZN => n15060);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_19_28_port, A2 => n15715, B1 => 
                           REGISTERS_21_28_port, B2 => n15499, ZN => n15058);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n15714, B1 => 
                           REGISTERS_24_28_port, B2 => n15670, ZN => n15057);
   U2179 : AOI22_X1 port map( A1 => REGISTERS_26_28_port, A2 => n15716, B1 => 
                           REGISTERS_31_28_port, B2 => n15707, ZN => n15056);
   U2180 : AOI22_X1 port map( A1 => REGISTERS_18_28_port, A2 => n15677, B1 => 
                           REGISTERS_28_28_port, B2 => n15619, ZN => n15055);
   U2181 : NAND4_X1 port map( A1 => n15058, A2 => n15057, A3 => n15056, A4 => 
                           n15055, ZN => n15059);
   U2182 : NOR2_X1 port map( A1 => n15060, A2 => n15059, ZN => n15074);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n15741, B1 => 
                           REGISTERS_6_28_port, B2 => n15690, ZN => n15065);
   U2184 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n15684, B1 => 
                           REGISTERS_0_28_port, B2 => n15637, ZN => n15064);
   U2185 : AOI22_X1 port map( A1 => REGISTERS_7_28_port, A2 => n15727, B1 => 
                           REGISTERS_2_28_port, B2 => n15742, ZN => n15063);
   U2186 : INV_X1 port map( A => n15061, ZN => n15560);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n15560, B1 => 
                           REGISTERS_5_28_port, B2 => n15630, ZN => n15062);
   U2188 : NAND4_X1 port map( A1 => n15065, A2 => n15064, A3 => n15063, A4 => 
                           n15062, ZN => n15072);
   U2189 : INV_X1 port map( A => n15066, ZN => n15740);
   U2190 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n15740, B1 => 
                           REGISTERS_8_28_port, B2 => n15730, ZN => n15070);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n15744, B1 => 
                           REGISTERS_9_28_port, B2 => n15660, ZN => n15069);
   U2192 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n15630, B1 => 
                           REGISTERS_10_28_port, B2 => n15742, ZN => n15068);
   U2193 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n15727, B1 => 
                           REGISTERS_14_28_port, B2 => n15690, ZN => n15067);
   U2194 : NAND4_X1 port map( A1 => n15070, A2 => n15069, A3 => n15068, A4 => 
                           n15067, ZN => n15071);
   U2195 : AOI22_X1 port map( A1 => n15567, A2 => n15072, B1 => n15591, B2 => 
                           n15071, ZN => n15073);
   U2196 : OAI21_X1 port map( B1 => n15700, B2 => n15074, A => n15073, ZN => 
                           N413);
   U2197 : AOI22_X1 port map( A1 => REGISTERS_22_27_port, A2 => n15676, B1 => 
                           REGISTERS_29_27_port, B2 => n15718, ZN => n15078);
   U2198 : AOI22_X1 port map( A1 => REGISTERS_30_27_port, A2 => n15713, B1 => 
                           REGISTERS_31_27_port, B2 => n15575, ZN => n15077);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n15719, B1 => 
                           REGISTERS_20_27_port, B2 => n15476, ZN => n15076);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_18_27_port, A2 => n15677, B1 => 
                           REGISTERS_27_27_port, B2 => n15675, ZN => n15075);
   U2201 : NAND4_X1 port map( A1 => n15078, A2 => n15077, A3 => n15076, A4 => 
                           n15075, ZN => n15084);
   U2202 : AOI22_X1 port map( A1 => REGISTERS_19_27_port, A2 => n15715, B1 => 
                           REGISTERS_28_27_port, B2 => n15619, ZN => n15082);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n15669, B1 => 
                           REGISTERS_25_27_port, B2 => n15412, ZN => n15081);
   U2204 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n15670, B1 => 
                           REGISTERS_17_27_port, B2 => n15407, ZN => n15080);
   U2205 : AOI22_X1 port map( A1 => REGISTERS_26_27_port, A2 => n15716, B1 => 
                           REGISTERS_23_27_port, B2 => n15453, ZN => n15079);
   U2206 : NAND4_X1 port map( A1 => n15082, A2 => n15081, A3 => n15080, A4 => 
                           n15079, ZN => n15083);
   U2207 : NOR2_X1 port map( A1 => n15084, A2 => n15083, ZN => n15097);
   U2208 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n15727, B1 => 
                           REGISTERS_4_27_port, B2 => n15732, ZN => n15089);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_2_27_port, A2 => n15685, B1 => 
                           REGISTERS_0_27_port, B2 => n15730, ZN => n15088);
   U2210 : INV_X1 port map( A => n15085, ZN => n15731);
   U2211 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n15731, B1 => 
                           REGISTERS_6_27_port, B2 => n15690, ZN => n15087);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n15741, B1 => 
                           REGISTERS_3_27_port, B2 => n15691, ZN => n15086);
   U2213 : NAND4_X1 port map( A1 => n15089, A2 => n15088, A3 => n15087, A4 => 
                           n15086, ZN => n15095);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_14_27_port, A2 => n15631, B1 => 
                           REGISTERS_13_27_port, B2 => n15630, ZN => n15093);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n15560, B1 => 
                           REGISTERS_15_27_port, B2 => n15739, ZN => n15092);
   U2216 : AOI22_X1 port map( A1 => REGISTERS_10_27_port, A2 => n15685, B1 => 
                           REGISTERS_11_27_port, B2 => n15691, ZN => n15091);
   U2217 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n15730, B1 => 
                           REGISTERS_9_27_port, B2 => n15660, ZN => n15090);
   U2218 : NAND4_X1 port map( A1 => n15093, A2 => n15092, A3 => n15091, A4 => 
                           n15090, ZN => n15094);
   U2219 : AOI22_X1 port map( A1 => n15567, A2 => n15095, B1 => n15591, B2 => 
                           n15094, ZN => n15096);
   U2220 : OAI21_X1 port map( B1 => n15700, B2 => n15097, A => n15096, ZN => 
                           N412);
   U2221 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n15669, B1 => 
                           REGISTERS_19_26_port, B2 => n15574, ZN => n15101);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n15714, B1 => 
                           REGISTERS_26_26_port, B2 => n15549, ZN => n15100);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n15701, B1 => 
                           REGISTERS_23_26_port, B2 => n15453, ZN => n15099);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_30_26_port, A2 => n15713, B1 => 
                           REGISTERS_24_26_port, B2 => n15670, ZN => n15098);
   U2225 : NAND4_X1 port map( A1 => n15101, A2 => n15100, A3 => n15099, A4 => 
                           n15098, ZN => n15107);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n15596, B1 => 
                           REGISTERS_20_26_port, B2 => n15476, ZN => n15105);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n15702, B1 => 
                           REGISTERS_22_26_port, B2 => n15706, ZN => n15104);
   U2228 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n15719, B1 => 
                           REGISTERS_31_26_port, B2 => n15575, ZN => n15103);
   U2229 : AOI22_X1 port map( A1 => REGISTERS_18_26_port, A2 => n15677, B1 => 
                           REGISTERS_17_26_port, B2 => n15407, ZN => n15102);
   U2230 : NAND4_X1 port map( A1 => n15105, A2 => n15104, A3 => n15103, A4 => 
                           n15102, ZN => n15106);
   U2231 : NOR2_X1 port map( A1 => n15107, A2 => n15106, ZN => n15119);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n15740, B1 => 
                           REGISTERS_4_26_port, B2 => n15560, ZN => n15111);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n15630, B1 => 
                           REGISTERS_1_26_port, B2 => n15728, ZN => n15110);
   U2234 : AOI22_X1 port map( A1 => REGISTERS_6_26_port, A2 => n15690, B1 => 
                           REGISTERS_2_26_port, B2 => n15742, ZN => n15109);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n15636, B1 => 
                           REGISTERS_0_26_port, B2 => n15730, ZN => n15108);
   U2236 : NAND4_X1 port map( A1 => n15111, A2 => n15110, A3 => n15109, A4 => 
                           n15108, ZN => n15117);
   U2237 : AOI22_X1 port map( A1 => REGISTERS_14_26_port, A2 => n15631, B1 => 
                           REGISTERS_9_26_port, B2 => n15660, ZN => n15115);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n15691, B1 => 
                           REGISTERS_12_26_port, B2 => n15560, ZN => n15114);
   U2239 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n15727, B1 => 
                           REGISTERS_10_26_port, B2 => n15742, ZN => n15113);
   U2240 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n15637, B1 => 
                           REGISTERS_13_26_port, B2 => n15731, ZN => n15112);
   U2241 : NAND4_X1 port map( A1 => n15115, A2 => n15114, A3 => n15113, A4 => 
                           n15112, ZN => n15116);
   U2242 : AOI22_X1 port map( A1 => n15567, A2 => n15117, B1 => n15591, B2 => 
                           n15116, ZN => n15118);
   U2243 : OAI21_X1 port map( B1 => n15700, B2 => n15119, A => n15118, ZN => 
                           N411);
   U2244 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n15714, B1 => 
                           REGISTERS_21_25_port, B2 => n15499, ZN => n15123);
   U2245 : AOI22_X1 port map( A1 => REGISTERS_23_25_port, A2 => n15708, B1 => 
                           REGISTERS_22_25_port, B2 => n15706, ZN => n15122);
   U2246 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n15715, B1 => 
                           REGISTERS_18_25_port, B2 => n15704, ZN => n15121);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_30_25_port, A2 => n15713, B1 => 
                           REGISTERS_29_25_port, B2 => n15596, ZN => n15120);
   U2248 : NAND4_X1 port map( A1 => n15123, A2 => n15122, A3 => n15121, A4 => 
                           n15120, ZN => n15129);
   U2249 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n15669, B1 => 
                           REGISTERS_20_25_port, B2 => n15476, ZN => n15127);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n15707, B1 => 
                           REGISTERS_26_25_port, B2 => n15549, ZN => n15126);
   U2251 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n15701, B1 => 
                           REGISTERS_28_25_port, B2 => n15619, ZN => n15125);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n15720, B1 => 
                           REGISTERS_17_25_port, B2 => n15407, ZN => n15124);
   U2253 : NAND4_X1 port map( A1 => n15127, A2 => n15126, A3 => n15125, A4 => 
                           n15124, ZN => n15128);
   U2254 : NOR2_X1 port map( A1 => n15129, A2 => n15128, ZN => n15142);
   U2255 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n15743, B1 => 
                           REGISTERS_0_25_port, B2 => n15730, ZN => n15133);
   U2256 : AOI22_X1 port map( A1 => REGISTERS_6_25_port, A2 => n15737, B1 => 
                           REGISTERS_2_25_port, B2 => n15742, ZN => n15132);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n15684, B1 => 
                           REGISTERS_4_25_port, B2 => n15560, ZN => n15131);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n15727, B1 => 
                           REGISTERS_1_25_port, B2 => n15728, ZN => n15130);
   U2259 : NAND4_X1 port map( A1 => n15133, A2 => n15132, A3 => n15131, A4 => 
                           n15130, ZN => n15140);
   U2260 : INV_X1 port map( A => n15134, ZN => n15729);
   U2261 : AOI22_X1 port map( A1 => REGISTERS_14_25_port, A2 => n15690, B1 => 
                           REGISTERS_10_25_port, B2 => n15729, ZN => n15138);
   U2262 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n15630, B1 => 
                           REGISTERS_12_25_port, B2 => n15560, ZN => n15137);
   U2263 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n15741, B1 => 
                           REGISTERS_15_25_port, B2 => n15636, ZN => n15136);
   U2264 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n15738, B1 => 
                           REGISTERS_11_25_port, B2 => n15691, ZN => n15135);
   U2265 : NAND4_X1 port map( A1 => n15138, A2 => n15137, A3 => n15136, A4 => 
                           n15135, ZN => n15139);
   U2266 : AOI22_X1 port map( A1 => n15567, A2 => n15140, B1 => n15591, B2 => 
                           n15139, ZN => n15141);
   U2267 : OAI21_X1 port map( B1 => n15700, B2 => n15142, A => n15141, ZN => 
                           N410);
   U2268 : AOI22_X1 port map( A1 => REGISTERS_31_24_port, A2 => n15707, B1 => 
                           REGISTERS_17_24_port, B2 => n15407, ZN => n15146);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n15701, B1 => 
                           REGISTERS_18_24_port, B2 => n15704, ZN => n15145);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n15702, B1 => 
                           REGISTERS_22_24_port, B2 => n15676, ZN => n15144);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n15705, B1 => 
                           REGISTERS_29_24_port, B2 => n15596, ZN => n15143);
   U2272 : NAND4_X1 port map( A1 => n15146, A2 => n15145, A3 => n15144, A4 => 
                           n15143, ZN => n15152);
   U2273 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n15708, B1 => 
                           REGISTERS_21_24_port, B2 => n15499, ZN => n15150);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n15669, B1 => 
                           REGISTERS_30_24_port, B2 => n15548, ZN => n15149);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_19_24_port, A2 => n15715, B1 => 
                           REGISTERS_24_24_port, B2 => n15720, ZN => n15148);
   U2276 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n15714, B1 => 
                           REGISTERS_26_24_port, B2 => n15549, ZN => n15147);
   U2277 : NAND4_X1 port map( A1 => n15150, A2 => n15149, A3 => n15148, A4 => 
                           n15147, ZN => n15151);
   U2278 : NOR2_X1 port map( A1 => n15152, A2 => n15151, ZN => n15164);
   U2279 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n15691, B1 => 
                           REGISTERS_1_24_port, B2 => n15660, ZN => n15156);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n15637, B1 => 
                           REGISTERS_7_24_port, B2 => n15739, ZN => n15155);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_6_24_port, A2 => n15631, B1 => 
                           REGISTERS_4_24_port, B2 => n15560, ZN => n15154);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_2_24_port, A2 => n15685, B1 => 
                           REGISTERS_5_24_port, B2 => n15731, ZN => n15153);
   U2283 : NAND4_X1 port map( A1 => n15156, A2 => n15155, A3 => n15154, A4 => 
                           n15153, ZN => n15162);
   U2284 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n15731, B1 => 
                           REGISTERS_12_24_port, B2 => n15560, ZN => n15160);
   U2285 : AOI22_X1 port map( A1 => REGISTERS_10_24_port, A2 => n15685, B1 => 
                           REGISTERS_9_24_port, B2 => n15728, ZN => n15159);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n15738, B1 => 
                           REGISTERS_15_24_port, B2 => n15636, ZN => n15158);
   U2287 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n15684, B1 => 
                           REGISTERS_14_24_port, B2 => n15631, ZN => n15157);
   U2288 : NAND4_X1 port map( A1 => n15160, A2 => n15159, A3 => n15158, A4 => 
                           n15157, ZN => n15161);
   U2289 : AOI22_X1 port map( A1 => n15567, A2 => n15162, B1 => n15591, B2 => 
                           n15161, ZN => n15163);
   U2290 : OAI21_X1 port map( B1 => n15700, B2 => n15164, A => n15163, ZN => 
                           N409);
   U2291 : AOI22_X1 port map( A1 => REGISTERS_27_23_port, A2 => n15675, B1 => 
                           REGISTERS_16_23_port, B2 => n15703, ZN => n15168);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n15702, B1 => 
                           REGISTERS_31_23_port, B2 => n15575, ZN => n15167);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n15705, B1 => 
                           REGISTERS_18_23_port, B2 => n15704, ZN => n15166);
   U2294 : AOI22_X1 port map( A1 => REGISTERS_22_23_port, A2 => n15676, B1 => 
                           REGISTERS_21_23_port, B2 => n15499, ZN => n15165);
   U2295 : NAND4_X1 port map( A1 => n15168, A2 => n15167, A3 => n15166, A4 => 
                           n15165, ZN => n15174);
   U2296 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n15720, B1 => 
                           REGISTERS_26_23_port, B2 => n15549, ZN => n15172);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n15717, B1 => 
                           REGISTERS_30_23_port, B2 => n15548, ZN => n15171);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n15701, B1 => 
                           REGISTERS_19_23_port, B2 => n15574, ZN => n15170);
   U2299 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n15718, B1 => 
                           REGISTERS_23_23_port, B2 => n15708, ZN => n15169);
   U2300 : NAND4_X1 port map( A1 => n15172, A2 => n15171, A3 => n15170, A4 => 
                           n15169, ZN => n15173);
   U2301 : NOR2_X1 port map( A1 => n15174, A2 => n15173, ZN => n15186);
   U2302 : AOI22_X1 port map( A1 => REGISTERS_6_23_port, A2 => n15631, B1 => 
                           REGISTERS_4_23_port, B2 => n15560, ZN => n15178);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_2_23_port, A2 => n15685, B1 => 
                           REGISTERS_1_23_port, B2 => n15660, ZN => n15177);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_3_23_port, A2 => n15740, B1 => 
                           REGISTERS_0_23_port, B2 => n15730, ZN => n15176);
   U2305 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n15743, B1 => 
                           REGISTERS_7_23_port, B2 => n15636, ZN => n15175);
   U2306 : NAND4_X1 port map( A1 => n15178, A2 => n15177, A3 => n15176, A4 => 
                           n15175, ZN => n15184);
   U2307 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n15636, B1 => 
                           REGISTERS_12_23_port, B2 => n15560, ZN => n15182);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n15731, B1 => 
                           REGISTERS_9_23_port, B2 => n15728, ZN => n15181);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n15730, B1 => 
                           REGISTERS_14_23_port, B2 => n15631, ZN => n15180);
   U2310 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n15691, B1 => 
                           REGISTERS_10_23_port, B2 => n15729, ZN => n15179);
   U2311 : NAND4_X1 port map( A1 => n15182, A2 => n15181, A3 => n15180, A4 => 
                           n15179, ZN => n15183);
   U2312 : AOI22_X1 port map( A1 => n15567, A2 => n15184, B1 => n15591, B2 => 
                           n15183, ZN => n15185);
   U2313 : OAI21_X1 port map( B1 => n15755, B2 => n15186, A => n15185, ZN => 
                           N408);
   U2314 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n15670, B1 => 
                           REGISTERS_18_22_port, B2 => n15704, ZN => n15190);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n15715, B1 => 
                           REGISTERS_22_22_port, B2 => n15676, ZN => n15189);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n15717, B1 => 
                           REGISTERS_21_22_port, B2 => n15499, ZN => n15188);
   U2317 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n15718, B1 => 
                           REGISTERS_16_22_port, B2 => n15703, ZN => n15187);
   U2318 : NAND4_X1 port map( A1 => n15190, A2 => n15189, A3 => n15188, A4 => 
                           n15187, ZN => n15196);
   U2319 : AOI22_X1 port map( A1 => REGISTERS_27_22_port, A2 => n15675, B1 => 
                           REGISTERS_20_22_port, B2 => n15476, ZN => n15194);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n15707, B1 => 
                           REGISTERS_30_22_port, B2 => n15548, ZN => n15193);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_26_22_port, A2 => n15716, B1 => 
                           REGISTERS_28_22_port, B2 => n15702, ZN => n15192);
   U2322 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n15453, B1 => 
                           REGISTERS_25_22_port, B2 => n15412, ZN => n15191);
   U2323 : NAND4_X1 port map( A1 => n15194, A2 => n15193, A3 => n15192, A4 => 
                           n15191, ZN => n15195);
   U2324 : NOR2_X1 port map( A1 => n15196, A2 => n15195, ZN => n15208);
   U2325 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n15738, B1 => 
                           REGISTERS_6_22_port, B2 => n15631, ZN => n15200);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n15727, B1 => 
                           REGISTERS_5_22_port, B2 => n15731, ZN => n15199);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n15741, B1 => 
                           REGISTERS_3_22_port, B2 => n15740, ZN => n15198);
   U2328 : AOI22_X1 port map( A1 => REGISTERS_2_22_port, A2 => n15685, B1 => 
                           REGISTERS_4_22_port, B2 => n15560, ZN => n15197);
   U2329 : NAND4_X1 port map( A1 => n15200, A2 => n15199, A3 => n15198, A4 => 
                           n15197, ZN => n15206);
   U2330 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n15741, B1 => 
                           REGISTERS_13_22_port, B2 => n15731, ZN => n15204);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n15684, B1 => 
                           REGISTERS_15_22_port, B2 => n15636, ZN => n15203);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_10_22_port, A2 => n15729, B1 => 
                           REGISTERS_14_22_port, B2 => n15631, ZN => n15202);
   U2333 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n15744, B1 => 
                           REGISTERS_8_22_port, B2 => n15637, ZN => n15201);
   U2334 : NAND4_X1 port map( A1 => n15204, A2 => n15203, A3 => n15202, A4 => 
                           n15201, ZN => n15205);
   U2335 : AOI22_X1 port map( A1 => n15567, A2 => n15206, B1 => n15591, B2 => 
                           n15205, ZN => n15207);
   U2336 : OAI21_X1 port map( B1 => n15755, B2 => n15208, A => n15207, ZN => 
                           N407);
   U2337 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n15701, B1 => 
                           REGISTERS_27_21_port, B2 => n15714, ZN => n15212);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n15676, B1 => 
                           REGISTERS_28_21_port, B2 => n15619, ZN => n15211);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n15717, B1 => 
                           REGISTERS_29_21_port, B2 => n15596, ZN => n15210);
   U2340 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n15669, B1 => 
                           REGISTERS_20_21_port, B2 => n15476, ZN => n15209);
   U2341 : NAND4_X1 port map( A1 => n15212, A2 => n15211, A3 => n15210, A4 => 
                           n15209, ZN => n15218);
   U2342 : AOI22_X1 port map( A1 => REGISTERS_26_21_port, A2 => n15716, B1 => 
                           REGISTERS_21_21_port, B2 => n15499, ZN => n15216);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_18_21_port, A2 => n15677, B1 => 
                           REGISTERS_24_21_port, B2 => n15720, ZN => n15215);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n15574, B1 => 
                           REGISTERS_23_21_port, B2 => n15453, ZN => n15214);
   U2345 : AOI22_X1 port map( A1 => REGISTERS_30_21_port, A2 => n15713, B1 => 
                           REGISTERS_31_21_port, B2 => n15575, ZN => n15213);
   U2346 : NAND4_X1 port map( A1 => n15216, A2 => n15215, A3 => n15214, A4 => 
                           n15213, ZN => n15217);
   U2347 : NOR2_X1 port map( A1 => n15218, A2 => n15217, ZN => n15230);
   U2348 : AOI22_X1 port map( A1 => REGISTERS_2_21_port, A2 => n15685, B1 => 
                           REGISTERS_3_21_port, B2 => n15740, ZN => n15222);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n15630, B1 => 
                           REGISTERS_0_21_port, B2 => n15730, ZN => n15221);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n15744, B1 => 
                           REGISTERS_6_21_port, B2 => n15631, ZN => n15220);
   U2351 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n15739, B1 => 
                           REGISTERS_1_21_port, B2 => n15660, ZN => n15219);
   U2352 : NAND4_X1 port map( A1 => n15222, A2 => n15221, A3 => n15220, A4 => 
                           n15219, ZN => n15228);
   U2353 : AOI22_X1 port map( A1 => REGISTERS_14_21_port, A2 => n15690, B1 => 
                           REGISTERS_8_21_port, B2 => n15738, ZN => n15226);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n15732, B1 => 
                           REGISTERS_15_21_port, B2 => n15636, ZN => n15225);
   U2355 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n15741, B1 => 
                           REGISTERS_11_21_port, B2 => n15740, ZN => n15224);
   U2356 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n15743, B1 => 
                           REGISTERS_10_21_port, B2 => n15729, ZN => n15223);
   U2357 : NAND4_X1 port map( A1 => n15226, A2 => n15225, A3 => n15224, A4 => 
                           n15223, ZN => n15227);
   U2358 : AOI22_X1 port map( A1 => n15567, A2 => n15228, B1 => n15591, B2 => 
                           n15227, ZN => n15229);
   U2359 : OAI21_X1 port map( B1 => n15755, B2 => n15230, A => n15229, ZN => 
                           N406);
   U2360 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n15499, B1 => 
                           REGISTERS_18_20_port, B2 => n15704, ZN => n15234);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n15702, B1 => 
                           REGISTERS_26_20_port, B2 => n15549, ZN => n15233);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n15596, B1 => 
                           REGISTERS_19_20_port, B2 => n15574, ZN => n15232);
   U2363 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n15412, B1 => 
                           REGISTERS_23_20_port, B2 => n15453, ZN => n15231);
   U2364 : NAND4_X1 port map( A1 => n15234, A2 => n15233, A3 => n15232, A4 => 
                           n15231, ZN => n15240);
   U2365 : AOI22_X1 port map( A1 => REGISTERS_22_20_port, A2 => n15676, B1 => 
                           REGISTERS_31_20_port, B2 => n15575, ZN => n15238);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n15669, B1 => 
                           REGISTERS_24_20_port, B2 => n15720, ZN => n15237);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n15714, B1 => 
                           REGISTERS_20_20_port, B2 => n15476, ZN => n15236);
   U2368 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n15407, B1 => 
                           REGISTERS_30_20_port, B2 => n15548, ZN => n15235);
   U2369 : NAND4_X1 port map( A1 => n15238, A2 => n15237, A3 => n15236, A4 => 
                           n15235, ZN => n15239);
   U2370 : NOR2_X1 port map( A1 => n15240, A2 => n15239, ZN => n15252);
   U2371 : AOI22_X1 port map( A1 => REGISTERS_3_20_port, A2 => n15691, B1 => 
                           REGISTERS_0_20_port, B2 => n15637, ZN => n15244);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n15744, B1 => 
                           REGISTERS_1_20_port, B2 => n15728, ZN => n15243);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_6_20_port, A2 => n15631, B1 => 
                           REGISTERS_2_20_port, B2 => n15685, ZN => n15242);
   U2374 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n15743, B1 => 
                           REGISTERS_7_20_port, B2 => n15739, ZN => n15241);
   U2375 : NAND4_X1 port map( A1 => n15244, A2 => n15243, A3 => n15242, A4 => 
                           n15241, ZN => n15250);
   U2376 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n15727, B1 => 
                           REGISTERS_13_20_port, B2 => n15731, ZN => n15248);
   U2377 : AOI22_X1 port map( A1 => REGISTERS_10_20_port, A2 => n15729, B1 => 
                           REGISTERS_9_20_port, B2 => n15660, ZN => n15247);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n15744, B1 => 
                           REGISTERS_11_20_port, B2 => n15740, ZN => n15246);
   U2379 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n15730, B1 => 
                           REGISTERS_14_20_port, B2 => n15631, ZN => n15245);
   U2380 : NAND4_X1 port map( A1 => n15248, A2 => n15247, A3 => n15246, A4 => 
                           n15245, ZN => n15249);
   U2381 : AOI22_X1 port map( A1 => n15567, A2 => n15250, B1 => n15750, B2 => 
                           n15249, ZN => n15251);
   U2382 : OAI21_X1 port map( B1 => n15755, B2 => n15252, A => n15251, ZN => 
                           N405);
   U2383 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n15412, B1 => 
                           REGISTERS_29_19_port, B2 => n15596, ZN => n15256);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n15407, B1 => 
                           REGISTERS_30_19_port, B2 => n15548, ZN => n15255);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n15705, B1 => 
                           REGISTERS_18_19_port, B2 => n15704, ZN => n15254);
   U2386 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n15720, B1 => 
                           REGISTERS_31_19_port, B2 => n15575, ZN => n15253);
   U2387 : NAND4_X1 port map( A1 => n15256, A2 => n15255, A3 => n15254, A4 => 
                           n15253, ZN => n15262);
   U2388 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n15715, B1 => 
                           REGISTERS_21_19_port, B2 => n15499, ZN => n15260);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n15703, B1 => 
                           REGISTERS_22_19_port, B2 => n15676, ZN => n15259);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_27_19_port, A2 => n15714, B1 => 
                           REGISTERS_26_19_port, B2 => n15549, ZN => n15258);
   U2391 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n15708, B1 => 
                           REGISTERS_28_19_port, B2 => n15702, ZN => n15257);
   U2392 : NAND4_X1 port map( A1 => n15260, A2 => n15259, A3 => n15258, A4 => 
                           n15257, ZN => n15261);
   U2393 : NOR2_X1 port map( A1 => n15262, A2 => n15261, ZN => n15274);
   U2394 : CLKBUF_X1 port map( A => n15752, Z => n15593);
   U2395 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n15728, B1 => 
                           REGISTERS_7_19_port, B2 => n15636, ZN => n15266);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n15731, B1 => 
                           REGISTERS_0_19_port, B2 => n15730, ZN => n15265);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_3_19_port, A2 => n15740, B1 => 
                           REGISTERS_6_19_port, B2 => n15631, ZN => n15264);
   U2398 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n15744, B1 => 
                           REGISTERS_2_19_port, B2 => n15729, ZN => n15263);
   U2399 : NAND4_X1 port map( A1 => n15266, A2 => n15265, A3 => n15264, A4 => 
                           n15263, ZN => n15272);
   U2400 : AOI22_X1 port map( A1 => REGISTERS_14_19_port, A2 => n15737, B1 => 
                           REGISTERS_10_19_port, B2 => n15742, ZN => n15270);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n15740, B1 => 
                           REGISTERS_15_19_port, B2 => n15636, ZN => n15269);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n15738, B1 => 
                           REGISTERS_9_19_port, B2 => n15728, ZN => n15268);
   U2403 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n15743, B1 => 
                           REGISTERS_12_19_port, B2 => n15560, ZN => n15267);
   U2404 : NAND4_X1 port map( A1 => n15270, A2 => n15269, A3 => n15268, A4 => 
                           n15267, ZN => n15271);
   U2405 : AOI22_X1 port map( A1 => n15593, A2 => n15272, B1 => n15591, B2 => 
                           n15271, ZN => n15273);
   U2406 : OAI21_X1 port map( B1 => n15755, B2 => n15274, A => n15273, ZN => 
                           N404);
   U2407 : AOI22_X1 port map( A1 => REGISTERS_26_18_port, A2 => n15549, B1 => 
                           REGISTERS_19_18_port, B2 => n15574, ZN => n15278);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_30_18_port, A2 => n15548, B1 => 
                           REGISTERS_25_18_port, B2 => n15412, ZN => n15277);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n15407, B1 => 
                           REGISTERS_21_18_port, B2 => n15499, ZN => n15276);
   U2410 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n15702, B1 => 
                           REGISTERS_29_18_port, B2 => n15596, ZN => n15275);
   U2411 : NAND4_X1 port map( A1 => n15278, A2 => n15277, A3 => n15276, A4 => 
                           n15275, ZN => n15284);
   U2412 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n15714, B1 => 
                           REGISTERS_24_18_port, B2 => n15720, ZN => n15282);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n15703, B1 => 
                           REGISTERS_23_18_port, B2 => n15453, ZN => n15281);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_18_18_port, A2 => n15677, B1 => 
                           REGISTERS_22_18_port, B2 => n15676, ZN => n15280);
   U2415 : AOI22_X1 port map( A1 => REGISTERS_31_18_port, A2 => n15575, B1 => 
                           REGISTERS_20_18_port, B2 => n15705, ZN => n15279);
   U2416 : NAND4_X1 port map( A1 => n15282, A2 => n15281, A3 => n15280, A4 => 
                           n15279, ZN => n15283);
   U2417 : NOR2_X1 port map( A1 => n15284, A2 => n15283, ZN => n15296);
   U2418 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n15731, B1 => 
                           REGISTERS_4_18_port, B2 => n15560, ZN => n15288);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n15739, B1 => 
                           REGISTERS_6_18_port, B2 => n15631, ZN => n15287);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n15691, B1 => 
                           REGISTERS_0_18_port, B2 => n15730, ZN => n15286);
   U2421 : AOI22_X1 port map( A1 => REGISTERS_2_18_port, A2 => n15685, B1 => 
                           REGISTERS_1_18_port, B2 => n15728, ZN => n15285);
   U2422 : NAND4_X1 port map( A1 => n15288, A2 => n15287, A3 => n15286, A4 => 
                           n15285, ZN => n15294);
   U2423 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n15744, B1 => 
                           REGISTERS_9_18_port, B2 => n15660, ZN => n15292);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n15637, B1 => 
                           REGISTERS_13_18_port, B2 => n15731, ZN => n15291);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n15727, B1 => 
                           REGISTERS_14_18_port, B2 => n15631, ZN => n15290);
   U2426 : AOI22_X1 port map( A1 => REGISTERS_10_18_port, A2 => n15742, B1 => 
                           REGISTERS_11_18_port, B2 => n15740, ZN => n15289);
   U2427 : NAND4_X1 port map( A1 => n15292, A2 => n15291, A3 => n15290, A4 => 
                           n15289, ZN => n15293);
   U2428 : AOI22_X1 port map( A1 => n15593, A2 => n15294, B1 => n15591, B2 => 
                           n15293, ZN => n15295);
   U2429 : OAI21_X1 port map( B1 => n15755, B2 => n15296, A => n15295, ZN => 
                           N403);
   U2430 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n15719, B1 => 
                           REGISTERS_30_17_port, B2 => n15548, ZN => n15300);
   U2431 : AOI22_X1 port map( A1 => REGISTERS_26_17_port, A2 => n15549, B1 => 
                           REGISTERS_25_17_port, B2 => n15412, ZN => n15299);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n15702, B1 => 
                           REGISTERS_19_17_port, B2 => n15574, ZN => n15298);
   U2433 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n15720, B1 => 
                           REGISTERS_18_17_port, B2 => n15704, ZN => n15297);
   U2434 : NAND4_X1 port map( A1 => n15300, A2 => n15299, A3 => n15298, A4 => 
                           n15297, ZN => n15306);
   U2435 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n15707, B1 => 
                           REGISTERS_27_17_port, B2 => n15714, ZN => n15304);
   U2436 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n15708, B1 => 
                           REGISTERS_20_17_port, B2 => n15705, ZN => n15303);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n15717, B1 => 
                           REGISTERS_22_17_port, B2 => n15676, ZN => n15302);
   U2438 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n15703, B1 => 
                           REGISTERS_29_17_port, B2 => n15596, ZN => n15301);
   U2439 : NAND4_X1 port map( A1 => n15304, A2 => n15303, A3 => n15302, A4 => 
                           n15301, ZN => n15305);
   U2440 : NOR2_X1 port map( A1 => n15306, A2 => n15305, ZN => n15318);
   U2441 : AOI22_X1 port map( A1 => REGISTERS_3_17_port, A2 => n15740, B1 => 
                           REGISTERS_5_17_port, B2 => n15731, ZN => n15310);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n15631, B1 => 
                           REGISTERS_2_17_port, B2 => n15742, ZN => n15309);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n15730, B1 => 
                           REGISTERS_7_17_port, B2 => n15636, ZN => n15308);
   U2444 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n15728, B1 => 
                           REGISTERS_4_17_port, B2 => n15560, ZN => n15307);
   U2445 : NAND4_X1 port map( A1 => n15310, A2 => n15309, A3 => n15308, A4 => 
                           n15307, ZN => n15316);
   U2446 : AOI22_X1 port map( A1 => REGISTERS_14_17_port, A2 => n15737, B1 => 
                           REGISTERS_13_17_port, B2 => n15731, ZN => n15314);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n15739, B1 => 
                           REGISTERS_9_17_port, B2 => n15728, ZN => n15313);
   U2448 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n15691, B1 => 
                           REGISTERS_8_17_port, B2 => n15738, ZN => n15312);
   U2449 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n15742, B1 => 
                           REGISTERS_12_17_port, B2 => n15732, ZN => n15311);
   U2450 : NAND4_X1 port map( A1 => n15314, A2 => n15313, A3 => n15312, A4 => 
                           n15311, ZN => n15315);
   U2451 : AOI22_X1 port map( A1 => n15593, A2 => n15316, B1 => n15591, B2 => 
                           n15315, ZN => n15317);
   U2452 : OAI21_X1 port map( B1 => n15755, B2 => n15318, A => n15317, ZN => 
                           N402);
   U2453 : AOI22_X1 port map( A1 => REGISTERS_30_16_port, A2 => n15713, B1 => 
                           REGISTERS_18_16_port, B2 => n15677, ZN => n15322);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n15669, B1 => 
                           REGISTERS_26_16_port, B2 => n15549, ZN => n15321);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n15705, B1 => 
                           REGISTERS_23_16_port, B2 => n15453, ZN => n15320);
   U2456 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n15706, B1 => 
                           REGISTERS_31_16_port, B2 => n15575, ZN => n15319);
   U2457 : NAND4_X1 port map( A1 => n15322, A2 => n15321, A3 => n15320, A4 => 
                           n15319, ZN => n15328);
   U2458 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n15596, B1 => 
                           REGISTERS_17_16_port, B2 => n15407, ZN => n15326);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n15675, B1 => 
                           REGISTERS_25_16_port, B2 => n15412, ZN => n15325);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n15715, B1 => 
                           REGISTERS_21_16_port, B2 => n15719, ZN => n15324);
   U2461 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n15619, B1 => 
                           REGISTERS_24_16_port, B2 => n15720, ZN => n15323);
   U2462 : NAND4_X1 port map( A1 => n15326, A2 => n15325, A3 => n15324, A4 => 
                           n15323, ZN => n15327);
   U2463 : NOR2_X1 port map( A1 => n15328, A2 => n15327, ZN => n15340);
   U2464 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n15691, B1 => 
                           REGISTERS_6_16_port, B2 => n15631, ZN => n15332);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_2_16_port, A2 => n15729, B1 => 
                           REGISTERS_5_16_port, B2 => n15731, ZN => n15331);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n15738, B1 => 
                           REGISTERS_4_16_port, B2 => n15732, ZN => n15330);
   U2467 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n15636, B1 => 
                           REGISTERS_1_16_port, B2 => n15660, ZN => n15329);
   U2468 : NAND4_X1 port map( A1 => n15332, A2 => n15331, A3 => n15330, A4 => 
                           n15329, ZN => n15338);
   U2469 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n15744, B1 => 
                           REGISTERS_13_16_port, B2 => n15731, ZN => n15336);
   U2470 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n15739, B1 => 
                           REGISTERS_8_16_port, B2 => n15637, ZN => n15335);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n15685, B1 => 
                           REGISTERS_9_16_port, B2 => n15728, ZN => n15334);
   U2472 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n15691, B1 => 
                           REGISTERS_14_16_port, B2 => n15631, ZN => n15333);
   U2473 : NAND4_X1 port map( A1 => n15336, A2 => n15335, A3 => n15334, A4 => 
                           n15333, ZN => n15337);
   U2474 : AOI22_X1 port map( A1 => n15593, A2 => n15338, B1 => n15591, B2 => 
                           n15337, ZN => n15339);
   U2475 : OAI21_X1 port map( B1 => n15755, B2 => n15340, A => n15339, ZN => 
                           N401);
   U2476 : AOI22_X1 port map( A1 => REGISTERS_26_15_port, A2 => n15716, B1 => 
                           REGISTERS_28_15_port, B2 => n15702, ZN => n15344);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n15720, B1 => 
                           REGISTERS_25_15_port, B2 => n15412, ZN => n15343);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_22_15_port, A2 => n15706, B1 => 
                           REGISTERS_17_15_port, B2 => n15407, ZN => n15342);
   U2479 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n15596, B1 => 
                           REGISTERS_20_15_port, B2 => n15705, ZN => n15341);
   U2480 : NAND4_X1 port map( A1 => n15344, A2 => n15343, A3 => n15342, A4 => 
                           n15341, ZN => n15350);
   U2481 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n15453, B1 => 
                           REGISTERS_27_15_port, B2 => n15714, ZN => n15348);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n15669, B1 => 
                           REGISTERS_21_15_port, B2 => n15719, ZN => n15347);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_18_15_port, A2 => n15677, B1 => 
                           REGISTERS_30_15_port, B2 => n15548, ZN => n15346);
   U2484 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n15707, B1 => 
                           REGISTERS_19_15_port, B2 => n15574, ZN => n15345);
   U2485 : NAND4_X1 port map( A1 => n15348, A2 => n15347, A3 => n15346, A4 => 
                           n15345, ZN => n15349);
   U2486 : NOR2_X1 port map( A1 => n15350, A2 => n15349, ZN => n15362);
   U2487 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n15637, B1 => 
                           REGISTERS_3_15_port, B2 => n15740, ZN => n15354);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n15741, B1 => 
                           REGISTERS_6_15_port, B2 => n15631, ZN => n15353);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n15560, B1 => 
                           REGISTERS_5_15_port, B2 => n15731, ZN => n15352);
   U2490 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n15727, B1 => 
                           REGISTERS_2_15_port, B2 => n15729, ZN => n15351);
   U2491 : NAND4_X1 port map( A1 => n15354, A2 => n15353, A3 => n15352, A4 => 
                           n15351, ZN => n15360);
   U2492 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n15744, B1 => 
                           REGISTERS_14_15_port, B2 => n15737, ZN => n15358);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n15630, B1 => 
                           REGISTERS_11_15_port, B2 => n15740, ZN => n15357);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n15660, B1 => 
                           REGISTERS_10_15_port, B2 => n15729, ZN => n15356);
   U2495 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n15727, B1 => 
                           REGISTERS_8_15_port, B2 => n15730, ZN => n15355);
   U2496 : NAND4_X1 port map( A1 => n15358, A2 => n15357, A3 => n15356, A4 => 
                           n15355, ZN => n15359);
   U2497 : AOI22_X1 port map( A1 => n15593, A2 => n15360, B1 => n15591, B2 => 
                           n15359, ZN => n15361);
   U2498 : OAI21_X1 port map( B1 => n15700, B2 => n15362, A => n15361, ZN => 
                           N400);
   U2499 : AOI22_X1 port map( A1 => REGISTERS_30_14_port, A2 => n15713, B1 => 
                           REGISTERS_19_14_port, B2 => n15574, ZN => n15366);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n15412, B1 => 
                           REGISTERS_21_14_port, B2 => n15719, ZN => n15365);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n15676, B1 => 
                           REGISTERS_17_14_port, B2 => n15407, ZN => n15364);
   U2502 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n15476, B1 => 
                           REGISTERS_16_14_port, B2 => n15703, ZN => n15363);
   U2503 : NAND4_X1 port map( A1 => n15366, A2 => n15365, A3 => n15364, A4 => 
                           n15363, ZN => n15372);
   U2504 : AOI22_X1 port map( A1 => REGISTERS_31_14_port, A2 => n15707, B1 => 
                           REGISTERS_23_14_port, B2 => n15453, ZN => n15370);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n15619, B1 => 
                           REGISTERS_29_14_port, B2 => n15596, ZN => n15369);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_26_14_port, A2 => n15716, B1 => 
                           REGISTERS_27_14_port, B2 => n15714, ZN => n15368);
   U2507 : AOI22_X1 port map( A1 => REGISTERS_18_14_port, A2 => n15704, B1 => 
                           REGISTERS_24_14_port, B2 => n15720, ZN => n15367);
   U2508 : NAND4_X1 port map( A1 => n15370, A2 => n15369, A3 => n15368, A4 => 
                           n15367, ZN => n15371);
   U2509 : NOR2_X1 port map( A1 => n15372, A2 => n15371, ZN => n15384);
   U2510 : AOI22_X1 port map( A1 => REGISTERS_2_14_port, A2 => n15729, B1 => 
                           REGISTERS_1_14_port, B2 => n15660, ZN => n15376);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n15636, B1 => 
                           REGISTERS_5_14_port, B2 => n15731, ZN => n15375);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_6_14_port, A2 => n15690, B1 => 
                           REGISTERS_4_14_port, B2 => n15732, ZN => n15374);
   U2513 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n15691, B1 => 
                           REGISTERS_0_14_port, B2 => n15637, ZN => n15373);
   U2514 : NAND4_X1 port map( A1 => n15376, A2 => n15375, A3 => n15374, A4 => 
                           n15373, ZN => n15382);
   U2515 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n15691, B1 => 
                           REGISTERS_15_14_port, B2 => n15636, ZN => n15380);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n15730, B1 => 
                           REGISTERS_14_14_port, B2 => n15737, ZN => n15379);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n15741, B1 => 
                           REGISTERS_12_14_port, B2 => n15732, ZN => n15378);
   U2518 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n15630, B1 => 
                           REGISTERS_10_14_port, B2 => n15729, ZN => n15377);
   U2519 : NAND4_X1 port map( A1 => n15380, A2 => n15379, A3 => n15378, A4 => 
                           n15377, ZN => n15381);
   U2520 : AOI22_X1 port map( A1 => n15593, A2 => n15382, B1 => n15591, B2 => 
                           n15381, ZN => n15383);
   U2521 : OAI21_X1 port map( B1 => n15755, B2 => n15384, A => n15383, ZN => 
                           N399);
   U2522 : AOI22_X1 port map( A1 => REGISTERS_27_13_port, A2 => n15714, B1 => 
                           REGISTERS_30_13_port, B2 => n15713, ZN => n15388);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n15499, B1 => 
                           REGISTERS_24_13_port, B2 => n15720, ZN => n15387);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n15669, B1 => 
                           REGISTERS_31_13_port, B2 => n15575, ZN => n15386);
   U2525 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n15717, B1 => 
                           REGISTERS_23_13_port, B2 => n15708, ZN => n15385);
   U2526 : NAND4_X1 port map( A1 => n15388, A2 => n15387, A3 => n15386, A4 => 
                           n15385, ZN => n15394);
   U2527 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n15715, B1 => 
                           REGISTERS_20_13_port, B2 => n15705, ZN => n15392);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n15701, B1 => 
                           REGISTERS_22_13_port, B2 => n15676, ZN => n15391);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_18_13_port, A2 => n15677, B1 => 
                           REGISTERS_28_13_port, B2 => n15702, ZN => n15390);
   U2530 : AOI22_X1 port map( A1 => REGISTERS_26_13_port, A2 => n15716, B1 => 
                           REGISTERS_29_13_port, B2 => n15596, ZN => n15389);
   U2531 : NAND4_X1 port map( A1 => n15392, A2 => n15391, A3 => n15390, A4 => 
                           n15389, ZN => n15393);
   U2532 : NOR2_X1 port map( A1 => n15394, A2 => n15393, ZN => n15406);
   U2533 : AOI22_X1 port map( A1 => REGISTERS_3_13_port, A2 => n15691, B1 => 
                           REGISTERS_6_13_port, B2 => n15737, ZN => n15398);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n15660, B1 => 
                           REGISTERS_7_13_port, B2 => n15636, ZN => n15397);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n15738, B1 => 
                           REGISTERS_5_13_port, B2 => n15743, ZN => n15396);
   U2536 : AOI22_X1 port map( A1 => REGISTERS_2_13_port, A2 => n15742, B1 => 
                           REGISTERS_4_13_port, B2 => n15732, ZN => n15395);
   U2537 : NAND4_X1 port map( A1 => n15398, A2 => n15397, A3 => n15396, A4 => 
                           n15395, ZN => n15404);
   U2538 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n15739, B1 => 
                           REGISTERS_12_13_port, B2 => n15732, ZN => n15402);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n15637, B1 => 
                           REGISTERS_11_13_port, B2 => n15740, ZN => n15401);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n15728, B1 => 
                           REGISTERS_10_13_port, B2 => n15729, ZN => n15400);
   U2541 : AOI22_X1 port map( A1 => REGISTERS_14_13_port, A2 => n15690, B1 => 
                           REGISTERS_13_13_port, B2 => n15743, ZN => n15399);
   U2542 : NAND4_X1 port map( A1 => n15402, A2 => n15401, A3 => n15400, A4 => 
                           n15399, ZN => n15403);
   U2543 : AOI22_X1 port map( A1 => n15593, A2 => n15404, B1 => n15591, B2 => 
                           n15403, ZN => n15405);
   U2544 : OAI21_X1 port map( B1 => n15700, B2 => n15406, A => n15405, ZN => 
                           N398);
   U2545 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n15705, B1 => 
                           REGISTERS_21_12_port, B2 => n15719, ZN => n15411);
   U2546 : AOI22_X1 port map( A1 => REGISTERS_26_12_port, A2 => n15716, B1 => 
                           REGISTERS_17_12_port, B2 => n15407, ZN => n15410);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n15669, B1 => 
                           REGISTERS_23_12_port, B2 => n15708, ZN => n15409);
   U2548 : AOI22_X1 port map( A1 => REGISTERS_22_12_port, A2 => n15676, B1 => 
                           REGISTERS_24_12_port, B2 => n15720, ZN => n15408);
   U2549 : NAND4_X1 port map( A1 => n15411, A2 => n15410, A3 => n15409, A4 => 
                           n15408, ZN => n15418);
   U2550 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n15714, B1 => 
                           REGISTERS_18_12_port, B2 => n15677, ZN => n15416);
   U2551 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n15619, B1 => 
                           REGISTERS_19_12_port, B2 => n15574, ZN => n15415);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_31_12_port, A2 => n15707, B1 => 
                           REGISTERS_30_12_port, B2 => n15713, ZN => n15414);
   U2553 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n15596, B1 => 
                           REGISTERS_25_12_port, B2 => n15412, ZN => n15413);
   U2554 : NAND4_X1 port map( A1 => n15416, A2 => n15415, A3 => n15414, A4 => 
                           n15413, ZN => n15417);
   U2555 : NOR2_X1 port map( A1 => n15418, A2 => n15417, ZN => n15430);
   U2556 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n15560, B1 => 
                           REGISTERS_7_12_port, B2 => n15636, ZN => n15422);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n15728, B1 => 
                           REGISTERS_2_12_port, B2 => n15729, ZN => n15421);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_6_12_port, A2 => n15737, B1 => 
                           REGISTERS_0_12_port, B2 => n15738, ZN => n15420);
   U2559 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n15691, B1 => 
                           REGISTERS_5_12_port, B2 => n15743, ZN => n15419);
   U2560 : NAND4_X1 port map( A1 => n15422, A2 => n15421, A3 => n15420, A4 => 
                           n15419, ZN => n15428);
   U2561 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n15727, B1 => 
                           REGISTERS_11_12_port, B2 => n15740, ZN => n15426);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n15744, B1 => 
                           REGISTERS_10_12_port, B2 => n15729, ZN => n15425);
   U2563 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n15728, B1 => 
                           REGISTERS_13_12_port, B2 => n15743, ZN => n15424);
   U2564 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n15637, B1 => 
                           REGISTERS_14_12_port, B2 => n15737, ZN => n15423);
   U2565 : NAND4_X1 port map( A1 => n15426, A2 => n15425, A3 => n15424, A4 => 
                           n15423, ZN => n15427);
   U2566 : AOI22_X1 port map( A1 => n15593, A2 => n15428, B1 => n15591, B2 => 
                           n15427, ZN => n15429);
   U2567 : OAI21_X1 port map( B1 => n15755, B2 => n15430, A => n15429, ZN => 
                           N397);
   U2568 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n15669, B1 => 
                           REGISTERS_23_11_port, B2 => n15708, ZN => n15434);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n15702, B1 => 
                           REGISTERS_19_11_port, B2 => n15715, ZN => n15433);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n15596, B1 => 
                           REGISTERS_21_11_port, B2 => n15719, ZN => n15432);
   U2571 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n15717, B1 => 
                           REGISTERS_25_11_port, B2 => n15701, ZN => n15431);
   U2572 : NAND4_X1 port map( A1 => n15434, A2 => n15433, A3 => n15432, A4 => 
                           n15431, ZN => n15440);
   U2573 : AOI22_X1 port map( A1 => REGISTERS_22_11_port, A2 => n15676, B1 => 
                           REGISTERS_18_11_port, B2 => n15677, ZN => n15438);
   U2574 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n15720, B1 => 
                           REGISTERS_27_11_port, B2 => n15714, ZN => n15437);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_31_11_port, A2 => n15707, B1 => 
                           REGISTERS_20_11_port, B2 => n15705, ZN => n15436);
   U2576 : AOI22_X1 port map( A1 => REGISTERS_26_11_port, A2 => n15716, B1 => 
                           REGISTERS_30_11_port, B2 => n15713, ZN => n15435);
   U2577 : NAND4_X1 port map( A1 => n15438, A2 => n15437, A3 => n15436, A4 => 
                           n15435, ZN => n15439);
   U2578 : NOR2_X1 port map( A1 => n15440, A2 => n15439, ZN => n15452);
   U2579 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n15636, B1 => 
                           REGISTERS_0_11_port, B2 => n15730, ZN => n15444);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n15684, B1 => 
                           REGISTERS_4_11_port, B2 => n15732, ZN => n15443);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_2_11_port, A2 => n15729, B1 => 
                           REGISTERS_5_11_port, B2 => n15743, ZN => n15442);
   U2582 : AOI22_X1 port map( A1 => REGISTERS_6_11_port, A2 => n15690, B1 => 
                           REGISTERS_1_11_port, B2 => n15741, ZN => n15441);
   U2583 : NAND4_X1 port map( A1 => n15444, A2 => n15443, A3 => n15442, A4 => 
                           n15441, ZN => n15450);
   U2584 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n15732, B1 => 
                           REGISTERS_14_11_port, B2 => n15737, ZN => n15448);
   U2585 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n15684, B1 => 
                           REGISTERS_8_11_port, B2 => n15637, ZN => n15447);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n15731, B1 => 
                           REGISTERS_9_11_port, B2 => n15660, ZN => n15446);
   U2587 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n15685, B1 => 
                           REGISTERS_15_11_port, B2 => n15636, ZN => n15445);
   U2588 : NAND4_X1 port map( A1 => n15448, A2 => n15447, A3 => n15446, A4 => 
                           n15445, ZN => n15449);
   U2589 : AOI22_X1 port map( A1 => n15593, A2 => n15450, B1 => n15591, B2 => 
                           n15449, ZN => n15451);
   U2590 : OAI21_X1 port map( B1 => n15755, B2 => n15452, A => n15451, ZN => 
                           N396);
   U2591 : AOI22_X1 port map( A1 => REGISTERS_18_10_port, A2 => n15677, B1 => 
                           REGISTERS_17_10_port, B2 => n15717, ZN => n15457);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n15707, B1 => 
                           REGISTERS_21_10_port, B2 => n15719, ZN => n15456);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n15476, B1 => 
                           REGISTERS_22_10_port, B2 => n15676, ZN => n15455);
   U2594 : AOI22_X1 port map( A1 => REGISTERS_23_10_port, A2 => n15453, B1 => 
                           REGISTERS_19_10_port, B2 => n15715, ZN => n15454);
   U2595 : NAND4_X1 port map( A1 => n15457, A2 => n15456, A3 => n15455, A4 => 
                           n15454, ZN => n15463);
   U2596 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n15701, B1 => 
                           REGISTERS_29_10_port, B2 => n15596, ZN => n15461);
   U2597 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n15702, B1 => 
                           REGISTERS_27_10_port, B2 => n15714, ZN => n15460);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_26_10_port, A2 => n15716, B1 => 
                           REGISTERS_24_10_port, B2 => n15720, ZN => n15459);
   U2599 : AOI22_X1 port map( A1 => REGISTERS_30_10_port, A2 => n15713, B1 => 
                           REGISTERS_16_10_port, B2 => n15703, ZN => n15458);
   U2600 : NAND4_X1 port map( A1 => n15461, A2 => n15460, A3 => n15459, A4 => 
                           n15458, ZN => n15462);
   U2601 : NOR2_X1 port map( A1 => n15463, A2 => n15462, ZN => n15475);
   U2602 : AOI22_X1 port map( A1 => REGISTERS_3_10_port, A2 => n15684, B1 => 
                           REGISTERS_4_10_port, B2 => n15560, ZN => n15467);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n15630, B1 => 
                           REGISTERS_7_10_port, B2 => n15739, ZN => n15466);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_6_10_port, A2 => n15737, B1 => 
                           REGISTERS_1_10_port, B2 => n15728, ZN => n15465);
   U2605 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n15738, B1 => 
                           REGISTERS_2_10_port, B2 => n15729, ZN => n15464);
   U2606 : NAND4_X1 port map( A1 => n15467, A2 => n15466, A3 => n15465, A4 => 
                           n15464, ZN => n15473);
   U2607 : AOI22_X1 port map( A1 => REGISTERS_10_10_port, A2 => n15685, B1 => 
                           REGISTERS_8_10_port, B2 => n15637, ZN => n15471);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n15739, B1 => 
                           REGISTERS_12_10_port, B2 => n15560, ZN => n15470);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n15630, B1 => 
                           REGISTERS_9_10_port, B2 => n15728, ZN => n15469);
   U2610 : AOI22_X1 port map( A1 => REGISTERS_14_10_port, A2 => n15690, B1 => 
                           REGISTERS_11_10_port, B2 => n15740, ZN => n15468);
   U2611 : NAND4_X1 port map( A1 => n15471, A2 => n15470, A3 => n15469, A4 => 
                           n15468, ZN => n15472);
   U2612 : AOI22_X1 port map( A1 => n15593, A2 => n15473, B1 => n15591, B2 => 
                           n15472, ZN => n15474);
   U2613 : OAI21_X1 port map( B1 => n15755, B2 => n15475, A => n15474, ZN => 
                           N395);
   U2614 : AOI22_X1 port map( A1 => REGISTERS_26_9_port, A2 => n15716, B1 => 
                           REGISTERS_17_9_port, B2 => n15717, ZN => n15480);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n15476, B1 => 
                           REGISTERS_30_9_port, B2 => n15713, ZN => n15479);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n15701, B1 => 
                           REGISTERS_24_9_port, B2 => n15720, ZN => n15478);
   U2617 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n15707, B1 => 
                           REGISTERS_23_9_port, B2 => n15708, ZN => n15477);
   U2618 : NAND4_X1 port map( A1 => n15480, A2 => n15479, A3 => n15478, A4 => 
                           n15477, ZN => n15486);
   U2619 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n15702, B1 => 
                           REGISTERS_29_9_port, B2 => n15596, ZN => n15484);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_18_9_port, A2 => n15704, B1 => 
                           REGISTERS_27_9_port, B2 => n15675, ZN => n15483);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n15669, B1 => 
                           REGISTERS_22_9_port, B2 => n15706, ZN => n15482);
   U2622 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n15719, B1 => 
                           REGISTERS_19_9_port, B2 => n15715, ZN => n15481);
   U2623 : NAND4_X1 port map( A1 => n15484, A2 => n15483, A3 => n15482, A4 => 
                           n15481, ZN => n15485);
   U2624 : NOR2_X1 port map( A1 => n15486, A2 => n15485, ZN => n15498);
   U2625 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n15684, B1 => 
                           REGISTERS_1_9_port, B2 => n15660, ZN => n15490);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n15738, B1 => 
                           REGISTERS_6_9_port, B2 => n15737, ZN => n15489);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n15727, B1 => 
                           REGISTERS_5_9_port, B2 => n15743, ZN => n15488);
   U2628 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n15744, B1 => 
                           REGISTERS_2_9_port, B2 => n15729, ZN => n15487);
   U2629 : NAND4_X1 port map( A1 => n15490, A2 => n15489, A3 => n15488, A4 => 
                           n15487, ZN => n15496);
   U2630 : AOI22_X1 port map( A1 => REGISTERS_10_9_port, A2 => n15742, B1 => 
                           REGISTERS_12_9_port, B2 => n15744, ZN => n15494);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n15636, B1 => 
                           REGISTERS_11_9_port, B2 => n15740, ZN => n15493);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_14_9_port, A2 => n15690, B1 => 
                           REGISTERS_8_9_port, B2 => n15637, ZN => n15492);
   U2633 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n15728, B1 => 
                           REGISTERS_13_9_port, B2 => n15743, ZN => n15491);
   U2634 : NAND4_X1 port map( A1 => n15494, A2 => n15493, A3 => n15492, A4 => 
                           n15491, ZN => n15495);
   U2635 : AOI22_X1 port map( A1 => n15593, A2 => n15496, B1 => n15591, B2 => 
                           n15495, ZN => n15497);
   U2636 : OAI21_X1 port map( B1 => n15700, B2 => n15498, A => n15497, ZN => 
                           N394);
   U2637 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n15702, B1 => 
                           REGISTERS_25_8_port, B2 => n15701, ZN => n15503);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n15499, B1 => 
                           REGISTERS_30_8_port, B2 => n15713, ZN => n15502);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n15714, B1 => 
                           REGISTERS_20_8_port, B2 => n15705, ZN => n15501);
   U2640 : AOI22_X1 port map( A1 => REGISTERS_26_8_port, A2 => n15716, B1 => 
                           REGISTERS_24_8_port, B2 => n15670, ZN => n15500);
   U2641 : NAND4_X1 port map( A1 => n15503, A2 => n15502, A3 => n15501, A4 => 
                           n15500, ZN => n15509);
   U2642 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n15596, B1 => 
                           REGISTERS_23_8_port, B2 => n15708, ZN => n15507);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n15715, B1 => 
                           REGISTERS_31_8_port, B2 => n15707, ZN => n15506);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_22_8_port, A2 => n15676, B1 => 
                           REGISTERS_17_8_port, B2 => n15717, ZN => n15505);
   U2645 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n15669, B1 => 
                           REGISTERS_18_8_port, B2 => n15677, ZN => n15504);
   U2646 : NAND4_X1 port map( A1 => n15507, A2 => n15506, A3 => n15505, A4 => 
                           n15504, ZN => n15508);
   U2647 : NOR2_X1 port map( A1 => n15509, A2 => n15508, ZN => n15521);
   U2648 : AOI22_X1 port map( A1 => REGISTERS_2_8_port, A2 => n15729, B1 => 
                           REGISTERS_1_8_port, B2 => n15728, ZN => n15513);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_6_8_port, A2 => n15690, B1 => 
                           REGISTERS_0_8_port, B2 => n15637, ZN => n15512);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n15739, B1 => 
                           REGISTERS_4_8_port, B2 => n15560, ZN => n15511);
   U2651 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n15630, B1 => 
                           REGISTERS_3_8_port, B2 => n15740, ZN => n15510);
   U2652 : NAND4_X1 port map( A1 => n15513, A2 => n15512, A3 => n15511, A4 => 
                           n15510, ZN => n15519);
   U2653 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n15630, B1 => 
                           REGISTERS_14_8_port, B2 => n15737, ZN => n15517);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_10_8_port, A2 => n15685, B1 => 
                           REGISTERS_12_8_port, B2 => n15732, ZN => n15516);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n15636, B1 => 
                           REGISTERS_9_8_port, B2 => n15660, ZN => n15515);
   U2656 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n15684, B1 => 
                           REGISTERS_8_8_port, B2 => n15637, ZN => n15514);
   U2657 : NAND4_X1 port map( A1 => n15517, A2 => n15516, A3 => n15515, A4 => 
                           n15514, ZN => n15518);
   U2658 : AOI22_X1 port map( A1 => n15593, A2 => n15519, B1 => n15591, B2 => 
                           n15518, ZN => n15520);
   U2659 : OAI21_X1 port map( B1 => n15755, B2 => n15521, A => n15520, ZN => 
                           N393);
   U2660 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n15719, B1 => 
                           REGISTERS_31_7_port, B2 => n15707, ZN => n15525);
   U2661 : AOI22_X1 port map( A1 => REGISTERS_30_7_port, A2 => n15548, B1 => 
                           REGISTERS_18_7_port, B2 => n15677, ZN => n15524);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n15717, B1 => 
                           REGISTERS_27_7_port, B2 => n15675, ZN => n15523);
   U2663 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n15669, B1 => 
                           REGISTERS_24_7_port, B2 => n15670, ZN => n15522);
   U2664 : NAND4_X1 port map( A1 => n15525, A2 => n15524, A3 => n15523, A4 => 
                           n15522, ZN => n15531);
   U2665 : AOI22_X1 port map( A1 => REGISTERS_19_7_port, A2 => n15715, B1 => 
                           REGISTERS_28_7_port, B2 => n15619, ZN => n15529);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n15701, B1 => 
                           REGISTERS_29_7_port, B2 => n15718, ZN => n15528);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n15676, B1 => 
                           REGISTERS_26_7_port, B2 => n15716, ZN => n15527);
   U2668 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n15705, B1 => 
                           REGISTERS_23_7_port, B2 => n15708, ZN => n15526);
   U2669 : NAND4_X1 port map( A1 => n15529, A2 => n15528, A3 => n15527, A4 => 
                           n15526, ZN => n15530);
   U2670 : NOR2_X1 port map( A1 => n15531, A2 => n15530, ZN => n15543);
   U2671 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n15741, B1 => 
                           REGISTERS_3_7_port, B2 => n15684, ZN => n15535);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n15744, B1 => 
                           REGISTERS_2_7_port, B2 => n15742, ZN => n15534);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n15727, B1 => 
                           REGISTERS_6_7_port, B2 => n15690, ZN => n15533);
   U2674 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n15738, B1 => 
                           REGISTERS_5_7_port, B2 => n15743, ZN => n15532);
   U2675 : NAND4_X1 port map( A1 => n15535, A2 => n15534, A3 => n15533, A4 => 
                           n15532, ZN => n15541);
   U2676 : AOI22_X1 port map( A1 => REGISTERS_10_7_port, A2 => n15742, B1 => 
                           REGISTERS_9_7_port, B2 => n15741, ZN => n15539);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n15738, B1 => 
                           REGISTERS_15_7_port, B2 => n15739, ZN => n15538);
   U2678 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n15684, B1 => 
                           REGISTERS_14_7_port, B2 => n15690, ZN => n15537);
   U2679 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n15630, B1 => 
                           REGISTERS_12_7_port, B2 => n15732, ZN => n15536);
   U2680 : NAND4_X1 port map( A1 => n15539, A2 => n15538, A3 => n15537, A4 => 
                           n15536, ZN => n15540);
   U2681 : AOI22_X1 port map( A1 => n15593, A2 => n15541, B1 => n15591, B2 => 
                           n15540, ZN => n15542);
   U2682 : OAI21_X1 port map( B1 => n15700, B2 => n15543, A => n15542, ZN => 
                           N392);
   U2683 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n15702, B1 => 
                           REGISTERS_17_6_port, B2 => n15717, ZN => n15547);
   U2684 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n15701, B1 => 
                           REGISTERS_23_6_port, B2 => n15708, ZN => n15546);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_31_6_port, A2 => n15575, B1 => 
                           REGISTERS_21_6_port, B2 => n15719, ZN => n15545);
   U2686 : AOI22_X1 port map( A1 => REGISTERS_22_6_port, A2 => n15676, B1 => 
                           REGISTERS_18_6_port, B2 => n15677, ZN => n15544);
   U2687 : NAND4_X1 port map( A1 => n15547, A2 => n15546, A3 => n15545, A4 => 
                           n15544, ZN => n15555);
   U2688 : AOI22_X1 port map( A1 => REGISTERS_30_6_port, A2 => n15548, B1 => 
                           REGISTERS_20_6_port, B2 => n15705, ZN => n15553);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_19_6_port, A2 => n15574, B1 => 
                           REGISTERS_24_6_port, B2 => n15670, ZN => n15552);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n15596, B1 => 
                           REGISTERS_16_6_port, B2 => n15669, ZN => n15551);
   U2691 : AOI22_X1 port map( A1 => REGISTERS_26_6_port, A2 => n15549, B1 => 
                           REGISTERS_27_6_port, B2 => n15675, ZN => n15550);
   U2692 : NAND4_X1 port map( A1 => n15553, A2 => n15552, A3 => n15551, A4 => 
                           n15550, ZN => n15554);
   U2693 : NOR2_X1 port map( A1 => n15555, A2 => n15554, ZN => n15569);
   U2694 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n15630, B1 => 
                           REGISTERS_6_6_port, B2 => n15690, ZN => n15559);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n15560, B1 => 
                           REGISTERS_1_6_port, B2 => n15741, ZN => n15558);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_2_6_port, A2 => n15729, B1 => 
                           REGISTERS_7_6_port, B2 => n15739, ZN => n15557);
   U2697 : AOI22_X1 port map( A1 => REGISTERS_3_6_port, A2 => n15684, B1 => 
                           REGISTERS_0_6_port, B2 => n15637, ZN => n15556);
   U2698 : NAND4_X1 port map( A1 => n15559, A2 => n15558, A3 => n15557, A4 => 
                           n15556, ZN => n15566);
   U2699 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n15660, B1 => 
                           REGISTERS_13_6_port, B2 => n15743, ZN => n15564);
   U2700 : AOI22_X1 port map( A1 => REGISTERS_14_6_port, A2 => n15631, B1 => 
                           REGISTERS_15_6_port, B2 => n15739, ZN => n15563);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n15691, B1 => 
                           REGISTERS_10_6_port, B2 => n15742, ZN => n15562);
   U2702 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n15738, B1 => 
                           REGISTERS_12_6_port, B2 => n15560, ZN => n15561);
   U2703 : NAND4_X1 port map( A1 => n15564, A2 => n15563, A3 => n15562, A4 => 
                           n15561, ZN => n15565);
   U2704 : AOI22_X1 port map( A1 => n15567, A2 => n15566, B1 => n15591, B2 => 
                           n15565, ZN => n15568);
   U2705 : OAI21_X1 port map( B1 => n15755, B2 => n15569, A => n15568, ZN => 
                           N391);
   U2706 : AOI22_X1 port map( A1 => REGISTERS_26_5_port, A2 => n15716, B1 => 
                           REGISTERS_18_5_port, B2 => n15677, ZN => n15573);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n15719, B1 => 
                           REGISTERS_29_5_port, B2 => n15718, ZN => n15572);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n15701, B1 => 
                           REGISTERS_23_5_port, B2 => n15708, ZN => n15571);
   U2709 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n15720, B1 => 
                           REGISTERS_27_5_port, B2 => n15675, ZN => n15570);
   U2710 : NAND4_X1 port map( A1 => n15573, A2 => n15572, A3 => n15571, A4 => 
                           n15570, ZN => n15581);
   U2711 : AOI22_X1 port map( A1 => REGISTERS_19_5_port, A2 => n15574, B1 => 
                           REGISTERS_22_5_port, B2 => n15706, ZN => n15579);
   U2712 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n15669, B1 => 
                           REGISTERS_30_5_port, B2 => n15713, ZN => n15578);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_31_5_port, A2 => n15575, B1 => 
                           REGISTERS_20_5_port, B2 => n15705, ZN => n15577);
   U2714 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n15702, B1 => 
                           REGISTERS_17_5_port, B2 => n15717, ZN => n15576);
   U2715 : NAND4_X1 port map( A1 => n15579, A2 => n15578, A3 => n15577, A4 => 
                           n15576, ZN => n15580);
   U2716 : NOR2_X1 port map( A1 => n15581, A2 => n15580, ZN => n15595);
   U2717 : AOI22_X1 port map( A1 => REGISTERS_6_5_port, A2 => n15737, B1 => 
                           REGISTERS_2_5_port, B2 => n15742, ZN => n15585);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n15741, B1 => 
                           REGISTERS_5_5_port, B2 => n15630, ZN => n15584);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n15744, B1 => 
                           REGISTERS_3_5_port, B2 => n15684, ZN => n15583);
   U2720 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n15738, B1 => 
                           REGISTERS_7_5_port, B2 => n15739, ZN => n15582);
   U2721 : NAND4_X1 port map( A1 => n15585, A2 => n15584, A3 => n15583, A4 => 
                           n15582, ZN => n15592);
   U2722 : AOI22_X1 port map( A1 => REGISTERS_14_5_port, A2 => n15737, B1 => 
                           REGISTERS_11_5_port, B2 => n15684, ZN => n15589);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n15738, B1 => 
                           REGISTERS_12_5_port, B2 => n15732, ZN => n15588);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_10_5_port, A2 => n15685, B1 => 
                           REGISTERS_9_5_port, B2 => n15728, ZN => n15587);
   U2725 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n15636, B1 => 
                           REGISTERS_13_5_port, B2 => n15743, ZN => n15586);
   U2726 : NAND4_X1 port map( A1 => n15589, A2 => n15588, A3 => n15587, A4 => 
                           n15586, ZN => n15590);
   U2727 : AOI22_X1 port map( A1 => n15593, A2 => n15592, B1 => n15591, B2 => 
                           n15590, ZN => n15594);
   U2728 : OAI21_X1 port map( B1 => n15700, B2 => n15595, A => n15594, ZN => 
                           N390);
   U2729 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n15719, B1 => 
                           REGISTERS_28_4_port, B2 => n15619, ZN => n15600);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n15596, B1 => 
                           REGISTERS_19_4_port, B2 => n15715, ZN => n15599);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n15676, B1 => 
                           REGISTERS_18_4_port, B2 => n15677, ZN => n15598);
   U2732 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n15701, B1 => 
                           REGISTERS_16_4_port, B2 => n15669, ZN => n15597);
   U2733 : NAND4_X1 port map( A1 => n15600, A2 => n15599, A3 => n15598, A4 => 
                           n15597, ZN => n15606);
   U2734 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n15717, B1 => 
                           REGISTERS_30_4_port, B2 => n15713, ZN => n15604);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n15670, B1 => 
                           REGISTERS_20_4_port, B2 => n15705, ZN => n15603);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n15714, B1 => 
                           REGISTERS_31_4_port, B2 => n15707, ZN => n15602);
   U2737 : AOI22_X1 port map( A1 => REGISTERS_23_4_port, A2 => n15708, B1 => 
                           REGISTERS_26_4_port, B2 => n15716, ZN => n15601);
   U2738 : NAND4_X1 port map( A1 => n15604, A2 => n15603, A3 => n15602, A4 => 
                           n15601, ZN => n15605);
   U2739 : NOR2_X1 port map( A1 => n15606, A2 => n15605, ZN => n15618);
   U2740 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n15731, B1 => 
                           REGISTERS_6_4_port, B2 => n15737, ZN => n15610);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n15732, B1 => 
                           REGISTERS_0_4_port, B2 => n15730, ZN => n15609);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n15684, B1 => 
                           REGISTERS_7_4_port, B2 => n15739, ZN => n15608);
   U2743 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n15660, B1 => 
                           REGISTERS_2_4_port, B2 => n15742, ZN => n15607);
   U2744 : NAND4_X1 port map( A1 => n15610, A2 => n15609, A3 => n15608, A4 => 
                           n15607, ZN => n15616);
   U2745 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n15741, B1 => 
                           REGISTERS_14_4_port, B2 => n15737, ZN => n15614);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n15738, B1 => 
                           REGISTERS_13_4_port, B2 => n15630, ZN => n15613);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n15739, B1 => 
                           REGISTERS_12_4_port, B2 => n15732, ZN => n15612);
   U2748 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n15684, B1 => 
                           REGISTERS_10_4_port, B2 => n15742, ZN => n15611);
   U2749 : NAND4_X1 port map( A1 => n15614, A2 => n15613, A3 => n15612, A4 => 
                           n15611, ZN => n15615);
   U2750 : AOI22_X1 port map( A1 => n15752, A2 => n15616, B1 => n15750, B2 => 
                           n15615, ZN => n15617);
   U2751 : OAI21_X1 port map( B1 => n15755, B2 => n15618, A => n15617, ZN => 
                           N389);
   U2752 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n15717, B1 => 
                           REGISTERS_22_3_port, B2 => n15706, ZN => n15623);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_31_3_port, A2 => n15707, B1 => 
                           REGISTERS_29_3_port, B2 => n15718, ZN => n15622);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n15719, B1 => 
                           REGISTERS_30_3_port, B2 => n15713, ZN => n15621);
   U2755 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n15720, B1 => 
                           REGISTERS_28_3_port, B2 => n15619, ZN => n15620);
   U2756 : NAND4_X1 port map( A1 => n15623, A2 => n15622, A3 => n15621, A4 => 
                           n15620, ZN => n15629);
   U2757 : AOI22_X1 port map( A1 => REGISTERS_26_3_port, A2 => n15716, B1 => 
                           REGISTERS_27_3_port, B2 => n15675, ZN => n15627);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n15669, B1 => 
                           REGISTERS_20_3_port, B2 => n15705, ZN => n15626);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n15708, B1 => 
                           REGISTERS_19_3_port, B2 => n15715, ZN => n15625);
   U2760 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n15701, B1 => 
                           REGISTERS_18_3_port, B2 => n15677, ZN => n15624);
   U2761 : NAND4_X1 port map( A1 => n15627, A2 => n15626, A3 => n15625, A4 => 
                           n15624, ZN => n15628);
   U2762 : NOR2_X1 port map( A1 => n15629, A2 => n15628, ZN => n15645);
   U2763 : AOI22_X1 port map( A1 => REGISTERS_7_3_port, A2 => n15727, B1 => 
                           REGISTERS_4_3_port, B2 => n15732, ZN => n15635);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n15630, B1 => 
                           REGISTERS_1_3_port, B2 => n15741, ZN => n15634);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n15742, B1 => 
                           REGISTERS_6_3_port, B2 => n15631, ZN => n15633);
   U2766 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n15684, B1 => 
                           REGISTERS_0_3_port, B2 => n15730, ZN => n15632);
   U2767 : NAND4_X1 port map( A1 => n15635, A2 => n15634, A3 => n15633, A4 => 
                           n15632, ZN => n15643);
   U2768 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n15741, B1 => 
                           REGISTERS_14_3_port, B2 => n15737, ZN => n15641);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_15_3_port, A2 => n15636, B1 => 
                           REGISTERS_13_3_port, B2 => n15743, ZN => n15640);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n15740, B1 => 
                           REGISTERS_8_3_port, B2 => n15637, ZN => n15639);
   U2771 : AOI22_X1 port map( A1 => REGISTERS_10_3_port, A2 => n15729, B1 => 
                           REGISTERS_12_3_port, B2 => n15744, ZN => n15638);
   U2772 : NAND4_X1 port map( A1 => n15641, A2 => n15640, A3 => n15639, A4 => 
                           n15638, ZN => n15642);
   U2773 : AOI22_X1 port map( A1 => n15752, A2 => n15643, B1 => n15750, B2 => 
                           n15642, ZN => n15644);
   U2774 : OAI21_X1 port map( B1 => n15700, B2 => n15645, A => n15644, ZN => 
                           N388);
   U2775 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n15714, B1 => 
                           REGISTERS_19_2_port, B2 => n15715, ZN => n15649);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n15669, B1 => 
                           REGISTERS_29_2_port, B2 => n15718, ZN => n15648);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_30_2_port, A2 => n15713, B1 => 
                           REGISTERS_25_2_port, B2 => n15701, ZN => n15647);
   U2778 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n15708, B1 => 
                           REGISTERS_20_2_port, B2 => n15705, ZN => n15646);
   U2779 : NAND4_X1 port map( A1 => n15649, A2 => n15648, A3 => n15647, A4 => 
                           n15646, ZN => n15655);
   U2780 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n15720, B1 => 
                           REGISTERS_26_2_port, B2 => n15716, ZN => n15653);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n15702, B1 => 
                           REGISTERS_21_2_port, B2 => n15719, ZN => n15652);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n15707, B1 => 
                           REGISTERS_22_2_port, B2 => n15706, ZN => n15651);
   U2783 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n15717, B1 => 
                           REGISTERS_18_2_port, B2 => n15677, ZN => n15650);
   U2784 : NAND4_X1 port map( A1 => n15653, A2 => n15652, A3 => n15651, A4 => 
                           n15650, ZN => n15654);
   U2785 : NOR2_X1 port map( A1 => n15655, A2 => n15654, ZN => n15668);
   U2786 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n15739, B1 => 
                           REGISTERS_4_2_port, B2 => n15744, ZN => n15659);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n15738, B1 => 
                           REGISTERS_2_2_port, B2 => n15742, ZN => n15658);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n15731, B1 => 
                           REGISTERS_1_2_port, B2 => n15741, ZN => n15657);
   U2789 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n15691, B1 => 
                           REGISTERS_6_2_port, B2 => n15690, ZN => n15656);
   U2790 : NAND4_X1 port map( A1 => n15659, A2 => n15658, A3 => n15657, A4 => 
                           n15656, ZN => n15666);
   U2791 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n15738, B1 => 
                           REGISTERS_15_2_port, B2 => n15727, ZN => n15664);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n15685, B1 => 
                           REGISTERS_9_2_port, B2 => n15660, ZN => n15663);
   U2793 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n15743, B1 => 
                           REGISTERS_12_2_port, B2 => n15732, ZN => n15662);
   U2794 : AOI22_X1 port map( A1 => REGISTERS_11_2_port, A2 => n15740, B1 => 
                           REGISTERS_14_2_port, B2 => n15737, ZN => n15661);
   U2795 : NAND4_X1 port map( A1 => n15664, A2 => n15663, A3 => n15662, A4 => 
                           n15661, ZN => n15665);
   U2796 : AOI22_X1 port map( A1 => n15752, A2 => n15666, B1 => n15750, B2 => 
                           n15665, ZN => n15667);
   U2797 : OAI21_X1 port map( B1 => n15755, B2 => n15668, A => n15667, ZN => 
                           N387);
   U2798 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n15702, B1 => 
                           REGISTERS_16_1_port, B2 => n15669, ZN => n15674);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n15715, B1 => 
                           REGISTERS_29_1_port, B2 => n15718, ZN => n15673);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_30_1_port, A2 => n15713, B1 => 
                           REGISTERS_24_1_port, B2 => n15670, ZN => n15672);
   U2801 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n15705, B1 => 
                           REGISTERS_31_1_port, B2 => n15707, ZN => n15671);
   U2802 : NAND4_X1 port map( A1 => n15674, A2 => n15673, A3 => n15672, A4 => 
                           n15671, ZN => n15683);
   U2803 : AOI22_X1 port map( A1 => REGISTERS_26_1_port, A2 => n15716, B1 => 
                           REGISTERS_25_1_port, B2 => n15701, ZN => n15681);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_23_1_port, A2 => n15708, B1 => 
                           REGISTERS_27_1_port, B2 => n15675, ZN => n15680);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_22_1_port, A2 => n15676, B1 => 
                           REGISTERS_17_1_port, B2 => n15717, ZN => n15679);
   U2806 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n15677, B1 => 
                           REGISTERS_21_1_port, B2 => n15719, ZN => n15678);
   U2807 : NAND4_X1 port map( A1 => n15681, A2 => n15680, A3 => n15679, A4 => 
                           n15678, ZN => n15682);
   U2808 : NOR2_X1 port map( A1 => n15683, A2 => n15682, ZN => n15699);
   U2809 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n15743, B1 => 
                           REGISTERS_6_1_port, B2 => n15737, ZN => n15689);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n15741, B1 => 
                           REGISTERS_7_1_port, B2 => n15727, ZN => n15688);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_3_1_port, A2 => n15684, B1 => 
                           REGISTERS_0_1_port, B2 => n15730, ZN => n15687);
   U2812 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n15744, B1 => 
                           REGISTERS_2_1_port, B2 => n15685, ZN => n15686);
   U2813 : NAND4_X1 port map( A1 => n15689, A2 => n15688, A3 => n15687, A4 => 
                           n15686, ZN => n15697);
   U2814 : AOI22_X1 port map( A1 => REGISTERS_10_1_port, A2 => n15742, B1 => 
                           REGISTERS_8_1_port, B2 => n15730, ZN => n15695);
   U2815 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n15741, B1 => 
                           REGISTERS_15_1_port, B2 => n15727, ZN => n15694);
   U2816 : AOI22_X1 port map( A1 => REGISTERS_14_1_port, A2 => n15690, B1 => 
                           REGISTERS_12_1_port, B2 => n15744, ZN => n15693);
   U2817 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n15691, B1 => 
                           REGISTERS_13_1_port, B2 => n15743, ZN => n15692);
   U2818 : NAND4_X1 port map( A1 => n15695, A2 => n15694, A3 => n15693, A4 => 
                           n15692, ZN => n15696);
   U2819 : AOI22_X1 port map( A1 => n15752, A2 => n15697, B1 => n15750, B2 => 
                           n15696, ZN => n15698);
   U2820 : OAI21_X1 port map( B1 => n15700, B2 => n15699, A => n15698, ZN => 
                           N386);
   U2821 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n15702, B1 => 
                           REGISTERS_25_0_port, B2 => n15701, ZN => n15712);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_18_0_port, A2 => n15704, B1 => 
                           REGISTERS_16_0_port, B2 => n15703, ZN => n15711);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_22_0_port, A2 => n15706, B1 => 
                           REGISTERS_20_0_port, B2 => n15705, ZN => n15710);
   U2824 : AOI22_X1 port map( A1 => REGISTERS_23_0_port, A2 => n15708, B1 => 
                           REGISTERS_31_0_port, B2 => n15707, ZN => n15709);
   U2825 : NAND4_X1 port map( A1 => n15712, A2 => n15711, A3 => n15710, A4 => 
                           n15709, ZN => n15726);
   U2826 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n15714, B1 => 
                           REGISTERS_30_0_port, B2 => n15713, ZN => n15724);
   U2827 : AOI22_X1 port map( A1 => REGISTERS_26_0_port, A2 => n15716, B1 => 
                           REGISTERS_19_0_port, B2 => n15715, ZN => n15723);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n15718, B1 => 
                           REGISTERS_17_0_port, B2 => n15717, ZN => n15722);
   U2829 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n15720, B1 => 
                           REGISTERS_21_0_port, B2 => n15719, ZN => n15721);
   U2830 : NAND4_X1 port map( A1 => n15724, A2 => n15723, A3 => n15722, A4 => 
                           n15721, ZN => n15725);
   U2831 : NOR2_X1 port map( A1 => n15726, A2 => n15725, ZN => n15754);
   U2832 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n15727, B1 => 
                           REGISTERS_6_0_port, B2 => n15737, ZN => n15736);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n15729, B1 => 
                           REGISTERS_1_0_port, B2 => n15728, ZN => n15735);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_3_0_port, A2 => n15740, B1 => 
                           REGISTERS_0_0_port, B2 => n15730, ZN => n15734);
   U2835 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n15732, B1 => 
                           REGISTERS_5_0_port, B2 => n15731, ZN => n15733);
   U2836 : NAND4_X1 port map( A1 => n15736, A2 => n15735, A3 => n15734, A4 => 
                           n15733, ZN => n15751);
   U2837 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n15738, B1 => 
                           REGISTERS_14_0_port, B2 => n15737, ZN => n15748);
   U2838 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n15740, B1 => 
                           REGISTERS_15_0_port, B2 => n15739, ZN => n15747);
   U2839 : AOI22_X1 port map( A1 => REGISTERS_10_0_port, A2 => n15742, B1 => 
                           REGISTERS_9_0_port, B2 => n15741, ZN => n15746);
   U2840 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n15744, B1 => 
                           REGISTERS_13_0_port, B2 => n15743, ZN => n15745);
   U2841 : NAND4_X1 port map( A1 => n15748, A2 => n15747, A3 => n15746, A4 => 
                           n15745, ZN => n15749);
   U2842 : AOI22_X1 port map( A1 => n15752, A2 => n15751, B1 => n15750, B2 => 
                           n15749, ZN => n15753);
   U2843 : OAI21_X1 port map( B1 => n15755, B2 => n15754, A => n15753, ZN => 
                           N385);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ENABLE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_28_port, 
      curr_instruction_to_cu_i_27_port, curr_instruction_to_cu_i_26_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_5_port, curr_instruction_to_cu_i_4_port, 
      curr_instruction_to_cu_i_3_port, curr_instruction_to_cu_i_2_port, 
      curr_instruction_to_cu_i_1_port, curr_instruction_to_cu_i_0_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n131, cu_i_n127, 
      cu_i_n126, cu_i_n125, cu_i_n124, cu_i_n123, cu_i_n210, cu_i_n209, 
      cu_i_n145, cu_i_n26, cu_i_n25, cu_i_n23, cu_i_cw1_i_4_port, 
      cu_i_cw1_i_7_port, cu_i_cw1_i_8_port, cu_i_cw3_6_port, cu_i_cw2_5_port, 
      cu_i_cw2_6_port, cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_0_port, 
      cu_i_cw1_1_port, cu_i_cw1_2_port, cu_i_cw1_3_port, cu_i_cw1_4_port, 
      cu_i_cw1_5_port, cu_i_cw1_6_port, cu_i_cw1_7_port, cu_i_cw1_8_port, 
      cu_i_cw1_10_port, cu_i_cw1_11_port, cu_i_cw1_12_port, cu_i_N279, 
      cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, 
      cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, 
      cu_i_cmd_word_4_port, cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, 
      cu_i_cmd_word_8_port, cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n78, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_n12, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n309, n311, n691, n697, n699,
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n737, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n756, 
      n758, n759, n760, n761, n762, n763, n764, n1152, n2319, n3092, n3486, 
      n3487, n3488, n3489, n3494, n3495, n3496, n3497, n3498, n3499, n3500, 
      n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
      n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, 
      n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, 
      n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, 
      n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
      n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, 
      n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, 
      n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, 
      n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, 
      n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, 
      n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, 
      n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, 
      n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
      n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, 
      n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, 
      n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, 
      n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, 
      n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, 
      n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, 
      n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, 
      n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, 
      n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, 
      n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, 
      n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, 
      n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, 
      n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, 
      n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, 
      n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, 
      n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, 
      n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, 
      n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, 
      n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, 
      n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, 
      n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, 
      n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, 
      n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
      n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
      n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, 
      n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, 
      n3891, n3892, n3893, DRAM_ENABLE_port, n3895, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => n_1413, QN => cu_i_n123);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n12, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n43, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1414, mul_exeception => 
                           n_1415, FUNC(0) => n3494, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1416, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n3893, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n3893, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n3893, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n309, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n3893, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n3893, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n3893, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n309, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n3893, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n3893, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n309, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n3893, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n3893, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n3893, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n3893, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n3893, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n309, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n3893, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n3893, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n3893, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n309, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n309, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n309, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n309, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n3893, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n3893, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n3893, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n3893, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n309, Z =>
                           DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n3893, Z 
                           => DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n3895, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n3895, Z =>
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n3895, Z =>
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n3895, Z =>
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n3895, Z =>
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n3895, Z =>
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n3895, Z =>
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n3895, Z =>
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n3895, Z =>
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n3895, Z =>
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n3895, Z =>
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n3895, Z =>
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => n3895, Z =>
                           DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => n3895, Z =>
                           DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => n3895, Z =>
                           DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => n3895, Z =>
                           DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => n3895, Z => 
                           DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1417);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n3891, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n3892, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n3892, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n3892, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n3891, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n3892, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n3891, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n3892, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n3890, D => datapath_i_n18, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n3890, D => datapath_i_n17, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n3890, D => datapath_i_n16, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n3890, D => datapath_i_n15, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n3890, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n3890, D => 
                           curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n3890, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n3890, D => datapath_i_n12, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n3890, D => datapath_i_n11, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n3890, D => datapath_i_n10, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n3890, D => datapath_i_n9, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n3495, CK => CLK, RN => RST
                           , Q => cu_i_cw3_6_port, QN => n_1418);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n131, CK => CLK, RN =>
                           RST, Q => n_1419, QN => n699);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1420);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1421);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1422);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n126, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n3889);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => n_1423, QN => n756);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n3892, CK => CLK, RN => RST
                           , Q => n_1424, QN => n2319);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1425)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1426)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1427)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1428);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1429);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n311, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1430);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1431);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => n1152, CK => CLK, RN => RST,
                           Q => cu_i_cw1_4_port, QN => n_1432);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1433);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1434);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1435);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1436);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1437);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1438);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1439);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1440);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1441);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1442);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1443);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1444);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1445);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1446);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1447);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1448);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1449);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1450);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1451);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1452);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1453);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1454);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1455);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1456);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1457);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1458);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1459);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1460);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1461);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1462);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1463);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1464);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1465);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1466);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1467);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1468)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1469)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1470)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1471)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1472)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1473)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1474)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1475)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1476)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1477)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1478)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1479)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1480)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1481)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1482)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1483)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1484)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1485)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1486)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1487)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1488)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1489)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1490);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1491);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1492);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1493);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1494);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1495);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1496);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1497);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1498);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1499);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1500);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1501);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1502);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1503);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1504);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1505);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1506);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1507);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1508);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1509);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1510);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1511);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1512);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1513);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1514);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1515);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1516);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1517);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1518);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1519);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1520);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1521);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1522);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1523);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1524);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1525);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1526);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1527);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1528);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1529);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1530);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1531);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1532);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1533);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1534);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1535);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1536);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1537);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1538);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1539);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1540);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1541);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1542);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1543);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1544);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1545);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1546);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1547);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1548);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1549);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1550);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1551);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1552);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1553);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1554);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1555);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1556);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1557);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1558);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1559);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1560);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1561);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1562);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1563);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1564, QN => n703);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1565, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1566, QN => n726);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1567, QN => n725);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1568, QN => n724);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1569, QN => n691);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1570, QN => n723);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1571, QN => n722);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1572, QN => n721);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1573, QN => n720);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1574, QN => n719);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1575, QN => n718);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1576, QN => n717);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1577, QN => n716);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1578, QN => n715);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1579, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1580, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1581, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1582, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1583, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1584, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1585, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1586, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1587, QN => n706);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1588, QN => n705);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1589, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1590, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1591, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1592, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1593, QN => n728);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1594, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1595, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1596);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1597);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1598);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1599);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1600);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1601);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1602);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1603);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1604);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1605);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1606);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1607);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1608);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1609);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1610);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1611);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1612);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1613);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1614);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1615);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1616);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1617);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1618);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1619);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1620);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1621);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1622);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1623);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1624);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1625);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1626);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1627);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n3890, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1628);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1629);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1630);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1631);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1632);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1633);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1634);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1635);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1636);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1637);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1638);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1639);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1640);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1641);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1642);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1643);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1644);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1645);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1646);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1647);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1648);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1649);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1650);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1651);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1652);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1653);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1654);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n764);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n763);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n762);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n761);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n760);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n759);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n758);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1655);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1656);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1657);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1658);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1659);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1660);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1661);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1662);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1663);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1664);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1665);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1666);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1667);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1668);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1669);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1670);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1671);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1672);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1673);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1674);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1675);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1676);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1677);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1678);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1679);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1680);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1681);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1682);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1683);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1684);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1685);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1686);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1687);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1688);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1689);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1690);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1691);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1692);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1693);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1694);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1695);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1696);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1697);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1698);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1699);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1700);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1701);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1702);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1703);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1704);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1705);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1706);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1707);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1708);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1709);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1710);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1711);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1712);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1713);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1714);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1715);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1716);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1717);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1718);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1719);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1720);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1721);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => n3489, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1722);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => n3488, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1723);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1724);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => n3487, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1725);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n3486, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1726);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n3880);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n3875);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => n3882, QN => n737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n3871);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n3883);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n3873);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1727);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1728);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1729);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1730);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1731);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1732);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1733);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n697);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1734);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1735);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1736);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1738);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1741);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1742);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1743);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1744);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n_1745);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n3877);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n3884);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n3872);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n3887);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n3876);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1746
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1747
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1748
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1749
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1750
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1751
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1752
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1753
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1754
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1755
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1756
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1757
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1758
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1759
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1760
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1761
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1762
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1763
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1764
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1765
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1766
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1767
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1768)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1769)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1770)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1771)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1772)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1773)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1774)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1775)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1776)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1777)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1778);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_30_port, QN => 
                           n_1779);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n753);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_28_port, QN => 
                           n_1780);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n751);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_26_port, QN => 
                           n_1781);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n750);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_24_port, QN => 
                           n_1782);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n749);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_22_port, QN => 
                           n_1783);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n748);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_20_port, QN => 
                           n_1784);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n747);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_18_port, QN => 
                           n_1785);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n746);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_16_port, QN => 
                           n_1786);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n745);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_14_port, QN => 
                           n_1787);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n752);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_12_port, QN => 
                           n_1788);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n744);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_10_port, QN => 
                           n_1789);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n743
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_8_port, QN => 
                           n_1790);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n742
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_6_port, QN => 
                           n_1791);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n741
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_1792);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_1793);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_1794);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1795);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1796);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => n3878, QN => n3092);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1797);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => n3881, QN => cu_i_n26);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => n3888, QN => cu_i_n25);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => n3885, QN => cu_i_n124);
   U3283 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   U3284 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(8), ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U3285 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U3286 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U3287 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U3288 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U3289 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U3290 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(31), ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U3291 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(30), ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U3292 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U3293 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(29), ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U3294 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(28), ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U3295 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(27), ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U3296 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(26), ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U3297 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(25), ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U3298 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(24), ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U3299 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(23), ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U3300 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(22), ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U3301 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(21), ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U3302 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U3303 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U3304 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U3305 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U3306 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U3307 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U3308 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(15), ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U3309 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(14), ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U3310 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(13), ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U3311 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(12), ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U3312 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(11), ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U3313 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(10), ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U3314 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(0), ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => n3874, QN => cu_i_n125);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => n3886, QN => cu_i_n23);
   cu_i_stall_reg : DFFR_X2 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n704, QN => n3879);
   U3315 : NAND2_X1 port map( A1 => n3523, A2 => n3885, ZN => n3631);
   U3316 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n3880, A3 => n3873, A4 => n3636, ZN => 
                           cu_i_cmd_word_4_port);
   U3317 : AOI21_X1 port map( B1 => n3762, B2 => n3761, A => cu_i_cw3_6_port, 
                           ZN => n3763);
   U3318 : OAI21_X1 port map( B1 => n3631, B2 => n3632, A => n699, ZN => 
                           write_rf_i);
   U3319 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_0_port, B1
                           => cu_i_cw1_0_port, B2 => n3879, ZN => n3587);
   U3320 : NAND2_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, ZN => n3523);
   U3321 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U3322 : NOR2_X1 port map( A1 => n3587, A2 => n3581, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U3323 : AOI211_X1 port map( C1 => n3568, C2 => n3639, A => 
                           cu_i_cmd_word_4_port, B => cu_i_cmd_word_7_port, ZN 
                           => n3583);
   U3324 : NOR2_X1 port map( A1 => cu_i_n123, A2 => n3886, ZN => n3568);
   U3325 : CLKBUF_X1 port map( A => n3870, Z => n3859);
   U3326 : CLKBUF_X1 port map( A => n3750, Z => n3576);
   U3327 : NAND2_X1 port map( A1 => n3092, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n3750);
   U3328 : CLKBUF_X1 port map( A => n3708, Z => n3756);
   U3329 : AOI21_X1 port map( B1 => n3569, B2 => n3584, A => n3596, ZN => n3759
                           );
   U3330 : NOR4_X1 port map( A1 => n3612, A2 => n3599, A3 => n3872, A4 => n3877
                           , ZN => n3584);
   U3331 : OR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n3522
                           , A3 => n3883, ZN => n3802);
   U3332 : NAND3_X1 port map( A1 => n3568, A2 => 
                           curr_instruction_to_cu_i_27_port, A3 => n3871, ZN =>
                           n3636);
   U3333 : OAI22_X1 port map( A1 => n3879, A2 => cu_i_cmd_word_4_port, B1 => 
                           cu_i_cw2_8_port, B2 => n704, ZN => n309);
   U3334 : INV_X1 port map( A => n309, ZN => DRAM_ENABLE_port);
   U3335 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n3893);
   U3336 : INV_X1 port map( A => cu_i_cmd_word_4_port, ZN => n3757);
   U3337 : NOR2_X1 port map( A1 => n3882, A2 => n3757, ZN => 
                           cu_i_cmd_word_3_port);
   U3338 : OAI22_X1 port map( A1 => n3879, A2 => cu_i_cmd_word_3_port, B1 => 
                           cu_i_cw2_7_port, B2 => n704, ZN => n3585);
   U3339 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n3585, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U3340 : CLKBUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n3895);
   U3341 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n3878, ZN => n3748);
   U3342 : CLKBUF_X1 port map( A => n3748, Z => n3574);
   U3343 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_27_port,
                           B2 => n3878, ZN => n3496);
   U3344 : OAI21_X1 port map( B1 => n724, B2 => n3750, A => n3496, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U3345 : CLKBUF_X1 port map( A => n3878, Z => n3747);
   U3346 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_25_port,
                           B2 => n3747, ZN => n3497);
   U3347 : OAI21_X1 port map( B1 => n723, B2 => n3576, A => n3497, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U3348 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_23_port,
                           B2 => n3878, ZN => n3498);
   U3349 : OAI21_X1 port map( B1 => n721, B2 => n3750, A => n3498, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U3350 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_21_port,
                           B2 => n3747, ZN => n3499);
   U3351 : OAI21_X1 port map( B1 => n719, B2 => n3576, A => n3499, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U3352 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_19_port,
                           B2 => n3878, ZN => n3500);
   U3353 : OAI21_X1 port map( B1 => n717, B2 => n3750, A => n3500, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U3354 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_17_port,
                           B2 => n3747, ZN => n3501);
   U3355 : OAI21_X1 port map( B1 => n715, B2 => n3576, A => n3501, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U3356 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_15_port,
                           B2 => n3878, ZN => n3502);
   U3357 : OAI21_X1 port map( B1 => n713, B2 => n3750, A => n3502, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U3358 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_13_port,
                           B2 => n3747, ZN => n3503);
   U3359 : OAI21_X1 port map( B1 => n711, B2 => n3576, A => n3503, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U3360 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_11_port,
                           B2 => n3878, ZN => n3504);
   U3361 : OAI21_X1 port map( B1 => n709, B2 => n3750, A => n3504, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U3362 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_9_port, 
                           B2 => n3878, ZN => n3505);
   U3363 : OAI21_X1 port map( B1 => n707, B2 => n3750, A => n3505, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U3364 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_7_port, 
                           B2 => n3747, ZN => n3506);
   U3365 : OAI21_X1 port map( B1 => n705, B2 => n3750, A => n3506, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U3366 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_5_port, 
                           B2 => n3878, ZN => n3507);
   U3367 : OAI21_X1 port map( B1 => n731, B2 => n3576, A => n3507, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U3368 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_4_port, 
                           B2 => n3747, ZN => n3508);
   U3369 : OAI21_X1 port map( B1 => n730, B2 => n3576, A => n3508, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U3370 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_2_port, 
                           B2 => n3878, ZN => n3509);
   U3371 : OAI21_X1 port map( B1 => n728, B2 => n3576, A => n3509, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U3372 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_3_port, 
                           B2 => n3747, ZN => n3510);
   U3373 : OAI21_X1 port map( B1 => n729, B2 => n3576, A => n3510, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U3374 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_6_port, 
                           B2 => n3878, ZN => n3511);
   U3375 : OAI21_X1 port map( B1 => n732, B2 => n3576, A => n3511, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U3376 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_8_port, 
                           B2 => n3878, ZN => n3512);
   U3377 : OAI21_X1 port map( B1 => n706, B2 => n3576, A => n3512, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U3378 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_10_port,
                           B2 => n3878, ZN => n3513);
   U3379 : OAI21_X1 port map( B1 => n708, B2 => n3576, A => n3513, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U3380 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_12_port,
                           B2 => n3878, ZN => n3514);
   U3381 : OAI21_X1 port map( B1 => n710, B2 => n3576, A => n3514, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U3382 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_14_port,
                           B2 => n3878, ZN => n3515);
   U3383 : OAI21_X1 port map( B1 => n712, B2 => n3576, A => n3515, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U3384 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_16_port,
                           B2 => n3878, ZN => n3516);
   U3385 : OAI21_X1 port map( B1 => n714, B2 => n3576, A => n3516, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U3386 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_18_port,
                           B2 => n3878, ZN => n3517);
   U3387 : OAI21_X1 port map( B1 => n716, B2 => n3576, A => n3517, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U3388 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_20_port,
                           B2 => n3747, ZN => n3518);
   U3389 : OAI21_X1 port map( B1 => n718, B2 => n3576, A => n3518, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U3390 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_22_port,
                           B2 => n3747, ZN => n3519);
   U3391 : OAI21_X1 port map( B1 => n720, B2 => n3750, A => n3519, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U3392 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_24_port,
                           B2 => n3747, ZN => n3520);
   U3393 : OAI21_X1 port map( B1 => n722, B2 => n3750, A => n3520, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U3394 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_26_port,
                           B2 => n3747, ZN => n3521);
   U3395 : OAI21_X1 port map( B1 => n691, B2 => n3750, A => n3521, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U3396 : NAND4_X1 port map( A1 => n737, A2 => n3568, A3 => n3880, A4 => n3875
                           , ZN => n3522);
   U3397 : NOR2_X1 port map( A1 => n3871, A2 => 
                           curr_instruction_to_cu_i_27_port, ZN => n3616);
   U3398 : INV_X1 port map( A => n3616, ZN => n3608);
   U3399 : OR2_X1 port map( A1 => n3522, A2 => n3608, ZN => n3803);
   U3400 : NAND2_X1 port map( A1 => n3802, A2 => n3803, ZN => n1152);
   U3401 : NAND4_X1 port map( A1 => cu_i_n26, A2 => cu_i_n25, A3 => n3874, A4 
                           => n3885, ZN => cu_i_n145);
   U3402 : NAND2_X1 port map( A1 => cu_i_n145, A2 => n3631, ZN => n3569);
   U3403 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_5_port, A2 => 
                           curr_instruction_to_cu_i_1_port, ZN => n3612);
   U3404 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_0_port, ZN => n3599);
   U3405 : NAND3_X1 port map( A1 => n737, A2 => n3880, A3 => n3873, ZN => n3567
                           );
   U3406 : NOR4_X2 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           curr_instruction_to_cu_i_28_port, A3 => 
                           curr_instruction_to_cu_i_27_port, A4 => n3567, ZN =>
                           n3644);
   U3407 : NAND2_X1 port map( A1 => n3584, A2 => n3644, ZN => n3606);
   U3408 : OAI21_X1 port map( B1 => n3569, B2 => n3606, A => n3568, ZN => n3524
                           );
   U3409 : NAND2_X1 port map( A1 => cu_i_n123, A2 => n3886, ZN => n3648);
   U3410 : AOI21_X1 port map( B1 => n3524, B2 => n3648, A => n704, ZN => 
                           IRAM_ENABLE_port);
   U3411 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, 
                           ZN => n3525);
   U3412 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, 
                           ZN => n3528);
   U3413 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, 
                           ZN => n3531);
   U3414 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, 
                           ZN => n3534);
   U3415 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, 
                           ZN => n3537);
   U3416 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, 
                           ZN => n3540);
   U3417 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, 
                           ZN => n3543);
   U3418 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, 
                           ZN => n3546);
   U3419 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, 
                           ZN => n3549);
   U3420 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN
                           => n3552);
   U3421 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN
                           => n3555);
   U3422 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN
                           => n3558);
   U3423 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_3_port, ZN =>
                           n3663);
   U3424 : NOR2_X1 port map( A1 => n3558, A2 => n3663, ZN => n3670);
   U3425 : NAND2_X1 port map( A1 => n3670, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n3669);
   U3426 : NOR2_X1 port map( A1 => n3555, A2 => n3669, ZN => n3676);
   U3427 : NAND2_X1 port map( A1 => n3676, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n3675);
   U3428 : NOR2_X1 port map( A1 => n3552, A2 => n3675, ZN => n3682);
   U3429 : NAND2_X1 port map( A1 => n3682, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n3681);
   U3430 : NOR2_X1 port map( A1 => n3549, A2 => n3681, ZN => n3688);
   U3431 : NAND2_X1 port map( A1 => n3688, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n3687);
   U3432 : NOR2_X1 port map( A1 => n3546, A2 => n3687, ZN => n3694);
   U3433 : NAND2_X1 port map( A1 => n3694, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n3693);
   U3434 : NOR2_X1 port map( A1 => n3543, A2 => n3693, ZN => n3700);
   U3435 : NAND2_X1 port map( A1 => n3700, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n3699);
   U3436 : NOR2_X1 port map( A1 => n3540, A2 => n3699, ZN => n3706);
   U3437 : NAND2_X1 port map( A1 => n3706, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n3705);
   U3438 : NOR2_X1 port map( A1 => n3537, A2 => n3705, ZN => n3713);
   U3439 : NAND2_X1 port map( A1 => n3713, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n3712);
   U3440 : NOR2_X1 port map( A1 => n3534, A2 => n3712, ZN => n3719);
   U3441 : NAND2_X1 port map( A1 => n3719, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n3718);
   U3442 : NOR2_X1 port map( A1 => n3531, A2 => n3718, ZN => n3725);
   U3443 : NAND2_X1 port map( A1 => n3725, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n3724);
   U3444 : NOR2_X1 port map( A1 => n3528, A2 => n3724, ZN => n3731);
   U3445 : NAND2_X1 port map( A1 => n3731, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n3730);
   U3446 : INV_X1 port map( A => n1152, ZN => n3649);
   U3447 : OAI221_X1 port map( B1 => n3879, B2 => n3649, C1 => n704, C2 => n756
                           , A => n3092, ZN => n3660);
   U3448 : INV_X1 port map( A => n3660, ZN => n3708);
   U3449 : NOR2_X1 port map( A1 => n3525, A2 => n3730, ZN => n3737);
   U3450 : AOI211_X1 port map( C1 => n3525, C2 => n3730, A => n3756, B => n3737
                           , ZN => n3527);
   U3451 : NAND2_X1 port map( A1 => IRAM_ENABLE_port, A2 => IRAM_ADDRESS_2_port
                           , ZN => n3657);
   U3452 : INV_X1 port map( A => n3657, ZN => n3659);
   U3453 : AND2_X1 port map( A1 => n3659, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n3666);
   U3454 : NAND2_X1 port map( A1 => n3666, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n3665);
   U3455 : NOR2_X1 port map( A1 => n741, A2 => n3665, ZN => n3672);
   U3456 : NAND2_X1 port map( A1 => n3672, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n3671);
   U3457 : NOR2_X1 port map( A1 => n742, A2 => n3671, ZN => n3678);
   U3458 : NAND2_X1 port map( A1 => n3678, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n3677);
   U3459 : NOR2_X1 port map( A1 => n743, A2 => n3677, ZN => n3684);
   U3460 : NAND2_X1 port map( A1 => n3684, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n3683);
   U3461 : NOR2_X1 port map( A1 => n744, A2 => n3683, ZN => n3690);
   U3462 : NAND2_X1 port map( A1 => n3690, A2 => IRAM_ADDRESS_12_port, ZN => 
                           n3689);
   U3463 : NOR2_X1 port map( A1 => n752, A2 => n3689, ZN => n3696);
   U3464 : NAND2_X1 port map( A1 => n3696, A2 => IRAM_ADDRESS_14_port, ZN => 
                           n3695);
   U3465 : NOR2_X1 port map( A1 => n745, A2 => n3695, ZN => n3702);
   U3466 : NAND2_X1 port map( A1 => n3702, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n3701);
   U3467 : NOR2_X1 port map( A1 => n746, A2 => n3701, ZN => n3709);
   U3468 : NAND2_X1 port map( A1 => n3709, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n3707);
   U3469 : NOR2_X1 port map( A1 => n747, A2 => n3707, ZN => n3715);
   U3470 : NAND2_X1 port map( A1 => n3715, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n3714);
   U3471 : NOR2_X1 port map( A1 => n748, A2 => n3714, ZN => n3721);
   U3472 : NAND2_X1 port map( A1 => n3721, A2 => IRAM_ADDRESS_22_port, ZN => 
                           n3720);
   U3473 : NOR2_X1 port map( A1 => n749, A2 => n3720, ZN => n3727);
   U3474 : NAND2_X1 port map( A1 => n3727, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n3726);
   U3475 : NOR2_X1 port map( A1 => n750, A2 => n3726, ZN => n3733);
   U3476 : NAND2_X1 port map( A1 => n3733, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n3732);
   U3477 : NOR2_X1 port map( A1 => n751, A2 => n3732, ZN => n3739);
   U3478 : AOI211_X1 port map( C1 => n751, C2 => n3732, A => n3739, B => n3660,
                           ZN => n3526);
   U3479 : OR2_X1 port map( A1 => n3527, A2 => n3526, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U3480 : AOI211_X1 port map( C1 => n3528, C2 => n3724, A => n3708, B => n3731
                           , ZN => n3530);
   U3481 : INV_X1 port map( A => n3756, ZN => n3753);
   U3482 : AOI211_X1 port map( C1 => n750, C2 => n3726, A => n3733, B => n3753,
                           ZN => n3529);
   U3483 : OR2_X1 port map( A1 => n3530, A2 => n3529, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U3484 : AOI211_X1 port map( C1 => n3531, C2 => n3718, A => n3708, B => n3725
                           , ZN => n3533);
   U3485 : AOI211_X1 port map( C1 => n749, C2 => n3720, A => n3727, B => n3753,
                           ZN => n3532);
   U3486 : OR2_X1 port map( A1 => n3533, A2 => n3532, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U3487 : AOI211_X1 port map( C1 => n3534, C2 => n3712, A => n3708, B => n3719
                           , ZN => n3536);
   U3488 : AOI211_X1 port map( C1 => n748, C2 => n3714, A => n3721, B => n3753,
                           ZN => n3535);
   U3489 : OR2_X1 port map( A1 => n3536, A2 => n3535, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U3490 : AOI211_X1 port map( C1 => n3537, C2 => n3705, A => n3708, B => n3713
                           , ZN => n3539);
   U3491 : AOI211_X1 port map( C1 => n747, C2 => n3707, A => n3715, B => n3753,
                           ZN => n3538);
   U3492 : OR2_X1 port map( A1 => n3539, A2 => n3538, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U3493 : AOI211_X1 port map( C1 => n3540, C2 => n3699, A => n3708, B => n3706
                           , ZN => n3542);
   U3494 : AOI211_X1 port map( C1 => n746, C2 => n3701, A => n3709, B => n3660,
                           ZN => n3541);
   U3495 : OR2_X1 port map( A1 => n3542, A2 => n3541, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U3496 : AOI211_X1 port map( C1 => n3543, C2 => n3693, A => n3756, B => n3700
                           , ZN => n3545);
   U3497 : AOI211_X1 port map( C1 => n745, C2 => n3695, A => n3702, B => n3660,
                           ZN => n3544);
   U3498 : OR2_X1 port map( A1 => n3545, A2 => n3544, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U3499 : AOI211_X1 port map( C1 => n3546, C2 => n3687, A => n3756, B => n3694
                           , ZN => n3548);
   U3500 : AOI211_X1 port map( C1 => n752, C2 => n3689, A => n3696, B => n3660,
                           ZN => n3547);
   U3501 : OR2_X1 port map( A1 => n3548, A2 => n3547, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U3502 : AOI211_X1 port map( C1 => n3549, C2 => n3681, A => n3756, B => n3688
                           , ZN => n3551);
   U3503 : AOI211_X1 port map( C1 => n744, C2 => n3683, A => n3690, B => n3753,
                           ZN => n3550);
   U3504 : OR2_X1 port map( A1 => n3551, A2 => n3550, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U3505 : AOI211_X1 port map( C1 => n3552, C2 => n3675, A => n3708, B => n3682
                           , ZN => n3554);
   U3506 : AOI211_X1 port map( C1 => n743, C2 => n3677, A => n3684, B => n3753,
                           ZN => n3553);
   U3507 : OR2_X1 port map( A1 => n3554, A2 => n3553, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U3508 : AOI211_X1 port map( C1 => n3555, C2 => n3669, A => n3708, B => n3676
                           , ZN => n3557);
   U3509 : AOI211_X1 port map( C1 => n742, C2 => n3671, A => n3678, B => n3660,
                           ZN => n3556);
   U3510 : OR2_X1 port map( A1 => n3557, A2 => n3556, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U3511 : AOI211_X1 port map( C1 => n3558, C2 => n3663, A => n3708, B => n3670
                           , ZN => n3560);
   U3512 : AOI211_X1 port map( C1 => n741, C2 => n3665, A => n3672, B => n3753,
                           ZN => n3559);
   U3513 : OR2_X1 port map( A1 => n3560, A2 => n3559, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U3514 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => n737
                           , A3 => curr_instruction_to_cu_i_27_port, ZN => 
                           n3561);
   U3515 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n3561, ZN => n3600);
   U3516 : AOI21_X1 port map( B1 => n3871, B2 => n3873, A => n3600, ZN => n3566
                           );
   U3517 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_5_port, A2 => 
                           n3644, A3 => n3877, A4 => n3887, ZN => n3613);
   U3518 : AOI211_X1 port map( C1 => n3876, C2 => n3872, A => n3884, B => n3613
                           , ZN => n3562);
   U3519 : OR2_X1 port map( A1 => n3566, A2 => n3562, ZN => cu_i_N267);
   U3520 : OAI22_X1 port map( A1 => n3879, A2 => cu_i_cw3_6_port, B1 => 
                           cu_i_cw2_6_port, B2 => n704, ZN => n3563);
   U3521 : INV_X1 port map( A => n3563, ZN => n3495);
   U3522 : NAND2_X1 port map( A1 => n3568, A2 => n3644, ZN => n3596);
   U3523 : INV_X1 port map( A => n3568, ZN => n3650);
   U3524 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => n737
                           , ZN => n3615);
   U3525 : NAND2_X1 port map( A1 => n3615, A2 => n3875, ZN => n3564);
   U3526 : NOR2_X1 port map( A1 => n3608, A2 => n3564, ZN => n3623);
   U3527 : OR2_X1 port map( A1 => n3564, A2 => curr_instruction_to_cu_i_26_port
                           , ZN => n3637);
   U3528 : NOR3_X1 port map( A1 => n3875, A2 => n3871, A3 => n3567, ZN => n3622
                           );
   U3529 : INV_X1 port map( A => n3622, ZN => n3565);
   U3530 : NAND2_X1 port map( A1 => n3637, A2 => n3565, ZN => n3614);
   U3531 : NOR3_X1 port map( A1 => n3623, A2 => n3566, A3 => n3614, ZN => n3641
                           );
   U3532 : OAI222_X1 port map( A1 => n3873, A2 => n3802, B1 => n3596, B2 => 
                           n3584, C1 => n3650, C2 => n3641, ZN => n311);
   U3533 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n311, ZN => 
                           cu_i_cmd_word_1_port);
   U3534 : NOR2_X1 port map( A1 => n3803, A2 => n3873, ZN => 
                           cu_i_cmd_word_7_port);
   U3535 : OAI21_X1 port map( B1 => n3608, B2 => n3567, A => n3641, ZN => n3639
                           );
   U3536 : AND2_X1 port map( A1 => n3583, A2 => n3802, ZN => n3828);
   U3537 : INV_X1 port map( A => n3828, ZN => n3891);
   U3538 : INV_X1 port map( A => n3802, ZN => n3890);
   U3539 : INV_X1 port map( A => n3759, ZN => n3758);
   U3540 : AOI221_X1 port map( B1 => n3758, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n3759, C2 =>
                           curr_instruction_to_cu_i_15_port, A => n3890, ZN => 
                           n3570);
   U3541 : INV_X1 port map( A => n3570, ZN => n3489);
   U3542 : AOI221_X1 port map( B1 => n3758, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n3759, C2 =>
                           curr_instruction_to_cu_i_14_port, A => n3890, ZN => 
                           n3571);
   U3543 : INV_X1 port map( A => n3571, ZN => n3488);
   U3544 : AOI221_X1 port map( B1 => n3758, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n3759, C2 =>
                           curr_instruction_to_cu_i_12_port, A => n3890, ZN => 
                           n3572);
   U3545 : INV_X1 port map( A => n3572, ZN => n3487);
   U3546 : AOI221_X1 port map( B1 => n3758, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n3759, C2 =>
                           curr_instruction_to_cu_i_11_port, A => n3890, ZN => 
                           n3573);
   U3547 : INV_X1 port map( A => n3573, ZN => n3486);
   U3548 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n3574, B1 => datapath_i_alu_output_val_i_29_port,
                           B2 => n3747, ZN => n3575);
   U3549 : OAI21_X1 port map( B1 => n726, B2 => n3576, A => n3575, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U3550 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_28_port,
                           B2 => n3747, ZN => n3577);
   U3551 : OAI21_X1 port map( B1 => n725, B2 => n3750, A => n3577, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U3552 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, 
                           ZN => n3578);
   U3553 : NAND2_X1 port map( A1 => n3737, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n3736);
   U3554 : NOR2_X1 port map( A1 => n3578, A2 => n3736, ZN => n3743);
   U3555 : AOI211_X1 port map( C1 => n3578, C2 => n3736, A => n3708, B => n3743
                           , ZN => n3580);
   U3556 : NAND2_X1 port map( A1 => n3739, A2 => IRAM_ADDRESS_28_port, ZN => 
                           n3738);
   U3557 : NOR2_X1 port map( A1 => n753, A2 => n3738, ZN => n3744);
   U3558 : AOI211_X1 port map( C1 => n753, C2 => n3738, A => n3744, B => n3660,
                           ZN => n3579);
   U3559 : OR2_X1 port map( A1 => n3580, A2 => n3579, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U3560 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_2_port, B1
                           => cu_i_cw1_2_port, B2 => n3879, ZN => n3595);
   U3561 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_1_port, B1
                           => cu_i_cw1_1_port, B2 => n3879, ZN => n3589);
   U3562 : INV_X1 port map( A => n704, ZN => n3654);
   U3563 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_3_port, B1
                           => cu_i_cw1_3_port, B2 => n3654, ZN => n3586);
   U3564 : AOI21_X1 port map( B1 => n3595, B2 => n3589, A => n3586, ZN => n3581
                           );
   U3565 : INV_X1 port map( A => n3586, ZN => n3594);
   U3566 : OAI211_X1 port map( C1 => n3587, C2 => n3589, A => n3594, B => n3595
                           , ZN => n3582);
   U3567 : INV_X1 port map( A => n3582, ZN => n3494);
   U3568 : NAND2_X1 port map( A1 => n3583, A2 => n3758, ZN => enable_rf_i);
   U3569 : INV_X1 port map( A => n3596, ZN => n3634);
   U3570 : NAND2_X1 port map( A1 => n3584, A2 => n3634, ZN => n3632);
   U3571 : INV_X1 port map( A => n3828, ZN => n3892);
   U3572 : AND2_X1 port map( A1 => n3892, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U3573 : INV_X1 port map( A => n3585, ZN => DRAM_READNOTWRITE);
   U3574 : AOI22_X1 port map( A1 => n704, A2 => n3828, B1 => n2319, B2 => n3654
                           , ZN => n3831);
   U3575 : CLKBUF_X1 port map( A => n3831, Z => n3833);
   U3576 : MUX2_X1 port map( A => datapath_i_val_b_i_2_port, B => 
                           datapath_i_val_immediate_i_2_port, S => n3833, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U3577 : MUX2_X1 port map( A => datapath_i_val_b_i_0_port, B => 
                           datapath_i_val_immediate_i_0_port, S => n3833, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U3578 : AOI21_X1 port map( B1 => n3595, B2 => n3587, A => n3586, ZN => n3588
                           );
   U3579 : NOR2_X1 port map( A1 => n3589, A2 => n3588, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U3580 : NOR2_X1 port map( A1 => n3874, A2 => n3632, ZN => cu_i_N273);
   U3581 : INV_X1 port map( A => n3632, ZN => n3761);
   U3582 : AOI221_X1 port map( B1 => cu_i_n25, B2 => n3761, C1 => cu_i_n26, C2 
                           => n3761, A => cu_i_N273, ZN => n3590);
   U3583 : INV_X1 port map( A => n3590, ZN => n3593);
   U3584 : NOR2_X1 port map( A1 => cu_i_n125, A2 => n3632, ZN => n3591);
   U3585 : NAND2_X1 port map( A1 => n3591, A2 => n3881, ZN => n3630);
   U3586 : NOR2_X1 port map( A1 => cu_i_n25, A2 => n3630, ZN => n3592);
   U3587 : MUX2_X1 port map( A => n3593, B => n3592, S => cu_i_n124, Z => 
                           cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U3589 : MUX2_X1 port map( A => datapath_i_val_b_i_1_port, B => 
                           datapath_i_val_immediate_i_1_port, S => n3831, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U3590 : NOR2_X1 port map( A1 => n3595, A2 => n3594, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U3591 : NAND2_X1 port map( A1 => n3828, A2 => n3596, ZN => cu_i_N278);
   U3592 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_4_port, ZN => n3597);
   U3593 : NAND2_X1 port map( A1 => n3644, A2 => n3597, ZN => n3598);
   U3594 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => n3872
                           , A3 => n3598, ZN => n3620);
   U3595 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n3599
                           , A3 => n3613, ZN => n3605);
   U3596 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n3873, ZN => n3602);
   U3597 : INV_X1 port map( A => n3600, ZN => n3601);
   U3598 : AOI21_X1 port map( B1 => n3602, B2 => n3601, A => n3622, ZN => n3603
                           );
   U3599 : INV_X1 port map( A => n3603, ZN => n3604);
   U3600 : AOI211_X1 port map( C1 => n3620, C2 => n3612, A => n3605, B => n3604
                           , ZN => n3607);
   U3601 : OAI211_X1 port map( C1 => n3608, C2 => n3637, A => n3607, B => n3606
                           , ZN => cu_i_N265);
   U3602 : MUX2_X1 port map( A => datapath_i_val_b_i_3_port, B => 
                           datapath_i_val_immediate_i_3_port, S => n3831, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U3603 : NOR2_X1 port map( A1 => n3879, A2 => n1152, ZN => n3609);
   U3604 : NOR2_X1 port map( A1 => n704, A2 => cu_i_cw1_4_port, ZN => n3638);
   U3605 : NOR2_X1 port map( A1 => n3609, A2 => n3638, ZN => n3610);
   U3606 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n3610, ZN => n3870);
   U3607 : INV_X1 port map( A => n3610, ZN => n3855);
   U3608 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n3855, ZN => n3868);
   U3609 : CLKBUF_X1 port map( A => n3868, Z => n3857);
   U3610 : CLKBUF_X1 port map( A => n3855, Z => n3867);
   U3611 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n3867, ZN => n3611);
   U3612 : OAI21_X1 port map( B1 => n691, B2 => n3859, A => n3611, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U3613 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_4_port, A3 => n3612, ZN => 
                           n3633);
   U3614 : NOR2_X1 port map( A1 => n3872, A2 => n3613, ZN => n3624);
   U3615 : AOI21_X1 port map( B1 => n3644, B2 => n3633, A => n3624, ZN => n3619
                           );
   U3616 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n3614, B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           n3620, ZN => n3618);
   U3617 : NAND3_X1 port map( A1 => n3616, A2 => n3615, A3 => n3873, ZN => 
                           n3617);
   U3618 : OAI211_X1 port map( C1 => curr_instruction_to_cu_i_0_port, C2 => 
                           n3619, A => n3618, B => n3617, ZN => cu_i_N264);
   U3619 : AND2_X1 port map( A1 => n3887, A2 => curr_instruction_to_cu_i_5_port
                           , ZN => n3628);
   U3620 : INV_X1 port map( A => n3620, ZN => n3627);
   U3621 : NOR3_X1 port map( A1 => n3871, A2 => n3883, A3 => n3637, ZN => n3621
                           );
   U3622 : AOI211_X1 port map( C1 => curr_instruction_to_cu_i_26_port, C2 => 
                           n3623, A => n3622, B => n3621, ZN => n3626);
   U3623 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           n3624, A3 => n3884, ZN => n3625);
   U3624 : OAI211_X1 port map( C1 => n3628, C2 => n3627, A => n3626, B => n3625
                           , ZN => cu_i_N266);
   U3625 : NAND2_X1 port map( A1 => n704, A2 => n3632, ZN => cu_i_N274);
   U3626 : AOI221_X1 port map( B1 => cu_i_n125, B2 => cu_i_n26, C1 => n3874, C2
                           => n3881, A => n3632, ZN => cu_i_N275);
   U3627 : OAI21_X1 port map( B1 => cu_i_n26, B2 => cu_i_n125, A => n3761, ZN 
                           => n3629);
   U3628 : AOI22_X1 port map( A1 => cu_i_n25, A2 => n3630, B1 => n3629, B2 => 
                           n3888, ZN => cu_i_N276);
   U3629 : INV_X1 port map( A => n3631, ZN => n3762);
   U3630 : AOI211_X1 port map( C1 => n704, C2 => cu_i_n145, A => n3762, B => 
                           n3632, ZN => cu_i_N279);
   U3631 : NAND4_X1 port map( A1 => n3634, A2 => n3633, A3 => n3876, A4 => 
                           n3872, ZN => n3635);
   U3632 : OAI21_X1 port map( B1 => n3637, B2 => n3636, A => n3635, ZN => 
                           cu_i_cmd_word_8_port);
   U3633 : MUX2_X1 port map( A => cu_i_cmd_word_8_port, B => cu_i_cw1_12_port, 
                           S => n3654, Z => alu_cin_i);
   U3634 : AOI21_X1 port map( B1 => n756, B2 => n704, A => n3638, ZN => 
                           cu_i_cw1_i_4_port);
   U3635 : MUX2_X1 port map( A => cu_i_cw2_7_port, B => cu_i_cw1_7_port, S => 
                           n3879, Z => cu_i_cw1_i_7_port);
   U3636 : MUX2_X1 port map( A => cu_i_cw2_8_port, B => cu_i_cw1_8_port, S => 
                           n3879, Z => cu_i_cw1_i_8_port);
   U3637 : INV_X1 port map( A => n3639, ZN => n3647);
   U3638 : INV_X1 port map( A => n3644, ZN => n3646);
   U3639 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_14_port, A2 => 
                           curr_instruction_to_cu_i_15_port, A3 => 
                           curr_instruction_to_cu_i_11_port, A4 => 
                           curr_instruction_to_cu_i_12_port, ZN => n3640);
   U3640 : NAND2_X1 port map( A1 => n740, A2 => n3640, ZN => n3645);
   U3641 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_19_port, A2 => 
                           curr_instruction_to_cu_i_20_port, A3 => 
                           curr_instruction_to_cu_i_16_port, A4 => 
                           curr_instruction_to_cu_i_17_port, ZN => n3642);
   U3642 : AOI21_X1 port map( B1 => n697, B2 => n3642, A => n3641, ZN => n3643)
                           ;
   U3643 : AOI221_X1 port map( B1 => n3647, B2 => n3646, C1 => n3645, C2 => 
                           n3644, A => n3643, ZN => n3651);
   U3644 : OAI211_X1 port map( C1 => n3651, C2 => n3650, A => n3649, B => n3648
                           , ZN => cu_i_n209);
   U3645 : NOR2_X1 port map( A1 => cu_i_n123, A2 => cu_i_n23, ZN => cu_i_n210);
   U3646 : AOI22_X1 port map( A1 => n704, A2 => n699, B1 => n3889, B2 => n3879,
                           ZN => cu_i_n131);
   U3647 : MUX2_X1 port map( A => cu_i_cw2_6_port, B => cu_i_cw1_6_port, S => 
                           n3654, Z => cu_i_n127);
   U3648 : MUX2_X1 port map( A => cu_i_cw2_5_port, B => cu_i_cw1_5_port, S => 
                           n3654, Z => cu_i_n126);
   U3649 : MUX2_X1 port map( A => curr_instruction_to_cu_i_31_port, B => 
                           IRAM_DATA(31), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U3650 : MUX2_X1 port map( A => curr_instruction_to_cu_i_30_port, B => 
                           IRAM_DATA(30), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U3651 : MUX2_X1 port map( A => n3882, B => IRAM_DATA(29), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U3652 : MUX2_X1 port map( A => curr_instruction_to_cu_i_28_port, B => 
                           IRAM_DATA(28), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U3653 : MUX2_X1 port map( A => curr_instruction_to_cu_i_27_port, B => 
                           IRAM_DATA(27), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U3654 : MUX2_X1 port map( A => curr_instruction_to_cu_i_26_port, B => 
                           IRAM_DATA(26), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U3655 : MUX2_X1 port map( A => datapath_i_n9, B => IRAM_DATA(25), S => n3654
                           , Z => datapath_i_fetch_stage_dp_n63);
   U3656 : MUX2_X1 port map( A => datapath_i_n10, B => IRAM_DATA(24), S => 
                           n3654, Z => datapath_i_fetch_stage_dp_n62);
   U3657 : MUX2_X1 port map( A => datapath_i_n11, B => IRAM_DATA(23), S => 
                           n3654, Z => datapath_i_fetch_stage_dp_n61);
   U3658 : MUX2_X1 port map( A => datapath_i_n12, B => IRAM_DATA(22), S => 
                           n3879, Z => datapath_i_fetch_stage_dp_n60);
   U3659 : MUX2_X1 port map( A => datapath_i_n13, B => IRAM_DATA(21), S => 
                           n3879, Z => datapath_i_fetch_stage_dp_n59);
   U3660 : MUX2_X1 port map( A => curr_instruction_to_cu_i_20_port, B => 
                           IRAM_DATA(20), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U3661 : MUX2_X1 port map( A => curr_instruction_to_cu_i_19_port, B => 
                           IRAM_DATA(19), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U3662 : NAND2_X1 port map( A1 => n3879, A2 => IRAM_DATA(18), ZN => n3652);
   U3663 : OAI21_X1 port map( B1 => n3879, B2 => n697, A => n3652, ZN => 
                           datapath_i_fetch_stage_dp_n56);
   U3664 : MUX2_X1 port map( A => curr_instruction_to_cu_i_17_port, B => 
                           IRAM_DATA(17), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U3665 : MUX2_X1 port map( A => curr_instruction_to_cu_i_16_port, B => 
                           IRAM_DATA(16), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U3666 : MUX2_X1 port map( A => curr_instruction_to_cu_i_15_port, B => 
                           IRAM_DATA(15), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U3667 : MUX2_X1 port map( A => curr_instruction_to_cu_i_14_port, B => 
                           IRAM_DATA(14), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U3668 : NAND2_X1 port map( A1 => n3879, A2 => IRAM_DATA(13), ZN => n3653);
   U3669 : OAI21_X1 port map( B1 => n3654, B2 => n740, A => n3653, ZN => 
                           datapath_i_fetch_stage_dp_n51);
   U3670 : MUX2_X1 port map( A => curr_instruction_to_cu_i_12_port, B => 
                           IRAM_DATA(12), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U3671 : MUX2_X1 port map( A => curr_instruction_to_cu_i_11_port, B => 
                           IRAM_DATA(11), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U3672 : MUX2_X1 port map( A => datapath_i_n14, B => IRAM_DATA(10), S => 
                           n3654, Z => datapath_i_fetch_stage_dp_n48);
   U3673 : MUX2_X1 port map( A => datapath_i_n15, B => IRAM_DATA(9), S => n3654
                           , Z => datapath_i_fetch_stage_dp_n47);
   U3674 : MUX2_X1 port map( A => datapath_i_n16, B => IRAM_DATA(8), S => n3879
                           , Z => datapath_i_fetch_stage_dp_n46);
   U3675 : MUX2_X1 port map( A => datapath_i_n17, B => IRAM_DATA(7), S => n3654
                           , Z => datapath_i_fetch_stage_dp_n45);
   U3676 : MUX2_X1 port map( A => datapath_i_n18, B => IRAM_DATA(6), S => n3654
                           , Z => datapath_i_fetch_stage_dp_n44);
   U3677 : MUX2_X1 port map( A => curr_instruction_to_cu_i_5_port, B => 
                           IRAM_DATA(5), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U3678 : MUX2_X1 port map( A => curr_instruction_to_cu_i_4_port, B => 
                           IRAM_DATA(4), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U3679 : MUX2_X1 port map( A => curr_instruction_to_cu_i_3_port, B => 
                           IRAM_DATA(3), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U3680 : MUX2_X1 port map( A => curr_instruction_to_cu_i_2_port, B => 
                           IRAM_DATA(2), S => n3879, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U3681 : MUX2_X1 port map( A => curr_instruction_to_cu_i_1_port, B => 
                           IRAM_DATA(1), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U3682 : MUX2_X1 port map( A => curr_instruction_to_cu_i_0_port, B => 
                           IRAM_DATA(0), S => n3654, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U3683 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_0_port, 
                           B2 => n3747, ZN => n3655);
   U3684 : OAI21_X1 port map( B1 => n733, B2 => n3750, A => n3655, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U3685 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N39_port, B => 
                           datapath_i_fetch_stage_dp_N5, S => n3660, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U3686 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_1_port, 
                           B2 => n3747, ZN => n3656);
   U3687 : OAI21_X1 port map( B1 => n734, B2 => n3750, A => n3656, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U3688 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N40_port, B => 
                           datapath_i_fetch_stage_dp_N6, S => n3660, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U3689 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n3657, ZN => n3658);
   U3690 : AOI22_X1 port map( A1 => n3756, A2 => n3658, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n3753, ZN => datapath_i_fetch_stage_dp_n35);
   U3691 : OAI21_X1 port map( B1 => n3659, B2 => IRAM_ADDRESS_3_port, A => 
                           n3708, ZN => n3662);
   U3692 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n3664);
   U3693 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           B2 => datapath_i_new_pc_value_mem_stage_i_3_port, A 
                           => n3660, ZN => n3661);
   U3694 : OAI22_X1 port map( A1 => n3666, A2 => n3662, B1 => n3664, B2 => 
                           n3661, ZN => datapath_i_fetch_stage_dp_n34);
   U3695 : OAI211_X1 port map( C1 => n3664, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n3753, B => n3663, ZN => n3668);
   U3696 : OAI211_X1 port map( C1 => n3666, C2 => IRAM_ADDRESS_4_port, A => 
                           n3756, B => n3665, ZN => n3667);
   U3697 : NAND2_X1 port map( A1 => n3668, A2 => n3667, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U3698 : OAI211_X1 port map( C1 => n3670, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n3753, B => n3669, ZN => n3674);
   U3699 : OAI211_X1 port map( C1 => n3672, C2 => IRAM_ADDRESS_6_port, A => 
                           n3756, B => n3671, ZN => n3673);
   U3700 : NAND2_X1 port map( A1 => n3674, A2 => n3673, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U3701 : OAI211_X1 port map( C1 => n3676, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n3753, B => n3675, ZN => n3680);
   U3702 : OAI211_X1 port map( C1 => n3678, C2 => IRAM_ADDRESS_8_port, A => 
                           n3756, B => n3677, ZN => n3679);
   U3703 : NAND2_X1 port map( A1 => n3680, A2 => n3679, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U3704 : OAI211_X1 port map( C1 => n3682, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n3753, B => n3681, ZN => n3686);
   U3705 : OAI211_X1 port map( C1 => n3684, C2 => IRAM_ADDRESS_10_port, A => 
                           n3756, B => n3683, ZN => n3685);
   U3706 : NAND2_X1 port map( A1 => n3686, A2 => n3685, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U3707 : OAI211_X1 port map( C1 => n3688, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n3753, B => n3687, ZN => n3692);
   U3708 : OAI211_X1 port map( C1 => n3690, C2 => IRAM_ADDRESS_12_port, A => 
                           n3708, B => n3689, ZN => n3691);
   U3709 : NAND2_X1 port map( A1 => n3692, A2 => n3691, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U3710 : OAI211_X1 port map( C1 => n3694, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n3753, B => n3693, ZN => n3698);
   U3711 : OAI211_X1 port map( C1 => n3696, C2 => IRAM_ADDRESS_14_port, A => 
                           n3708, B => n3695, ZN => n3697);
   U3712 : NAND2_X1 port map( A1 => n3698, A2 => n3697, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U3713 : OAI211_X1 port map( C1 => n3700, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n3753, B => n3699, ZN => n3704);
   U3714 : OAI211_X1 port map( C1 => n3702, C2 => IRAM_ADDRESS_16_port, A => 
                           n3708, B => n3701, ZN => n3703);
   U3715 : NAND2_X1 port map( A1 => n3704, A2 => n3703, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U3716 : OAI211_X1 port map( C1 => n3706, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n3753, B => n3705, ZN => n3711);
   U3717 : OAI211_X1 port map( C1 => n3709, C2 => IRAM_ADDRESS_18_port, A => 
                           n3708, B => n3707, ZN => n3710);
   U3718 : NAND2_X1 port map( A1 => n3711, A2 => n3710, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U3719 : OAI211_X1 port map( C1 => n3713, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n3753, B => n3712, ZN => n3717);
   U3720 : OAI211_X1 port map( C1 => n3715, C2 => IRAM_ADDRESS_20_port, A => 
                           n3756, B => n3714, ZN => n3716);
   U3721 : NAND2_X1 port map( A1 => n3717, A2 => n3716, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U3722 : OAI211_X1 port map( C1 => n3719, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n3753, B => n3718, ZN => n3723);
   U3723 : OAI211_X1 port map( C1 => n3721, C2 => IRAM_ADDRESS_22_port, A => 
                           n3756, B => n3720, ZN => n3722);
   U3724 : NAND2_X1 port map( A1 => n3723, A2 => n3722, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U3725 : OAI211_X1 port map( C1 => n3725, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n3753, B => n3724, ZN => n3729);
   U3726 : OAI211_X1 port map( C1 => n3727, C2 => IRAM_ADDRESS_24_port, A => 
                           n3756, B => n3726, ZN => n3728);
   U3727 : NAND2_X1 port map( A1 => n3729, A2 => n3728, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U3728 : OAI211_X1 port map( C1 => n3731, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n3753, B => n3730, ZN => n3735);
   U3729 : OAI211_X1 port map( C1 => n3733, C2 => IRAM_ADDRESS_26_port, A => 
                           n3756, B => n3732, ZN => n3734);
   U3730 : NAND2_X1 port map( A1 => n3735, A2 => n3734, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U3731 : OAI211_X1 port map( C1 => n3737, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n3753, B => n3736, ZN => n3741);
   U3732 : OAI211_X1 port map( C1 => n3739, C2 => IRAM_ADDRESS_28_port, A => 
                           n3756, B => n3738, ZN => n3740);
   U3733 : NAND2_X1 port map( A1 => n3741, A2 => n3740, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U3734 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n3748, B1 => datapath_i_alu_output_val_i_30_port,
                           B2 => n3747, ZN => n3742);
   U3735 : OAI21_X1 port map( B1 => n727, B2 => n3750, A => n3742, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   U3736 : NAND2_X1 port map( A1 => n3743, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n3752);
   U3737 : OAI211_X1 port map( C1 => n3743, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n3753, B => n3752, ZN => n3746);
   U3738 : NAND2_X1 port map( A1 => n3744, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n3751);
   U3739 : OAI211_X1 port map( C1 => n3744, C2 => IRAM_ADDRESS_30_port, A => 
                           n3756, B => n3751, ZN => n3745);
   U3740 : NAND2_X1 port map( A1 => n3746, A2 => n3745, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U3741 : AOI22_X1 port map( A1 => n3748, A2 => 
                           datapath_i_new_pc_value_decode_31_port, B1 => 
                           datapath_i_alu_output_val_i_31_port, B2 => n3747, ZN
                           => n3749);
   U3742 : OAI21_X1 port map( B1 => n703, B2 => n3750, A => n3749, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U3743 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n3751, Z => n3755)
                           ;
   U3744 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n3752, Z => n3754);
   U3745 : AOI22_X1 port map( A1 => n3756, A2 => n3755, B1 => n3754, B2 => 
                           n3753, ZN => datapath_i_fetch_stage_dp_n2);
   U3746 : OAI21_X1 port map( B1 => n737, B2 => n3757, A => n3758, ZN => 
                           read_rf_p2_i);
   U3747 : OAI221_X1 port map( B1 => n3759, B2 => n697, C1 => n3758, C2 => n740
                           , A => n3802, ZN => datapath_i_decode_stage_dp_n78);
   U3748 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ZN => n3760);
   U3749 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n3760, ZN => n3776);
   U3750 : INV_X1 port map( A => n3776, ZN => n3785);
   U3751 : AND2_X2 port map( A1 => n3785, A2 => n3763, ZN => n3799);
   U3752 : NOR2_X1 port map( A1 => n3776, A2 => n3763, ZN => n3798);
   U3753 : CLKBUF_X1 port map( A => n3798, Z => n3789);
   U3754 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_0_port, ZN => n3764
                           );
   U3755 : OAI21_X1 port map( B1 => n733, B2 => n3785, A => n3764, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U3756 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_1_port, ZN => n3765
                           );
   U3757 : OAI21_X1 port map( B1 => n734, B2 => n3785, A => n3765, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U3758 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_2_port, ZN => n3766
                           );
   U3759 : OAI21_X1 port map( B1 => n728, B2 => n3785, A => n3766, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U3760 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_3_port, ZN => n3767
                           );
   U3761 : OAI21_X1 port map( B1 => n729, B2 => n3785, A => n3767, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U3762 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_4_port, ZN => n3768
                           );
   U3763 : OAI21_X1 port map( B1 => n730, B2 => n3785, A => n3768, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U3764 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_5_port, ZN => n3769
                           );
   U3765 : OAI21_X1 port map( B1 => n731, B2 => n3785, A => n3769, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U3766 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_6_port, ZN => n3770
                           );
   U3767 : OAI21_X1 port map( B1 => n732, B2 => n3785, A => n3770, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U3768 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_7_port, ZN => n3771
                           );
   U3769 : OAI21_X1 port map( B1 => n705, B2 => n3785, A => n3771, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U3770 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_8_port, ZN => n3772
                           );
   U3771 : OAI21_X1 port map( B1 => n706, B2 => n3785, A => n3772, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U3772 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_9_port, ZN => n3773
                           );
   U3773 : OAI21_X1 port map( B1 => n707, B2 => n3785, A => n3773, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U3774 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => 
                           n3774);
   U3775 : OAI21_X1 port map( B1 => n708, B2 => n3785, A => n3774, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U3776 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => 
                           n3775);
   U3777 : OAI21_X1 port map( B1 => n709, B2 => n3785, A => n3775, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U3778 : INV_X1 port map( A => n3776, ZN => n3801);
   U3779 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => 
                           n3777);
   U3780 : OAI21_X1 port map( B1 => n710, B2 => n3801, A => n3777, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U3781 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => 
                           n3778);
   U3782 : OAI21_X1 port map( B1 => n711, B2 => n3785, A => n3778, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U3783 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => 
                           n3779);
   U3784 : OAI21_X1 port map( B1 => n712, B2 => n3801, A => n3779, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U3785 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => 
                           n3780);
   U3786 : OAI21_X1 port map( B1 => n713, B2 => n3785, A => n3780, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U3787 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => 
                           n3781);
   U3788 : OAI21_X1 port map( B1 => n714, B2 => n3801, A => n3781, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U3789 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => 
                           n3782);
   U3790 : OAI21_X1 port map( B1 => n715, B2 => n3785, A => n3782, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U3791 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => 
                           n3783);
   U3792 : OAI21_X1 port map( B1 => n716, B2 => n3801, A => n3783, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U3793 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => 
                           n3784);
   U3794 : OAI21_X1 port map( B1 => n717, B2 => n3785, A => n3784, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U3795 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => 
                           n3786);
   U3796 : OAI21_X1 port map( B1 => n718, B2 => n3801, A => n3786, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U3797 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => 
                           n3787);
   U3798 : OAI21_X1 port map( B1 => n719, B2 => n3801, A => n3787, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U3799 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => 
                           n3788);
   U3800 : OAI21_X1 port map( B1 => n720, B2 => n3801, A => n3788, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U3801 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n3789, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => 
                           n3790);
   U3802 : OAI21_X1 port map( B1 => n721, B2 => n3801, A => n3790, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U3803 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => 
                           n3791);
   U3804 : OAI21_X1 port map( B1 => n722, B2 => n3801, A => n3791, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U3805 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => 
                           n3792);
   U3806 : OAI21_X1 port map( B1 => n723, B2 => n3801, A => n3792, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U3807 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => 
                           n3793);
   U3808 : OAI21_X1 port map( B1 => n691, B2 => n3801, A => n3793, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U3809 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => 
                           n3794);
   U3810 : OAI21_X1 port map( B1 => n724, B2 => n3801, A => n3794, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U3811 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => 
                           n3795);
   U3812 : OAI21_X1 port map( B1 => n725, B2 => n3801, A => n3795, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U3813 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => 
                           n3796);
   U3814 : OAI21_X1 port map( B1 => n726, B2 => n3801, A => n3796, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U3815 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => 
                           n3797);
   U3816 : OAI21_X1 port map( B1 => n727, B2 => n3801, A => n3797, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U3817 : AOI22_X1 port map( A1 => n3799, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n3798, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => 
                           n3800);
   U3818 : OAI21_X1 port map( B1 => n703, B2 => n3801, A => n3800, ZN => 
                           datapath_i_decode_stage_dp_n12);
   U3819 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n3803, A => n3802, ZN => cu_i_cmd_word_6_port);
   U3820 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_6_port, B1 => 
                           cu_i_cw1_10_port, B2 => n3879, ZN => n3817);
   U3821 : NOR4_X1 port map( A1 => datapath_i_val_a_i_14_port, A2 => 
                           datapath_i_val_a_i_15_port, A3 => 
                           datapath_i_val_a_i_16_port, A4 => 
                           datapath_i_val_a_i_17_port, ZN => n3807);
   U3822 : NOR4_X1 port map( A1 => datapath_i_val_a_i_18_port, A2 => 
                           datapath_i_val_a_i_19_port, A3 => 
                           datapath_i_val_a_i_20_port, A4 => 
                           datapath_i_val_a_i_21_port, ZN => n3806);
   U3823 : NOR4_X1 port map( A1 => datapath_i_val_a_i_26_port, A2 => 
                           datapath_i_val_a_i_7_port, A3 => 
                           datapath_i_val_a_i_8_port, A4 => 
                           datapath_i_val_a_i_9_port, ZN => n3805);
   U3824 : NOR4_X1 port map( A1 => datapath_i_val_a_i_10_port, A2 => 
                           datapath_i_val_a_i_11_port, A3 => 
                           datapath_i_val_a_i_12_port, A4 => 
                           datapath_i_val_a_i_13_port, ZN => n3804);
   U3825 : NAND4_X1 port map( A1 => n3807, A2 => n3806, A3 => n3805, A4 => 
                           n3804, ZN => n3813);
   U3826 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n3811);
   U3827 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n3810);
   U3828 : NOR4_X1 port map( A1 => datapath_i_val_a_i_22_port, A2 => 
                           datapath_i_val_a_i_23_port, A3 => 
                           datapath_i_val_a_i_24_port, A4 => 
                           datapath_i_val_a_i_25_port, ZN => n3809);
   U3829 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n3808);
   U3830 : NAND4_X1 port map( A1 => n3811, A2 => n3810, A3 => n3809, A4 => 
                           n3808, ZN => n3812);
   U3831 : NOR2_X1 port map( A1 => n3813, A2 => n3812, ZN => n3815);
   U3832 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_7_port, B1 => 
                           cu_i_cw1_11_port, B2 => n3879, ZN => n3814);
   U3833 : NAND2_X1 port map( A1 => n3815, A2 => n3814, ZN => n3816);
   U3834 : OAI22_X1 port map( A1 => n3817, A2 => n3816, B1 => n3815, B2 => 
                           n3814, ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U3835 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, S 
                           => n3892, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U3836 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U3837 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, S 
                           => n3892, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U3838 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U3839 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, S 
                           => n3892, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U3840 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U3841 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U3842 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U3843 : NAND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
                           A2 => n3892, ZN => n3830);
   U3844 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
                           ZN => n3818);
   U3845 : NAND2_X1 port map( A1 => n3830, A2 => n3818, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U3846 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
                           ZN => n3819);
   U3847 : NAND2_X1 port map( A1 => n3830, A2 => n3819, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U3848 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
                           ZN => n3820);
   U3849 : NAND2_X1 port map( A1 => n3830, A2 => n3820, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U3850 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
                           ZN => n3821);
   U3851 : NAND2_X1 port map( A1 => n3830, A2 => n3821, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U3852 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
                           ZN => n3822);
   U3853 : NAND2_X1 port map( A1 => n3830, A2 => n3822, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U3854 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
                           ZN => n3823);
   U3855 : NAND2_X1 port map( A1 => n3830, A2 => n3823, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U3856 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
                           ZN => n3824);
   U3857 : NAND2_X1 port map( A1 => n3830, A2 => n3824, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U3858 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
                           ZN => n3825);
   U3859 : NAND2_X1 port map( A1 => n3830, A2 => n3825, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U3860 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
                           ZN => n3826);
   U3861 : NAND2_X1 port map( A1 => n3830, A2 => n3826, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U3862 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
                           ZN => n3827);
   U3863 : NAND2_X1 port map( A1 => n3830, A2 => n3827, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U3864 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U3865 : NAND2_X1 port map( A1 => n3828, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
                           ZN => n3829);
   U3866 : NAND2_X1 port map( A1 => n3830, A2 => n3829, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U3867 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U3868 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U3869 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U3870 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U3871 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U3872 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, S 
                           => n3891, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U3873 : MUX2_X1 port map( A => datapath_i_val_b_i_7_port, B => 
                           datapath_i_val_immediate_i_7_port, S => n3831, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U3874 : MUX2_X1 port map( A => datapath_i_val_b_i_8_port, B => 
                           datapath_i_val_immediate_i_8_port, S => n3831, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U3875 : MUX2_X1 port map( A => datapath_i_val_b_i_9_port, B => 
                           datapath_i_val_immediate_i_9_port, S => n3831, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U3876 : MUX2_X1 port map( A => datapath_i_val_b_i_10_port, B => 
                           datapath_i_val_immediate_i_10_port, S => n3831, Z =>
                           datapath_i_execute_stage_dp_opb_10_port);
   U3877 : MUX2_X1 port map( A => datapath_i_val_b_i_11_port, B => 
                           datapath_i_val_immediate_i_11_port, S => n3831, Z =>
                           datapath_i_execute_stage_dp_opb_11_port);
   U3878 : MUX2_X1 port map( A => datapath_i_val_b_i_12_port, B => 
                           datapath_i_val_immediate_i_12_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_12_port);
   U3879 : MUX2_X1 port map( A => datapath_i_val_b_i_13_port, B => 
                           datapath_i_val_immediate_i_13_port, S => n3831, Z =>
                           datapath_i_execute_stage_dp_opb_13_port);
   U3880 : MUX2_X1 port map( A => datapath_i_val_b_i_14_port, B => 
                           datapath_i_val_immediate_i_14_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_14_port);
   U3881 : MUX2_X1 port map( A => datapath_i_val_b_i_15_port, B => 
                           datapath_i_val_immediate_i_15_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_15_port);
   U3882 : MUX2_X1 port map( A => datapath_i_val_b_i_16_port, B => 
                           datapath_i_val_immediate_i_16_port, S => n3831, Z =>
                           datapath_i_execute_stage_dp_opb_16_port);
   U3883 : MUX2_X1 port map( A => datapath_i_val_b_i_17_port, B => 
                           datapath_i_val_immediate_i_17_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_17_port);
   U3884 : MUX2_X1 port map( A => datapath_i_val_b_i_18_port, B => 
                           datapath_i_val_immediate_i_18_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_18_port);
   U3885 : MUX2_X1 port map( A => datapath_i_val_b_i_19_port, B => 
                           datapath_i_val_immediate_i_19_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_19_port);
   U3886 : MUX2_X1 port map( A => datapath_i_val_b_i_20_port, B => 
                           datapath_i_val_immediate_i_20_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_20_port);
   U3887 : MUX2_X1 port map( A => datapath_i_val_b_i_21_port, B => 
                           datapath_i_val_immediate_i_21_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_21_port);
   U3888 : MUX2_X1 port map( A => datapath_i_val_b_i_22_port, B => 
                           datapath_i_val_immediate_i_22_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_22_port);
   U3889 : MUX2_X1 port map( A => datapath_i_val_b_i_23_port, B => 
                           datapath_i_val_immediate_i_23_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_23_port);
   U3890 : MUX2_X1 port map( A => datapath_i_val_b_i_24_port, B => 
                           datapath_i_val_immediate_i_24_port, S => n3833, Z =>
                           datapath_i_execute_stage_dp_opb_24_port);
   U3891 : NAND2_X1 port map( A1 => n3833, A2 => 
                           datapath_i_val_immediate_i_25_port, ZN => n3832);
   U3892 : OAI21_X1 port map( B1 => n3833, B2 => n758, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U3893 : OAI21_X1 port map( B1 => n3833, B2 => n759, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U3894 : OAI21_X1 port map( B1 => n3833, B2 => n760, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U3895 : OAI21_X1 port map( B1 => n3833, B2 => n761, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U3896 : OAI21_X1 port map( B1 => n3833, B2 => n762, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U3897 : OAI21_X1 port map( B1 => n3833, B2 => n763, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U3898 : OAI21_X1 port map( B1 => n3833, B2 => n764, A => n3832, ZN => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U3899 : MUX2_X1 port map( A => datapath_i_val_b_i_4_port, B => 
                           datapath_i_val_immediate_i_4_port, S => n3833, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U3900 : MUX2_X1 port map( A => datapath_i_val_b_i_5_port, B => 
                           datapath_i_val_immediate_i_5_port, S => n3833, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U3901 : MUX2_X1 port map( A => datapath_i_val_b_i_6_port, B => 
                           datapath_i_val_immediate_i_6_port, S => n3833, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U3902 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_7_port, B2 => 
                           n3855, ZN => n3834);
   U3903 : OAI21_X1 port map( B1 => n705, B2 => n3870, A => n3834, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U3904 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_8_port, B2 => 
                           n3867, ZN => n3835);
   U3905 : OAI21_X1 port map( B1 => n706, B2 => n3859, A => n3835, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U3906 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_9_port, B2 => 
                           n3855, ZN => n3836);
   U3907 : OAI21_X1 port map( B1 => n707, B2 => n3870, A => n3836, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U3908 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n3867, ZN => n3837);
   U3909 : OAI21_X1 port map( B1 => n708, B2 => n3859, A => n3837, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U3910 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n3855, ZN => n3838);
   U3911 : OAI21_X1 port map( B1 => n709, B2 => n3870, A => n3838, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U3912 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n3867, ZN => n3839);
   U3913 : OAI21_X1 port map( B1 => n710, B2 => n3859, A => n3839, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U3914 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n3855, ZN => n3840);
   U3915 : OAI21_X1 port map( B1 => n711, B2 => n3870, A => n3840, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U3916 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n3867, ZN => n3841);
   U3917 : OAI21_X1 port map( B1 => n712, B2 => n3859, A => n3841, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U3918 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n3855, ZN => n3842);
   U3919 : OAI21_X1 port map( B1 => n713, B2 => n3870, A => n3842, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U3920 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n3855, ZN => n3843);
   U3921 : OAI21_X1 port map( B1 => n714, B2 => n3870, A => n3843, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U3922 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n3867, ZN => n3844);
   U3923 : OAI21_X1 port map( B1 => n715, B2 => n3870, A => n3844, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U3924 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n3855, ZN => n3845);
   U3925 : OAI21_X1 port map( B1 => n716, B2 => n3859, A => n3845, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U3926 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n3867, ZN => n3846);
   U3927 : OAI21_X1 port map( B1 => n717, B2 => n3859, A => n3846, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U3928 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n3855, ZN => n3847);
   U3929 : OAI21_X1 port map( B1 => n718, B2 => n3859, A => n3847, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U3930 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n3867, ZN => n3848);
   U3931 : OAI21_X1 port map( B1 => n719, B2 => n3859, A => n3848, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U3932 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n3855, ZN => n3849);
   U3933 : OAI21_X1 port map( B1 => n720, B2 => n3859, A => n3849, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U3934 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n3855, ZN => n3850);
   U3935 : OAI21_X1 port map( B1 => n721, B2 => n3859, A => n3850, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U3936 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n3855, ZN => n3851);
   U3937 : OAI21_X1 port map( B1 => n722, B2 => n3859, A => n3851, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U3938 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n3855, ZN => n3852);
   U3939 : OAI21_X1 port map( B1 => n723, B2 => n3859, A => n3852, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U3940 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_0_port, B2 => 
                           n3855, ZN => n3853);
   U3941 : OAI21_X1 port map( B1 => n733, B2 => n3859, A => n3853, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U3942 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n3855, ZN => n3854);
   U3943 : OAI21_X1 port map( B1 => n724, B2 => n3859, A => n3854, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U3944 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n3855, ZN => n3856);
   U3945 : OAI21_X1 port map( B1 => n725, B2 => n3859, A => n3856, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U3946 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n3857, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n3867, ZN => n3858);
   U3947 : OAI21_X1 port map( B1 => n726, B2 => n3859, A => n3858, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U3948 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n3867, ZN => n3860);
   U3949 : OAI21_X1 port map( B1 => n727, B2 => n3870, A => n3860, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U3950 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n3867, ZN => n3861);
   U3951 : OAI21_X1 port map( B1 => n703, B2 => n3870, A => n3861, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U3952 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_1_port, B2 => 
                           n3867, ZN => n3862);
   U3953 : OAI21_X1 port map( B1 => n734, B2 => n3870, A => n3862, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U3954 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_2_port, B2 => 
                           n3867, ZN => n3863);
   U3955 : OAI21_X1 port map( B1 => n728, B2 => n3870, A => n3863, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U3956 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_3_port, B2 => 
                           n3867, ZN => n3864);
   U3957 : OAI21_X1 port map( B1 => n729, B2 => n3870, A => n3864, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U3958 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_4_port, B2 => 
                           n3867, ZN => n3865);
   U3959 : OAI21_X1 port map( B1 => n730, B2 => n3870, A => n3865, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U3960 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_5_port, B2 => 
                           n3867, ZN => n3866);
   U3961 : OAI21_X1 port map( B1 => n731, B2 => n3870, A => n3866, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U3962 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n3868, B1 => datapath_i_val_a_i_6_port, B2 => 
                           n3867, ZN => n3869);
   U3963 : OAI21_X1 port map( B1 => n732, B2 => n3870, A => n3869, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);

end SYN_dlx_rtl;
