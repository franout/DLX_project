
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal DATA2_I_30_port, DATA2_I_28_port, DATA2_I_27_port, DATA2_I_26_port, 
      DATA2_I_25_port, DATA2_I_24_port, DATA2_I_23_port, DATA2_I_22_port, 
      DATA2_I_21_port, DATA2_I_20_port, DATA2_I_19_port, DATA2_I_18_port, 
      DATA2_I_17_port, DATA2_I_16_port, DATA2_I_15_port, DATA2_I_14_port, 
      DATA2_I_13_port, DATA2_I_12_port, DATA2_I_11_port, DATA2_I_10_port, 
      DATA2_I_9_port, DATA2_I_8_port, DATA2_I_7_port, DATA2_I_6_port, 
      DATA2_I_5_port, DATA2_I_4_port, DATA2_I_3_port, DATA2_I_2_port, 
      DATA2_I_1_port, DATA2_I_0_port, data1_mul_15_port, data1_mul_0_port, 
      data2_mul_2_port, data2_mul_1_port, N2517, N2518, N2519, N2520, N2521, 
      N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n554, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1429, 
      n2808, n3020, n3026, n3027, n3028, n3029, n3030, n3036, n3940, n3957, 
      n3958, n3973, n3974, n3990, n3991, n3992, n3993, n3994, n3995, n3996, 
      n4007, n4008, n4009, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4293, n4295, n4302, n4395, n6095, n7769, n7822, n8528, n8534, n8535, 
      n8547, n8548, n8549, n8550, n8551, n8553, n8555, n8565, n8566, n8567, 
      n8571, n8572, n8573, n8574, n8578, n8579, n8581, n8584, n8587, n8588, 
      n8591, n8595, n8596, n8599, n8600, n8601, n8604, n8612, n8626, n8631, 
      n8632, n8634, n8635, n8636, n8638, n8639, n8640, n8642, n8646, n8647, 
      n8649, n8673, n8674, n8675, n8679, n8681, n8682, n8683, n8685, n8686, 
      n8689, n8690, n8692, n8694, n8696, n8698, n8700, n8702, n8704, n8706, 
      n8708, n8710, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, 
      n8721, n8722, n8723, n8724, n8725, n8727, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8744, 
      n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8757, n8762, 
      n8763, n8764, n8765, n8770, n8771, n8772, n8773, n8779, n8780, n8781, 
      n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, 
      n8792, n8793, n8800, n8810, n8811, n8812, n8813, n8814, n8818, n8819, 
      n8820, n8821, n8823, n8824, n8826, n8828, n8830, n8831, n8832, n8834, 
      n8837, n8838, n8847, n8859, n8861, n8867, n8871, n8875, n8880, n8887, 
      n8892, n8900, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, 
      n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, 
      n8929, n8931, n8932, n8933, n8940, n8942, n8943, n8944, n8945, n8946, 
      n8956, n8957, n8978, n8980, n8984, n8990, n9011, n9020, n9045, n9048, 
      n9051, n9054, n9057, n9060, n9063, n9066, n9069, n9072, n9075, n9078, 
      n9081, n9084, n11435, n11436, n11437, n11444, n11447, n11449, n11453, 
      n11457, n11458, n11459, n11469, n11473, n11485, n11526, n11540, n11714, 
      n11729, n11754, n11755, n11789, n11811, n11849, n11927, n11946, n11952, 
      n11955, n11959, n11960, n11966, n11979, n11981, n11996, n12004, n12031, 
      n12032, n12042, n12045, n12047, n12086, n12087, n12088, n12151, n12158, 
      n12162, n12189, n12212, n12213, n12229, n12230, n12246, n12254, n12255, 
      n12263, n12273, n12292, n12306, n12313, n12325, n12392, n12400, n12423, 
      n12446, n12473, n12474, n12487, n12509, n12526, n12527, n12721, n12722, 
      n12750, n12751, n12754, n12924, n12927, n13096, n13099, n13151, n13174, 
      n13175, n13182, n13186, n13848, n13849, n13850, n13851, n13852, n13853, 
      n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, 
      n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, 
      n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, 
      n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13890, 
      n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, 
      n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, 
      n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, 
      n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, 
      n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, 
      n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, 
      n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, 
      n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, 
      n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, 
      n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, 
      n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, 
      n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, 
      n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, 
      n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, 
      n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, 
      n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, 
      n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, 
      n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, 
      n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, 
      n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14070, n14071, 
      n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14080, n14081, 
      n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, 
      n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, 
      n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, 
      n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, 
      n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, 
      n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, 
      n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, 
      n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, 
      n14154, n14155, n14157, n14158, n14159, n14160, n14161, n14162, n14163, 
      n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, 
      n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, 
      n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, 
      n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, 
      n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, 
      n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, 
      n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, 
      n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, 
      n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, 
      n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, 
      n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, 
      n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, 
      n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, 
      n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, 
      n14290, n14291, n14292, n14293, n14294, n14296, n14297, n14298, n14299, 
      n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, 
      n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, 
      n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, 
      n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, 
      n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, 
      n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, 
      n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, 
      n14364, n14365, n14366, n14367, n14368, n14372, n14373, n14374, n14375, 
      n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, 
      n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, 
      n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, 
      n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, 
      n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, 
      n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, 
      n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, 
      n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, 
      n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, 
      n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, 
      n14466, n14467, n14469, n16389, n16390, n16391, n16393, n16394, n16396, 
      n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, 
      n16406, n16407, n16408, n16409, n16410, n16412, n16413, n16414, n16415, 
      n16416, n16417, n16418, n16419, n1808, n1809, n1810, n1811, n1812, n1813,
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
      n1864, n1865, n1866, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, 
      n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, 
      n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, 
      n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, 
      n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, 
      n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, 
      n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, 
      n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, 
      n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, 
      n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, 
      n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, 
      n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, 
      n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, 
      n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, 
      n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, 
      n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, 
      n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, 
      n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, 
      n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, 
      n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, 
      n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, 
      n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, 
      n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, 
      n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, 
      n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, 
      n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, 
      n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, 
      n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, 
      n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, 
      n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, 
      n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, 
      n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, 
      n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, 
      n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, 
      n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, 
      n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, 
      n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, 
      n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, 
      n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, 
      n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, 
      n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, 
      n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, 
      n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, 
      n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, 
      n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, 
      n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, 
      n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, 
      n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, 
      n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, 
      n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, 
      n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, 
      n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, 
      n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, 
      n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, 
      n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, 
      n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, 
      n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, 
      n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, 
      n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, 
      n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, 
      n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, 
      n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, 
      n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, 
      n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, 
      n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, 
      n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, 
      n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, 
      n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, 
      n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, 
      n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, 
      n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, 
      n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, 
      n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, 
      n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, 
      n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, 
      n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, 
      n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, 
      n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, 
      n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, 
      n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, 
      n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, 
      n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, 
      n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, 
      n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, 
      n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, 
      n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, 
      n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, 
      n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, 
      n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, 
      n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, 
      n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, 
      n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, 
      n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, 
      n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, 
      n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, 
      n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, 
      n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, 
      n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, 
      n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, 
      n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, 
      n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, 
      n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, 
      n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, 
      n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, 
      n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, 
      n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, 
      n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, 
      n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, 
      n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, 
      n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, 
      n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, 
      n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, 
      n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, 
      n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, 
      n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, 
      n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, 
      n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, 
      n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, 
      n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, 
      n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, 
      n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, 
      n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, 
      n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, 
      n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, 
      n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, 
      n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, 
      n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, 
      n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, 
      n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, 
      n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, 
      n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, 
      n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, 
      n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, 
      n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, 
      n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, 
      n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, 
      n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, 
      n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, 
      n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, 
      n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, 
      n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, 
      n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, 
      n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, 
      n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, 
      n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, 
      n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, 
      n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, 
      n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, 
      n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, 
      n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, 
      n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, 
      n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, 
      n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, 
      n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, 
      n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, 
      n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, 
      n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, 
      n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, 
      n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, 
      n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, 
      n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, 
      n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, 
      n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, 
      n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, 
      n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, 
      n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, 
      n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, 
      n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, 
      n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, 
      n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, 
      n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, 
      n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, 
      n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, 
      n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, 
      n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, 
      n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, 
      n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, 
      n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, 
      n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, 
      n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, 
      n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, 
      n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, 
      n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, 
      n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, 
      n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, 
      n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, 
      n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, 
      n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, 
      n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, 
      n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, 
      n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, 
      n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, 
      n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, 
      n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, 
      n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, 
      n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, 
      n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, 
      n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, 
      n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, 
      n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, 
      n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, 
      n18229, n18230, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575 : std_logic;

begin
   
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n18230, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n554, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n554, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n554, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n18230, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n554, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n554, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n18230, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n554, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n554, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n554, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n554, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n554, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n554, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n18230, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n554, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n554, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n554, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n554, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n554, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n554, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n554, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n554, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n554, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n18230, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n18230, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n18230, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n18230, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n7822, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n7822, Q => 
                           n9045);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n7822, Q => 
                           n9048);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n7822, Q => 
                           n9051);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n7822, Q => 
                           n9054);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n7822, Q => 
                           n9057);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n7822, Q => 
                           n9060);
   data1_mul_reg_8_inst : DLL_X1 port map( D => n14469, GN => n7822, Q => n9063
                           );
   data1_mul_reg_7_inst : DLL_X1 port map( D => n14467, GN => n7822, Q => n9066
                           );
   data1_mul_reg_6_inst : DLL_X1 port map( D => n14466, GN => n7822, Q => n9069
                           );
   data1_mul_reg_5_inst : DLL_X1 port map( D => n14465, GN => n7822, Q => n9072
                           );
   data1_mul_reg_4_inst : DLL_X1 port map( D => n14464, GN => n7822, Q => n9075
                           );
   data1_mul_reg_3_inst : DLL_X1 port map( D => n14326, GN => n7822, Q => n9078
                           );
   data1_mul_reg_2_inst : DLL_X1 port map( D => n14327, GN => n7822, Q => n9081
                           );
   data1_mul_reg_1_inst : DLL_X1 port map( D => n14463, GN => n7822, Q => n9084
                           );
   data1_mul_reg_0_inst : DLL_X1 port map( D => n14461, GN => n7822, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n7822, Q => 
                           n13182);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n7822, Q => 
                           n8990);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n7822, Q => 
                           n13175);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n7822, Q => 
                           n8984);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n7822, Q => 
                           n13174);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n7822, Q => 
                           n8980);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n7822, Q => 
                           n4302);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n7822, Q => 
                           n8978);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n7822, Q => 
                           n7769);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n7822, Q => 
                           n4295);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n7822, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n7822, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n554, Q => n4293);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1843, B => n1844, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1841, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1839, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1837, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1834, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1832, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1830, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1828, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1826, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1824, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1822, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1820, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1818, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1816, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1814, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3036,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => n8793);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => n8792);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => n8791);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => n8790);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => n8789);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => n8788);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => n8787);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => n8786);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => n8785);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => n8784);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => n8783);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => n8782);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => n8781);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => n8780);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1004, S => n8779);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => n14122, 
                           CI => n3026, CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => n8773);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => n14121, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => n14120, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => n14119, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => n14118, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => n14117,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => n14116,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => n14115,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => n14114,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => n14113,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => n14112,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => n14111,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => n14110,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => n14109,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => n8772);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => n14109,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => n8771, S => n8770);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n13855, B => n14108, CI => n14101, CO => n_1005, S 
                           => boothmul_pipelined_i_sum_B_in_3_22_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3030,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => n8765);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => n4018);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => n4017);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => n4016);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => n4015);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => n4014);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => n4013);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => n4012);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => n8764);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => n8763, S => n8762);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n14145, B => n14102, CI => n14094, CO => n4009, S =>
                           n4008);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n14144, B => n14100, CI => n4009, CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n14143, B => boothmul_pipelined_i_sum_B_in_3_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n14142, B => boothmul_pipelined_i_sum_B_in_3_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n13854, B => boothmul_pipelined_i_sum_B_in_3_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1006, S => n4007);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => n4018, 
                           CI => n3029, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => n8757);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => n4017, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => n4016, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => n8755);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => n4015, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => n8754);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => n4014, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => n8753);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => n4013, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => n8752);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => n4012, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => n8751, S => n8750);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n8928, B => n8764, CI => n8751, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => n3996);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n13904, B => n14093, CI => n14086, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => n3995);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n13903, B => n4008, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => n3994);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n13902, B => boothmul_pipelined_i_sum_B_in_4_19_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => n3993);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n13901, B => boothmul_pipelined_i_sum_B_in_4_20_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => n3992);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n13900, B => boothmul_pipelined_i_sum_B_in_4_21_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => n3991, S => n3990);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n13899, B => n4007, CI => n3991, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n13898, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => n8749);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n13861, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1007, S => n8748);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => n8755, 
                           CI => n3028, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => n8744);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => n8754, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => n8753, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => n8742);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => n8752, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => n8741);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           n14249, B => n14087, CI => n14077, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => n8740);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n14248, B => n14085, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => n8739);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n14247, B => n3995, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => n8738);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n14246, B => n3994, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => n8737);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n14245, B => n3993, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => n8736);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n14244, B => n3992, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => n8735);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n14243, B => n3990, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => n8734);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n14242, B => boothmul_pipelined_i_sum_B_in_5_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => n8733, S => n8732);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n14241, B => n8749, CI => n8733, CO => n3974, S => 
                           n3973);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n14240, B => n8748, CI => n3974, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n13897, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => n8731);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n13860, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1008, S => n8730);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => n14078,
                           CI => n3027, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => n8727);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => n14076,
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => n8740, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => n8725);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => n8739, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => n8724);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => n8738, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => n8723);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => n8737, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => n8722);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => n8736, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => n8721);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => n8735, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => n8720);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => n8734, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => n8719);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => n8732, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => n8718);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => n3973, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => n8717);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => n8716, S => n8715);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n14239, B => n14075, CI => n14059, CO => n3958, S =>
                           n3957);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n14238, B => n14074, CI => n3958, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n13896, B => n14074, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => n8714);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n13859, B => n14074, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1009, S => n8713);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => n14068,
                           CI => n3020, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => n8710);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => n14067,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => n8708);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => n14066,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => n8706);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => n14065,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => n8704);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => n14064,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => n8702);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => n14063,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => n8700);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => n14062,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => n8698);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => n14061,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => n8696);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => n14060,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => n8694);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => n14058,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => n8692);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => n3957, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => n8690);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => n8689, S => n8686);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n14237, B => n14057, CI => n14022, CO => n3940, S =>
                           n8685);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n14236, B => n14056, CI => n3940, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => n8683);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           n14235, B => n14056, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => n8682);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           n14234, B => n14056, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => n8681);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           n14234, B => n14056, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1010, S => n8679);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n7822, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n18230, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n554, Q => n4395);
   clk_r_REG7407_S3 : DFFR_X1 port map( D => DATA1(8), CK => clk, RN => rst_BAR
                           , Q => n14469, QN => n18193);
   clk_r_REG7561_S3 : DFFR_X1 port map( D => DATA1(7), CK => clk, RN => rst_BAR
                           , Q => n14467, QN => n16393);
   clk_r_REG7652_S3 : DFFS_X1 port map( D => n1888, CK => clk, SN => rst_BAR, Q
                           => n_1011, QN => n14466);
   clk_r_REG7937_S6 : DFFS_X1 port map( D => n1889, CK => clk, SN => rst_BAR, Q
                           => n18219, QN => n14465);
   clk_r_REG7528_S8 : DFFS_X1 port map( D => n1890, CK => clk, SN => rst_BAR, Q
                           => n_1012, QN => n14464);
   clk_r_REG8347_S3 : DFFS_X1 port map( D => n1891, CK => clk, SN => rst_BAR, Q
                           => n_1013, QN => n14463);
   clk_r_REG8349_S4 : DFFS_X1 port map( D => n14463, CK => clk, SN => rst_BAR, 
                           Q => n14462, QN => n_1014);
   clk_r_REG9901_S7 : DFFS_X1 port map( D => n1892, CK => clk, SN => rst_BAR, Q
                           => n_1015, QN => n14461);
   clk_r_REG10107_S2 : DFFR_X1 port map( D => cin, CK => clk, RN => rst_BAR, Q 
                           => n14460, QN => n_1016);
   clk_r_REG8019_S10 : DFFS_X1 port map( D => n1835, CK => clk, SN => rst_BAR, 
                           Q => n14459, QN => n_1017);
   clk_r_REG7869_S3 : DFFR_X1 port map( D => n13096, CK => clk, RN => rst_BAR, 
                           Q => n18192, QN => n14458);
   clk_r_REG7821_S3 : DFFR_X1 port map( D => n13099, CK => clk, RN => rst_BAR, 
                           Q => n18186, QN => n14457);
   clk_r_REG7820_S3 : DFFS_X1 port map( D => n13099, CK => clk, SN => rst_BAR, 
                           Q => n18180, QN => n14456);
   clk_r_REG7857_S3 : DFFR_X1 port map( D => n9011, CK => clk, RN => rst_BAR, Q
                           => n_1018, QN => n14455);
   clk_r_REG7800_S3 : DFFR_X1 port map( D => n11927, CK => clk, RN => rst_BAR, 
                           Q => n_1019, QN => n14454);
   clk_r_REG7938_S6 : DFFS_X1 port map( D => n1889, CK => clk, SN => rst_BAR, Q
                           => n14453, QN => n18213);
   clk_r_REG7250_S4 : DFFS_X1 port map( D => n1810, CK => clk, SN => rst_BAR, Q
                           => n14452, QN => n_1020);
   clk_r_REG8205_S3 : DFFR_X1 port map( D => DATA1(2), CK => clk, RN => rst_BAR
                           , Q => n_1021, QN => n14451);
   clk_r_REG9374_S5 : DFFS_X1 port map( D => n11946, CK => clk, SN => rst_BAR, 
                           Q => n_1022, QN => n14450);
   clk_r_REG9825_S7 : DFFR_X1 port map( D => DATA1(3), CK => clk, RN => rst_BAR
                           , Q => n18206, QN => n14449);
   clk_r_REG9184_S4 : DFFR_X1 port map( D => n1880, CK => clk, RN => rst_BAR, Q
                           => n14448, QN => n_1023);
   clk_r_REG7840_S3 : DFFR_X1 port map( D => n1883, CK => clk, RN => rst_BAR, Q
                           => n14447, QN => n_1024);
   clk_r_REG7844_S4 : DFFR_X1 port map( D => n1876, CK => clk, RN => rst_BAR, Q
                           => n14446, QN => n_1025);
   clk_r_REG8676_S4 : DFFR_X1 port map( D => n1877, CK => clk, RN => rst_BAR, Q
                           => n14445, QN => n_1026);
   clk_r_REG7846_S4 : DFFS_X1 port map( D => n1874, CK => clk, SN => rst_BAR, Q
                           => n14444, QN => n_1027);
   clk_r_REG7837_S3 : DFFS_X1 port map( D => n1886, CK => clk, SN => rst_BAR, Q
                           => n14443, QN => n_1028);
   clk_r_REG7838_S4 : DFFS_X1 port map( D => n1887, CK => clk, SN => rst_BAR, Q
                           => n14442, QN => n_1029);
   clk_r_REG7848_S3 : DFFS_X1 port map( D => n1871, CK => clk, SN => rst_BAR, Q
                           => n14441, QN => n_1030);
   clk_r_REG7115_S4 : DFFS_X1 port map( D => n1872, CK => clk, SN => rst_BAR, Q
                           => n14440, QN => n_1031);
   clk_r_REG9185_S4 : DFFS_X1 port map( D => n1882, CK => clk, SN => rst_BAR, Q
                           => n14439, QN => n_1032);
   clk_r_REG7529_S8 : DFFS_X1 port map( D => n1890, CK => clk, SN => rst_BAR, Q
                           => n14438, QN => n_1033);
   clk_r_REG7653_S3 : DFFS_X1 port map( D => n1888, CK => clk, SN => rst_BAR, Q
                           => n14437, QN => n18202);
   clk_r_REG7807_S3 : DFFS_X1 port map( D => n13151, CK => clk, SN => rst_BAR, 
                           Q => n_1034, QN => n14436);
   clk_r_REG7812_S3 : DFFR_X1 port map( D => n9020, CK => clk, RN => rst_BAR, Q
                           => n_1035, QN => n14435);
   clk_r_REG7811_S3 : DFFS_X1 port map( D => n9020, CK => clk, SN => rst_BAR, Q
                           => n_1036, QN => n14434);
   clk_r_REG7404_S5 : DFFR_X1 port map( D => n1846, CK => clk, RN => rst_BAR, Q
                           => n14433, QN => n_1037);
   clk_r_REG7307_S4 : DFFS_X1 port map( D => n1864, CK => clk, SN => rst_BAR, Q
                           => n14432, QN => n_1038);
   clk_r_REG7432_S4 : DFFR_X1 port map( D => n1860, CK => clk, RN => rst_BAR, Q
                           => n14431, QN => n_1039);
   clk_r_REG7438_S4 : DFFS_X1 port map( D => n1854, CK => clk, SN => rst_BAR, Q
                           => n14430, QN => n_1040);
   clk_r_REG7161_S4 : DFFR_X1 port map( D => n1878, CK => clk, RN => rst_BAR, Q
                           => n14429, QN => n_1041);
   clk_r_REG7155_S4 : DFFR_X1 port map( D => n1879, CK => clk, RN => rst_BAR, Q
                           => n14428, QN => n_1042);
   clk_r_REG7303_S4 : DFFR_X1 port map( D => n1885, CK => clk, RN => rst_BAR, Q
                           => n14427, QN => n_1043);
   clk_r_REG7038_S4 : DFFS_X1 port map( D => n1873, CK => clk, SN => rst_BAR, Q
                           => n14426, QN => n_1044);
   clk_r_REG7041_S4 : DFFS_X1 port map( D => n1875, CK => clk, SN => rst_BAR, Q
                           => n14425, QN => n_1045);
   clk_r_REG7001_S5 : DFFR_X1 port map( D => n1808, CK => clk, RN => rst_BAR, Q
                           => n14424, QN => n_1046);
   clk_r_REG7422_S4 : DFFS_X1 port map( D => n1858, CK => clk, SN => rst_BAR, Q
                           => n14423, QN => n_1047);
   clk_r_REG7343_S5 : DFFS_X1 port map( D => n16416, CK => clk, SN => rst_BAR, 
                           Q => n14422, QN => n_1048);
   clk_r_REG7335_S5 : DFFR_X1 port map( D => n16415, CK => clk, RN => rst_BAR, 
                           Q => n14421, QN => n_1049);
   clk_r_REG7796_S3 : DFFR_X1 port map( D => n16408, CK => clk, RN => rst_BAR, 
                           Q => n14420, QN => n18177);
   clk_r_REG7953_S3 : DFFR_X1 port map( D => n1868, CK => clk, RN => rst_BAR, Q
                           => n14418, QN => n18212);
   clk_r_REG7761_S3 : DFFS_X1 port map( D => n16400, CK => clk, SN => rst_BAR, 
                           Q => n14417, QN => n18197);
   clk_r_REG7359_S5 : DFFS_X1 port map( D => n1811, CK => clk, SN => rst_BAR, Q
                           => n14416, QN => n_1050);
   clk_r_REG7183_S10 : DFFR_X1 port map( D => n1851, CK => clk, RN => rst_BAR, 
                           Q => n14415, QN => n_1051);
   clk_r_REG7151_S3 : DFFR_X1 port map( D => n1849, CK => clk, RN => rst_BAR, Q
                           => n14414, QN => n_1052);
   clk_r_REG7096_S11 : DFFR_X1 port map( D => n1850, CK => clk, RN => rst_BAR, 
                           Q => n14413, QN => n_1053);
   clk_r_REG7426_S4 : DFFS_X1 port map( D => n1856, CK => clk, SN => rst_BAR, Q
                           => n14412, QN => n_1054);
   clk_r_REG7431_S4 : DFFS_X1 port map( D => n1852, CK => clk, SN => rst_BAR, Q
                           => n14411, QN => n_1055);
   clk_r_REG7437_S4 : DFFS_X1 port map( D => n1854, CK => clk, SN => rst_BAR, Q
                           => n14410, QN => n_1056);
   clk_r_REG7436_S4 : DFFR_X1 port map( D => n1855, CK => clk, RN => rst_BAR, Q
                           => n14409, QN => n_1057);
   clk_r_REG7162_S4 : DFFR_X1 port map( D => n1881, CK => clk, RN => rst_BAR, Q
                           => n14408, QN => n18201);
   clk_r_REG7163_S4 : DFFS_X1 port map( D => n1884, CK => clk, SN => rst_BAR, Q
                           => n14407, QN => n_1058);
   clk_r_REG7433_S4 : DFFR_X1 port map( D => n1859, CK => clk, RN => rst_BAR, Q
                           => n14406, QN => n_1059);
   clk_r_REG7383_S4 : DFFS_X1 port map( D => n1863, CK => clk, SN => rst_BAR, Q
                           => n14405, QN => n_1060);
   clk_r_REG8421_S4 : DFFR_X1 port map( D => n1865, CK => clk, RN => rst_BAR, Q
                           => n14404, QN => n_1061);
   clk_r_REG7767_S3 : DFFR_X1 port map( D => n16401, CK => clk, RN => rst_BAR, 
                           Q => n14403, QN => n18178);
   clk_r_REG7768_S3 : DFFS_X1 port map( D => n16401, CK => clk, SN => rst_BAR, 
                           Q => n14402, QN => n_1062);
   clk_r_REG7759_S3 : DFFS_X1 port map( D => n1901, CK => clk, SN => rst_BAR, Q
                           => n14401, QN => n18189);
   clk_r_REG7776_S3 : DFFS_X1 port map( D => n1902, CK => clk, SN => rst_BAR, Q
                           => n14400, QN => n18190);
   clk_r_REG7539_S4 : DFFR_X1 port map( D => n16418, CK => clk, RN => rst_BAR, 
                           Q => n14399, QN => n_1063);
   clk_r_REG7774_S3 : DFFS_X1 port map( D => n16406, CK => clk, SN => rst_BAR, 
                           Q => n14398, QN => n18215);
   clk_r_REG7782_S3 : DFFR_X1 port map( D => n16403, CK => clk, RN => rst_BAR, 
                           Q => n14397, QN => n18225);
   clk_r_REG7803_S3 : DFFR_X1 port map( D => n11927, CK => clk, RN => rst_BAR, 
                           Q => n14396, QN => n_1064);
   clk_r_REG7770_S3 : DFFR_X1 port map( D => n16412, CK => clk, RN => rst_BAR, 
                           Q => n14395, QN => n18226);
   clk_r_REG7791_S3 : DFFR_X1 port map( D => n16413, CK => clk, RN => rst_BAR, 
                           Q => n14394, QN => n_1065);
   clk_r_REG7831_S3 : DFFR_X1 port map( D => n1898, CK => clk, RN => rst_BAR, Q
                           => n14393, QN => n_1066);
   clk_r_REG7424_S4 : DFFR_X1 port map( D => n1857, CK => clk, RN => rst_BAR, Q
                           => n14392, QN => n_1067);
   clk_r_REG7798_S3 : DFFR_X1 port map( D => n1895, CK => clk, RN => rst_BAR, Q
                           => n14391, QN => n_1068);
   clk_r_REG7860_S3 : DFFR_X1 port map( D => n1899, CK => clk, RN => rst_BAR, Q
                           => n14390, QN => n_1069);
   clk_r_REG7824_S3 : DFFR_X1 port map( D => n1893, CK => clk, RN => rst_BAR, Q
                           => n14389, QN => n18211);
   clk_r_REG7754_S3 : DFFR_X1 port map( D => n16405, CK => clk, RN => rst_BAR, 
                           Q => n14388, QN => n_1070);
   clk_r_REG7753_S3 : DFFS_X1 port map( D => n16405, CK => clk, SN => rst_BAR, 
                           Q => n14387, QN => n_1071);
   clk_r_REG7741_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, Q
                           => n14386, QN => n18208);
   clk_r_REG7793_S3 : DFFS_X1 port map( D => n16407, CK => clk, SN => rst_BAR, 
                           Q => n14385, QN => n_1072);
   clk_r_REG7827_S3 : DFFR_X1 port map( D => n16404, CK => clk, RN => rst_BAR, 
                           Q => n14384, QN => n_1073);
   clk_r_REG7852_S3 : DFFR_X1 port map( D => n1897, CK => clk, RN => rst_BAR, Q
                           => n14383, QN => n_1074);
   clk_r_REG7784_S3 : DFFR_X1 port map( D => n16402, CK => clk, RN => rst_BAR, 
                           Q => n14382, QN => n_1075);
   clk_r_REG7780_S3 : DFFR_X1 port map( D => n1904, CK => clk, RN => rst_BAR, Q
                           => n14381, QN => n18224);
   clk_r_REG7779_S3 : DFFS_X1 port map( D => n1904, CK => clk, SN => rst_BAR, Q
                           => n14380, QN => n18216);
   clk_r_REG7558_S5 : DFFR_X1 port map( D => n1847, CK => clk, RN => rst_BAR, Q
                           => n14379, QN => n_1076);
   clk_r_REG7150_S4 : DFFS_X1 port map( D => n1809, CK => clk, SN => rst_BAR, Q
                           => n14378, QN => n_1077);
   clk_r_REG7789_S3 : DFFR_X1 port map( D => n16409, CK => clk, RN => rst_BAR, 
                           Q => n14377, QN => n_1078);
   clk_r_REG7813_S3 : DFFR_X1 port map( D => n9020, CK => clk, RN => rst_BAR, Q
                           => n14376, QN => n_1079);
   clk_r_REG7870_S3 : DFFR_X1 port map( D => n13096, CK => clk, RN => rst_BAR, 
                           Q => n14375, QN => n_1080);
   clk_r_REG7867_S3 : DFFR_X1 port map( D => n13099, CK => clk, RN => rst_BAR, 
                           Q => n14374, QN => n_1081);
   clk_r_REG7868_S3 : DFFS_X1 port map( D => n13099, CK => clk, SN => rst_BAR, 
                           Q => n14373, QN => n_1082);
   clk_r_REG6942_S4 : DFFS_X1 port map( D => n16417, CK => clk, SN => rst_BAR, 
                           Q => n14372, QN => n_1083);
   clk_r_REG7333_S5 : DFFS_X1 port map( D => n1845, CK => clk, SN => rst_BAR, Q
                           => n_1084, QN => n16410);
   clk_r_REG7070_S6 : DFFS_X1 port map( D => n16391, CK => clk, SN => rst_BAR, 
                           Q => n_1085, QN => n16396);
   clk_r_REG7192_S6 : DFFS_X1 port map( D => n16390, CK => clk, SN => rst_BAR, 
                           Q => n_1086, QN => n16394);
   clk_r_REG7949_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, Q
                           => n14368, QN => n_1087);
   clk_r_REG7856_S3 : DFFR_X1 port map( D => n1899, CK => clk, RN => rst_BAR, Q
                           => n14367, QN => n_1088);
   clk_r_REG7819_S3 : DFFR_X1 port map( D => n1895, CK => clk, RN => rst_BAR, Q
                           => n14366, QN => n_1089);
   clk_r_REG7808_S3 : DFFS_X1 port map( D => n13151, CK => clk, SN => rst_BAR, 
                           Q => n14365, QN => n_1090);
   clk_r_REG7810_S3 : DFFR_X1 port map( D => n1894, CK => clk, RN => rst_BAR, Q
                           => n14364, QN => n_1091);
   clk_r_REG7802_S3 : DFFR_X1 port map( D => n11927, CK => clk, RN => rst_BAR, 
                           Q => n14363, QN => n_1092);
   clk_r_REG7853_S3 : DFFR_X1 port map( D => n1897, CK => clk, RN => rst_BAR, Q
                           => n14362, QN => n_1093);
   clk_r_REG7825_S3 : DFFR_X1 port map( D => n1893, CK => clk, RN => rst_BAR, Q
                           => n14361, QN => n18205);
   clk_r_REG7757_S3 : DFFS_X1 port map( D => n1900, CK => clk, SN => rst_BAR, Q
                           => n14360, QN => n_1094);
   clk_r_REG7871_S3 : DFFR_X1 port map( D => n13096, CK => clk, RN => rst_BAR, 
                           Q => n14359, QN => n_1095);
   clk_r_REG7795_S3 : DFFR_X1 port map( D => n16408, CK => clk, RN => rst_BAR, 
                           Q => n14358, QN => n18228);
   clk_r_REG7858_S3 : DFFR_X1 port map( D => n9011, CK => clk, RN => rst_BAR, Q
                           => n14357, QN => n_1096);
   clk_r_REG7828_S3 : DFFR_X1 port map( D => n16404, CK => clk, RN => rst_BAR, 
                           Q => n14356, QN => n_1097);
   clk_r_REG8160_S7 : DFFS_X1 port map( D => n1814, CK => clk, SN => rst_BAR, Q
                           => n14355, QN => n_1098);
   clk_r_REG8161_S8 : DFFS_X1 port map( D => n14355, CK => clk, SN => rst_BAR, 
                           Q => n_1099, QN => n16414);
   clk_r_REG9903_S9 : DFFS_X1 port map( D => n1844, CK => clk, SN => rst_BAR, Q
                           => n14353, QN => n_1100);
   clk_r_REG9904_S10 : DFFS_X1 port map( D => n14353, CK => clk, SN => rst_BAR,
                           Q => n14352, QN => n_1101);
   clk_r_REG7950_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, Q
                           => n14351, QN => n_1102);
   clk_r_REG7763_S3 : DFFR_X1 port map( D => n1900, CK => clk, RN => rst_BAR, Q
                           => n14350, QN => n_1103);
   clk_r_REG7815_S3 : DFFR_X1 port map( D => n9020, CK => clk, RN => rst_BAR, Q
                           => n14349, QN => n_1104);
   clk_r_REG7829_S3 : DFFR_X1 port map( D => n16404, CK => clk, RN => rst_BAR, 
                           Q => n14348, QN => n_1105);
   clk_r_REG7771_S3 : DFFR_X1 port map( D => n16412, CK => clk, RN => rst_BAR, 
                           Q => n14347, QN => n_1106);
   clk_r_REG7952_S3 : DFFR_X1 port map( D => n1868, CK => clk, RN => rst_BAR, Q
                           => n14346, QN => n_1107);
   clk_r_REG7762_S3 : DFFS_X1 port map( D => n16400, CK => clk, SN => rst_BAR, 
                           Q => n14345, QN => n_1108);
   clk_r_REG7805_S3 : DFFR_X1 port map( D => n11927, CK => clk, RN => rst_BAR, 
                           Q => n14344, QN => n_1109);
   clk_r_REG7752_S3 : DFFR_X1 port map( D => n16405, CK => clk, RN => rst_BAR, 
                           Q => n14343, QN => n18227);
   clk_r_REG7773_S3 : DFFR_X1 port map( D => n16406, CK => clk, RN => rst_BAR, 
                           Q => n14342, QN => n18203);
   clk_r_REG7834_S3 : DFFR_X1 port map( D => n1898, CK => clk, RN => rst_BAR, Q
                           => n14341, QN => n_1110);
   clk_r_REG7854_S3 : DFFR_X1 port map( D => n1897, CK => clk, RN => rst_BAR, Q
                           => n14340, QN => n_1111);
   clk_r_REG7823_S3 : DFFR_X1 port map( D => n1893, CK => clk, RN => rst_BAR, Q
                           => n14339, QN => n18184);
   clk_r_REG9375_S5 : DFFS_X1 port map( D => n11946, CK => clk, SN => rst_BAR, 
                           Q => n14338, QN => n_1112);
   clk_r_REG7416_S4 : DFFR_X1 port map( D => n1853, CK => clk, RN => rst_BAR, Q
                           => n14337, QN => n_1113);
   clk_r_REG8206_S3 : DFFR_X1 port map( D => DATA1(2), CK => clk, RN => rst_BAR
                           , Q => n14336, QN => n_1114);
   clk_r_REG10254_S7 : DFFR_X1 port map( D => n1870, CK => clk, RN => rst_BAR, 
                           Q => n14335, QN => n_1115);
   clk_r_REG7818_S3 : DFFS_X1 port map( D => n13151, CK => clk, SN => rst_BAR, 
                           Q => n14334, QN => n18204);
   clk_r_REG7816_S3 : DFFR_X1 port map( D => n1894, CK => clk, RN => rst_BAR, Q
                           => n14333, QN => n_1116);
   clk_r_REG7764_S3 : DFFS_X1 port map( D => n1900, CK => clk, SN => rst_BAR, Q
                           => n14332, QN => n_1117);
   clk_r_REG7859_S3 : DFFR_X1 port map( D => n9011, CK => clk, RN => rst_BAR, Q
                           => n14331, QN => n18198);
   clk_r_REG7787_S3 : DFFS_X1 port map( D => n1903, CK => clk, SN => rst_BAR, Q
                           => n14330, QN => n_1118);
   clk_r_REG9902_S7 : DFFS_X1 port map( D => n1892, CK => clk, SN => rst_BAR, Q
                           => n14329, QN => n_1119);
   clk_r_REG8348_S3 : DFFS_X1 port map( D => n1891, CK => clk, SN => rst_BAR, Q
                           => n14328, QN => n18194);
   clk_r_REG8207_S3 : DFFR_X1 port map( D => DATA1(2), CK => clk, RN => rst_BAR
                           , Q => n14327, QN => n_1120);
   clk_r_REG9826_S7 : DFFR_X1 port map( D => DATA1(3), CK => clk, RN => rst_BAR
                           , Q => n14326, QN => n_1121);
   clk_r_REG7269_S5 : DFFS_X1 port map( D => n1816, CK => clk, SN => rst_BAR, Q
                           => n_1122, QN => n14325);
   clk_r_REG7299_S6 : DFFR_X1 port map( D => n14325, CK => clk, RN => rst_BAR, 
                           Q => n14324, QN => n_1123);
   clk_r_REG8173_S8 : DFFS_X1 port map( D => n1818, CK => clk, SN => rst_BAR, Q
                           => n_1124, QN => n14323);
   clk_r_REG8174_S9 : DFFR_X1 port map( D => n14323, CK => clk, RN => rst_BAR, 
                           Q => n14322, QN => n_1125);
   clk_r_REG8041_S8 : DFFS_X1 port map( D => n1820, CK => clk, SN => rst_BAR, Q
                           => n_1126, QN => n14321);
   clk_r_REG8042_S9 : DFFR_X1 port map( D => n14321, CK => clk, RN => rst_BAR, 
                           Q => n14320, QN => n_1127);
   clk_r_REG8033_S8 : DFFS_X1 port map( D => n1822, CK => clk, SN => rst_BAR, Q
                           => n_1128, QN => n14319);
   clk_r_REG8034_S9 : DFFR_X1 port map( D => n14319, CK => clk, RN => rst_BAR, 
                           Q => n14318, QN => n_1129);
   clk_r_REG7517_S9 : DFFS_X1 port map( D => n1824, CK => clk, SN => rst_BAR, Q
                           => n_1130, QN => n14317);
   clk_r_REG7518_S10 : DFFR_X1 port map( D => n14317, CK => clk, RN => rst_BAR,
                           Q => n14316, QN => n_1131);
   clk_r_REG7368_S5 : DFFS_X1 port map( D => n1826, CK => clk, SN => rst_BAR, Q
                           => n_1132, QN => n14315);
   clk_r_REG7381_S6 : DFFR_X1 port map( D => n14315, CK => clk, RN => rst_BAR, 
                           Q => n14314, QN => n_1133);
   clk_r_REG7439_S5 : DFFS_X1 port map( D => n1828, CK => clk, SN => rst_BAR, Q
                           => n_1134, QN => n14313);
   clk_r_REG7442_S6 : DFFR_X1 port map( D => n14313, CK => clk, RN => rst_BAR, 
                           Q => n14312, QN => n_1135);
   clk_r_REG7562_S5 : DFFS_X1 port map( D => n1830, CK => clk, SN => rst_BAR, Q
                           => n_1136, QN => n14311);
   clk_r_REG7566_S6 : DFFR_X1 port map( D => n14311, CK => clk, RN => rst_BAR, 
                           Q => n14310, QN => n_1137);
   clk_r_REG7654_S5 : DFFS_X1 port map( D => n1832, CK => clk, SN => rst_BAR, Q
                           => n_1138, QN => n14309);
   clk_r_REG7658_S6 : DFFR_X1 port map( D => n14309, CK => clk, RN => rst_BAR, 
                           Q => n14308, QN => n_1139);
   clk_r_REG7939_S8 : DFFS_X1 port map( D => n1834, CK => clk, SN => rst_BAR, Q
                           => n_1140, QN => n14307);
   clk_r_REG7943_S9 : DFFR_X1 port map( D => n14307, CK => clk, RN => rst_BAR, 
                           Q => n14306, QN => n_1141);
   clk_r_REG8017_S10 : DFFS_X1 port map( D => n1837, CK => clk, SN => rst_BAR, 
                           Q => n_1142, QN => n14305);
   clk_r_REG8026_S11 : DFFR_X1 port map( D => n14305, CK => clk, RN => rst_BAR,
                           Q => n14304, QN => n_1143);
   clk_r_REG9827_S9 : DFFS_X1 port map( D => n1839, CK => clk, SN => rst_BAR, Q
                           => n_1144, QN => n14303);
   clk_r_REG9828_S10 : DFFR_X1 port map( D => n14303, CK => clk, RN => rst_BAR,
                           Q => n14302, QN => n_1145);
   clk_r_REG8208_S5 : DFFS_X1 port map( D => n1841, CK => clk, SN => rst_BAR, Q
                           => n_1146, QN => n14301);
   clk_r_REG8213_S6 : DFFR_X1 port map( D => n14301, CK => clk, RN => rst_BAR, 
                           Q => n14300, QN => n_1147);
   clk_r_REG8350_S5 : DFFS_X1 port map( D => n1843, CK => clk, SN => rst_BAR, Q
                           => n_1148, QN => n14299);
   clk_r_REG8353_S6 : DFFR_X1 port map( D => n14299, CK => clk, RN => rst_BAR, 
                           Q => n14298, QN => n_1149);
   clk_r_REG7241_S4 : DFFR_X1 port map( D => n13182, CK => clk, RN => rst_BAR, 
                           Q => n14297, QN => n_1150);
   clk_r_REG7242_S5 : DFFR_X1 port map( D => n14297, CK => clk, RN => rst_BAR, 
                           Q => n14296, QN => n_1151);
   clk_r_REG7243_S6 : DFFR_X1 port map( D => n14296, CK => clk, RN => rst_BAR, 
                           Q => n18199, QN => n16389);
   clk_r_REG7260_S4 : DFFR_X1 port map( D => n8990, CK => clk, RN => rst_BAR, Q
                           => n14294, QN => n_1152);
   clk_r_REG7261_S5 : DFFR_X1 port map( D => n14294, CK => clk, RN => rst_BAR, 
                           Q => n14293, QN => n_1153);
   clk_r_REG7262_S6 : DFFR_X1 port map( D => n14293, CK => clk, RN => rst_BAR, 
                           Q => n14292, QN => n_1154);
   clk_r_REG7190_S4 : DFFR_X1 port map( D => n13175, CK => clk, RN => rst_BAR, 
                           Q => n14291, QN => n_1155);
   clk_r_REG7191_S5 : DFFR_X1 port map( D => n14291, CK => clk, RN => rst_BAR, 
                           Q => n14290, QN => n16390);
   clk_r_REG7172_S4 : DFFR_X1 port map( D => n8984, CK => clk, RN => rst_BAR, Q
                           => n14289, QN => n_1156);
   clk_r_REG7173_S5 : DFFR_X1 port map( D => n14289, CK => clk, RN => rst_BAR, 
                           Q => n14288, QN => n_1157);
   clk_r_REG7069_S5 : DFFR_X1 port map( D => n13174, CK => clk, RN => rst_BAR, 
                           Q => n14287, QN => n16391);
   clk_r_REG7050_S5 : DFFR_X1 port map( D => n8980, CK => clk, RN => rst_BAR, Q
                           => n14286, QN => n_1158);
   clk_r_REG7555_S5 : DFFS_X1 port map( D => n8814, CK => clk, SN => rst_BAR, Q
                           => n14282, QN => n_1159);
   clk_r_REG7556_S5 : DFFS_X1 port map( D => n8929, CK => clk, SN => rst_BAR, Q
                           => n14281, QN => n_1160);
   clk_r_REG7297_S5 : DFFS_X1 port map( D => n1812, CK => clk, SN => rst_BAR, Q
                           => n_1161, QN => n14280);
   clk_r_REG7298_S6 : DFFR_X1 port map( D => n14280, CK => clk, RN => rst_BAR, 
                           Q => n14279, QN => n_1162);
   clk_r_REG7251_S4 : DFFR_X1 port map( D => n8943, CK => clk, RN => rst_BAR, Q
                           => n14278, QN => n_1163);
   clk_r_REG10108_S3 : DFFR_X1 port map( D => n1866, CK => clk, RN => rst_BAR, 
                           Q => n_1164, QN => n14277);
   clk_r_REG7951_S3 : DFFR_X1 port map( D => n1868, CK => clk, RN => rst_BAR, Q
                           => n18210, QN => n14276);
   clk_r_REG7739_S3 : DFFR_X1 port map( D => n1869, CK => clk, RN => rst_BAR, Q
                           => n18179, QN => n14275);
   clk_r_REG7809_S3 : DFFR_X1 port map( D => n1894, CK => clk, RN => rst_BAR, Q
                           => n_1165, QN => n14274);
   clk_r_REG7778_S3 : DFFS_X1 port map( D => n11755, CK => clk, SN => rst_BAR, 
                           Q => n14273, QN => n_1166);
   clk_r_REG7648_S4 : DFFS_X1 port map( D => n8957, CK => clk, SN => rst_BAR, Q
                           => n14272, QN => n_1167);
   clk_r_REG8203_S4 : DFFS_X1 port map( D => n8956, CK => clk, SN => rst_BAR, Q
                           => n14271, QN => n_1168);
   clk_r_REG7737_S3 : DFFS_X1 port map( D => n8626, CK => clk, SN => rst_BAR, Q
                           => n14270, QN => n_1169);
   clk_r_REG7000_S5 : DFFR_X1 port map( D => n12158, CK => clk, RN => rst_BAR, 
                           Q => n14269, QN => n_1170);
   clk_r_REG7015_S4 : DFFS_X1 port map( D => n12255, CK => clk, SN => rst_BAR, 
                           Q => n14268, QN => n_1171);
   clk_r_REG6962_S5 : DFFS_X1 port map( D => n8946, CK => clk, SN => rst_BAR, Q
                           => n14267, QN => n_1172);
   clk_r_REG7110_S5 : DFFS_X1 port map( D => n8945, CK => clk, SN => rst_BAR, Q
                           => n14266, QN => n_1173);
   clk_r_REG7201_S10 : DFFS_X1 port map( D => n8944, CK => clk, SN => rst_BAR, 
                           Q => n14265, QN => n_1174);
   clk_r_REG7024_S4 : DFFR_X1 port map( D => n12292, CK => clk, RN => rst_BAR, 
                           Q => n14264, QN => n_1175);
   clk_r_REG6948_S10 : DFFS_X1 port map( D => n12325, CK => clk, SN => rst_BAR,
                           Q => n14263, QN => n_1176);
   clk_r_REG7129_S4 : DFFS_X1 port map( D => n12400, CK => clk, SN => rst_BAR, 
                           Q => n14262, QN => n_1177);
   clk_r_REG8175_S7 : DFFS_X1 port map( D => n12474, CK => clk, SN => rst_BAR, 
                           Q => n14261, QN => n_1178);
   clk_r_REG7056_S11 : DFFS_X1 port map( D => n8940, CK => clk, SN => rst_BAR, 
                           Q => n14260, QN => n_1179);
   clk_r_REG7738_S3 : DFFS_X1 port map( D => n12754, CK => clk, SN => rst_BAR, 
                           Q => n14259, QN => n_1180);
   clk_r_REG6914_S4 : DFFR_X1 port map( D => n8933, CK => clk, RN => rst_BAR, Q
                           => n14258, QN => n_1181);
   clk_r_REG6915_S5 : DFFR_X1 port map( D => n14258, CK => clk, RN => rst_BAR, 
                           Q => n14257, QN => n_1182);
   clk_r_REG6916_S6 : DFFR_X1 port map( D => n14257, CK => clk, RN => rst_BAR, 
                           Q => n14256, QN => n_1183);
   clk_r_REG6917_S7 : DFFR_X1 port map( D => n14256, CK => clk, RN => rst_BAR, 
                           Q => n14255, QN => n_1184);
   clk_r_REG6918_S8 : DFFR_X1 port map( D => n14255, CK => clk, RN => rst_BAR, 
                           Q => n14254, QN => n_1185);
   clk_r_REG6919_S9 : DFFR_X1 port map( D => n14254, CK => clk, RN => rst_BAR, 
                           Q => n14253, QN => n_1186);
   clk_r_REG7733_S4 : DFFS_X1 port map( D => n8932, CK => clk, SN => rst_BAR, Q
                           => n14252, QN => n_1187);
   clk_r_REG7334_S5 : DFFR_X1 port map( D => n16415, CK => clk, RN => rst_BAR, 
                           Q => n_1188, QN => n14250);
   clk_r_REG7353_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_15_port, CK => clk, 
                           RN => rst_BAR, Q => n14249, QN => n_1189);
   clk_r_REG7352_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_16_port, CK => clk, 
                           RN => rst_BAR, Q => n14248, QN => n_1190);
   clk_r_REG7351_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_17_port, CK => clk, 
                           RN => rst_BAR, Q => n14247, QN => n_1191);
   clk_r_REG7350_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_18_port, CK => clk, 
                           RN => rst_BAR, Q => n14246, QN => n_1192);
   clk_r_REG7349_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_19_port, CK => clk, 
                           RN => rst_BAR, Q => n14245, QN => n_1193);
   clk_r_REG7348_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_20_port, CK => clk, 
                           RN => rst_BAR, Q => n14244, QN => n_1194);
   clk_r_REG7347_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_21_port, CK => clk, 
                           RN => rst_BAR, Q => n14243, QN => n_1195);
   clk_r_REG7346_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_22_port, CK => clk, 
                           RN => rst_BAR, Q => n14242, QN => n_1196);
   clk_r_REG7345_S6 : DFFR_X1 port map( D => n8920, CK => clk, RN => rst_BAR, Q
                           => n14241, QN => n_1197);
   clk_r_REG7097_S6 : DFFR_X1 port map( D => n8919, CK => clk, RN => rst_BAR, Q
                           => n14240, QN => n_1198);
   clk_r_REG7196_S6 : DFFR_X1 port map( D => n8917, CK => clk, RN => rst_BAR, Q
                           => n14239, QN => n_1199);
   clk_r_REG7195_S6 : DFFR_X1 port map( D => n8916, CK => clk, RN => rst_BAR, Q
                           => n14238, QN => n_1200);
   clk_r_REG7247_S7 : DFFR_X1 port map( D => n8914, CK => clk, RN => rst_BAR, Q
                           => n14237, QN => n_1201);
   clk_r_REG7246_S7 : DFFR_X1 port map( D => n8913, CK => clk, RN => rst_BAR, Q
                           => n14236, QN => n_1202);
   clk_r_REG7245_S7 : DFFR_X1 port map( D => n8912, CK => clk, RN => rst_BAR, Q
                           => n14235, QN => n_1203);
   clk_r_REG7244_S7 : DFFR_X1 port map( D => n8911, CK => clk, RN => rst_BAR, Q
                           => n14234, QN => n_1204);
   clk_r_REG7552_S5 : DFFR_X1 port map( D => n16419, CK => clk, RN => rst_BAR, 
                           Q => n_1205, QN => n14233);
   clk_r_REG7792_S3 : DFFS_X1 port map( D => n16407, CK => clk, SN => rst_BAR, 
                           Q => n18220, QN => n14232);
   clk_r_REG7786_S3 : DFFR_X1 port map( D => n1903, CK => clk, RN => rst_BAR, Q
                           => n_1206, QN => n14230);
   clk_r_REG7785_S3 : DFFS_X1 port map( D => n1903, CK => clk, SN => rst_BAR, Q
                           => n_1207, QN => n14229);
   clk_r_REG7790_S3 : DFFR_X1 port map( D => n16413, CK => clk, RN => rst_BAR, 
                           Q => n18207, QN => n14227);
   clk_r_REG7830_S3 : DFFR_X1 port map( D => n1898, CK => clk, RN => rst_BAR, Q
                           => n18185, QN => n14226);
   clk_r_REG7769_S3 : DFFR_X1 port map( D => n16412, CK => clk, RN => rst_BAR, 
                           Q => n18176, QN => n14225);
   clk_r_REG7538_S4 : DFFR_X1 port map( D => n16418, CK => clk, RN => rst_BAR, 
                           Q => n_1208, QN => n14224);
   clk_r_REG7788_S3 : DFFR_X1 port map( D => n16409, CK => clk, RN => rst_BAR, 
                           Q => n_1209, QN => n14222);
   clk_r_REG7756_S3 : DFFR_X1 port map( D => n1900, CK => clk, RN => rst_BAR, Q
                           => n18200, QN => n14221);
   clk_r_REG7755_S3 : DFFS_X1 port map( D => n1900, CK => clk, SN => rst_BAR, Q
                           => n18218, QN => n14220);
   clk_r_REG8351_S5 : DFFS_X1 port map( D => n1842, CK => clk, SN => rst_BAR, Q
                           => n_1210, QN => n14219);
   clk_r_REG8352_S6 : DFFR_X1 port map( D => n14219, CK => clk, RN => rst_BAR, 
                           Q => n14218, QN => n_1211);
   clk_r_REG8209_S5 : DFFS_X1 port map( D => n1840, CK => clk, SN => rst_BAR, Q
                           => n_1212, QN => n14217);
   clk_r_REG8210_S6 : DFFR_X1 port map( D => n14217, CK => clk, RN => rst_BAR, 
                           Q => n14216, QN => n_1213);
   clk_r_REG8211_S5 : DFFS_X1 port map( D => n1838, CK => clk, SN => rst_BAR, Q
                           => n_1214, QN => n14215);
   clk_r_REG8212_S6 : DFFR_X1 port map( D => n14215, CK => clk, RN => rst_BAR, 
                           Q => n14214, QN => n_1215);
   clk_r_REG8018_S10 : DFFS_X1 port map( D => n1836, CK => clk, SN => rst_BAR, 
                           Q => n_1216, QN => n14213);
   clk_r_REG8025_S11 : DFFR_X1 port map( D => n14213, CK => clk, RN => rst_BAR,
                           Q => n14212, QN => n_1217);
   clk_r_REG7940_S8 : DFFS_X1 port map( D => n1833, CK => clk, SN => rst_BAR, Q
                           => n_1218, QN => n14211);
   clk_r_REG7942_S9 : DFFR_X1 port map( D => n14211, CK => clk, RN => rst_BAR, 
                           Q => n14210, QN => n_1219);
   clk_r_REG7655_S5 : DFFS_X1 port map( D => n1831, CK => clk, SN => rst_BAR, Q
                           => n_1220, QN => n14209);
   clk_r_REG7657_S6 : DFFR_X1 port map( D => n14209, CK => clk, RN => rst_BAR, 
                           Q => n14208, QN => n_1221);
   clk_r_REG7563_S5 : DFFS_X1 port map( D => n1829, CK => clk, SN => rst_BAR, Q
                           => n_1222, QN => n14207);
   clk_r_REG7565_S6 : DFFR_X1 port map( D => n14207, CK => clk, RN => rst_BAR, 
                           Q => n14206, QN => n_1223);
   clk_r_REG7440_S5 : DFFS_X1 port map( D => n1827, CK => clk, SN => rst_BAR, Q
                           => n_1224, QN => n14205);
   clk_r_REG7441_S6 : DFFR_X1 port map( D => n14205, CK => clk, RN => rst_BAR, 
                           Q => n14204, QN => n_1225);
   clk_r_REG7369_S5 : DFFS_X1 port map( D => n1825, CK => clk, SN => rst_BAR, Q
                           => n_1226, QN => n14203);
   clk_r_REG7370_S6 : DFFR_X1 port map( D => n14203, CK => clk, RN => rst_BAR, 
                           Q => n14202, QN => n_1227);
   clk_r_REG7371_S5 : DFFS_X1 port map( D => n1823, CK => clk, SN => rst_BAR, Q
                           => n_1228, QN => n14201);
   clk_r_REG7372_S6 : DFFR_X1 port map( D => n14201, CK => clk, RN => rst_BAR, 
                           Q => n14200, QN => n_1229);
   clk_r_REG7373_S5 : DFFS_X1 port map( D => n1821, CK => clk, SN => rst_BAR, Q
                           => n_1230, QN => n14199);
   clk_r_REG7375_S6 : DFFR_X1 port map( D => n14199, CK => clk, RN => rst_BAR, 
                           Q => n14198, QN => n_1231);
   clk_r_REG7376_S5 : DFFS_X1 port map( D => n1819, CK => clk, SN => rst_BAR, Q
                           => n_1232, QN => n14197);
   clk_r_REG7378_S6 : DFFR_X1 port map( D => n14197, CK => clk, RN => rst_BAR, 
                           Q => n14196, QN => n_1233);
   clk_r_REG7379_S5 : DFFS_X1 port map( D => n1817, CK => clk, SN => rst_BAR, Q
                           => n_1234, QN => n14195);
   clk_r_REG7380_S6 : DFFR_X1 port map( D => n14195, CK => clk, RN => rst_BAR, 
                           Q => n14194, QN => n_1235);
   clk_r_REG7270_S5 : DFFS_X1 port map( D => n1815, CK => clk, SN => rst_BAR, Q
                           => n_1236, QN => n14193);
   clk_r_REG7292_S6 : DFFR_X1 port map( D => n14193, CK => clk, RN => rst_BAR, 
                           Q => n14192, QN => n_1237);
   clk_r_REG7293_S5 : DFFS_X1 port map( D => n1813, CK => clk, SN => rst_BAR, Q
                           => n_1238, QN => n14191);
   clk_r_REG7296_S6 : DFFR_X1 port map( D => n14191, CK => clk, RN => rst_BAR, 
                           Q => n14190, QN => n_1239);
   clk_r_REG7647_S4 : DFFR_X1 port map( D => n1848, CK => clk, RN => rst_BAR, Q
                           => n_1240, QN => n14189);
   clk_r_REG7855_S3 : DFFR_X1 port map( D => n1899, CK => clk, RN => rst_BAR, Q
                           => n18195, QN => n14188);
   clk_r_REG7797_S3 : DFFR_X1 port map( D => n1895, CK => clk, RN => rst_BAR, Q
                           => n_1241, QN => n14187);
   clk_r_REG7799_S3 : DFFS_X1 port map( D => n1896, CK => clk, SN => rst_BAR, Q
                           => n_1242, QN => n14186);
   clk_r_REG7748_S4 : DFFS_X1 port map( D => n1429, CK => clk, SN => rst_BAR, Q
                           => n14185, QN => n_1243);
   clk_r_REG8073_S6 : DFFR_X1 port map( D => n8892, CK => clk, RN => rst_BAR, Q
                           => n14184, QN => n_1244);
   clk_r_REG7734_S4 : DFFS_X1 port map( D => n2808, CK => clk, SN => rst_BAR, Q
                           => n14183, QN => n_1245);
   clk_r_REG7735_S4 : DFFR_X1 port map( D => n8887, CK => clk, RN => rst_BAR, Q
                           => n14182, QN => n_1246);
   clk_r_REG7403_S5 : DFFR_X1 port map( D => n1846, CK => clk, RN => rst_BAR, Q
                           => n_1247, QN => n14181);
   clk_r_REG7391_S5 : DFFR_X1 port map( D => n8875, CK => clk, RN => rst_BAR, Q
                           => n14180, QN => n_1248);
   clk_r_REG7392_S6 : DFFR_X1 port map( D => n14180, CK => clk, RN => rst_BAR, 
                           Q => n14179, QN => n_1249);
   clk_r_REG7393_S7 : DFFR_X1 port map( D => n14179, CK => clk, RN => rst_BAR, 
                           Q => n14178, QN => n_1250);
   clk_r_REG7394_S8 : DFFR_X1 port map( D => n14178, CK => clk, RN => rst_BAR, 
                           Q => n14177, QN => n_1251);
   clk_r_REG7395_S9 : DFFR_X1 port map( D => n14177, CK => clk, RN => rst_BAR, 
                           Q => n14176, QN => n_1252);
   clk_r_REG8193_S4 : DFFR_X1 port map( D => n8861, CK => clk, RN => rst_BAR, Q
                           => n14175, QN => n_1253);
   clk_r_REG8194_S5 : DFFR_X1 port map( D => n14175, CK => clk, RN => rst_BAR, 
                           Q => n14174, QN => n_1254);
   clk_r_REG8195_S6 : DFFR_X1 port map( D => n14174, CK => clk, RN => rst_BAR, 
                           Q => n14173, QN => n_1255);
   clk_r_REG8196_S7 : DFFR_X1 port map( D => n14173, CK => clk, RN => rst_BAR, 
                           Q => n14172, QN => n_1256);
   clk_r_REG8197_S8 : DFFR_X1 port map( D => n14172, CK => clk, RN => rst_BAR, 
                           Q => n14171, QN => n_1257);
   clk_r_REG8198_S9 : DFFR_X1 port map( D => n14171, CK => clk, RN => rst_BAR, 
                           Q => n14170, QN => n_1258);
   clk_r_REG7365_S4 : DFFS_X1 port map( D => n8859, CK => clk, SN => rst_BAR, Q
                           => n14169, QN => n_1259);
   clk_r_REG7427_S4 : DFFS_X1 port map( D => n11714, CK => clk, SN => rst_BAR, 
                           Q => n14168, QN => n_1260);
   clk_r_REG6991_S5 : DFFS_X1 port map( D => n8847, CK => clk, SN => rst_BAR, Q
                           => n14167, QN => n_1261);
   clk_r_REG7160_S4 : DFFR_X1 port map( D => n1878, CK => clk, RN => rst_BAR, Q
                           => n_1262, QN => n14166);
   clk_r_REG7002_S5 : DFFS_X1 port map( D => n12151, CK => clk, SN => rst_BAR, 
                           Q => n14165, QN => n_1263);
   clk_r_REG6992_S5 : DFFR_X1 port map( D => n12212, CK => clk, RN => rst_BAR, 
                           Q => n14164, QN => n_1264);
   clk_r_REG7013_S4 : DFFS_X1 port map( D => n12230, CK => clk, SN => rst_BAR, 
                           Q => n14163, QN => n_1265);
   clk_r_REG8123_S4 : DFFS_X1 port map( D => n8838, CK => clk, SN => rst_BAR, Q
                           => n14162, QN => n_1266);
   clk_r_REG7861_S3 : DFFS_X1 port map( D => n12263, CK => clk, SN => rst_BAR, 
                           Q => n14161, QN => n_1267);
   clk_r_REG7111_S5 : DFFS_X1 port map( D => n8837, CK => clk, SN => rst_BAR, Q
                           => n14160, QN => n_1268);
   clk_r_REG7031_S3 : DFFS_X1 port map( D => n8834, CK => clk, SN => rst_BAR, Q
                           => n14159, QN => n_1269);
   clk_r_REG7023_S4 : DFFR_X1 port map( D => n8587, CK => clk, RN => rst_BAR, Q
                           => n14158, QN => n_1270);
   clk_r_REG7016_S4 : DFFR_X1 port map( D => n12306, CK => clk, RN => rst_BAR, 
                           Q => n14157, QN => n_1271);
   clk_r_REG7850_S3 : DFFS_X1 port map( D => n12313, CK => clk, SN => rst_BAR, 
                           Q => n_1272, QN => n18229);
   clk_r_REG7865_S3 : DFFR_X1 port map( D => n8832, CK => clk, RN => rst_BAR, Q
                           => n14155, QN => n_1273);
   clk_r_REG7866_S3 : DFFS_X1 port map( D => n8831, CK => clk, SN => rst_BAR, Q
                           => n14154, QN => n_1274);
   clk_r_REG8145_S6 : DFFS_X1 port map( D => n8830, CK => clk, SN => rst_BAR, Q
                           => n14153, QN => n_1275);
   clk_r_REG8153_S3 : DFFS_X1 port map( D => n8828, CK => clk, SN => rst_BAR, Q
                           => n14152, QN => n_1276);
   clk_r_REG7249_S4 : DFFS_X1 port map( D => n12423, CK => clk, SN => rst_BAR, 
                           Q => n14151, QN => n_1277);
   clk_r_REG7266_S4 : DFFR_X1 port map( D => n8826, CK => clk, RN => rst_BAR, Q
                           => n14150, QN => n_1278);
   clk_r_REG7361_S5 : DFFR_X1 port map( D => n8821, CK => clk, RN => rst_BAR, Q
                           => n14149, QN => n_1279);
   clk_r_REG7357_S5 : DFFR_X1 port map( D => n8566, CK => clk, RN => rst_BAR, Q
                           => n14148, QN => n_1280);
   clk_r_REG7356_S5 : DFFS_X1 port map( D => n8820, CK => clk, SN => rst_BAR, Q
                           => n14147, QN => n_1281);
   clk_r_REG7418_S4 : DFFS_X1 port map( D => n12527, CK => clk, SN => rst_BAR, 
                           Q => n14146, QN => n_1282);
   clk_r_REG7374_S5 : DFFR_X1 port map( D => n8813, CK => clk, RN => rst_BAR, Q
                           => n14145, QN => n_1283);
   clk_r_REG7377_S5 : DFFR_X1 port map( D => n8812, CK => clk, RN => rst_BAR, Q
                           => n14144, QN => n_1284);
   clk_r_REG7291_S5 : DFFR_X1 port map( D => n8811, CK => clk, RN => rst_BAR, Q
                           => n14143, QN => n_1285);
   clk_r_REG7290_S5 : DFFR_X1 port map( D => n8810, CK => clk, RN => rst_BAR, Q
                           => n14142, QN => n_1286);
   clk_r_REG8200_S4 : DFFR_X1 port map( D => n8800, CK => clk, RN => rst_BAR, Q
                           => n14140, QN => n_1287);
   clk_r_REG7783_S3 : DFFR_X1 port map( D => n16402, CK => clk, RN => rst_BAR, 
                           Q => n18191, QN => n14139);
   clk_r_REG7781_S3 : DFFR_X1 port map( D => n16403, CK => clk, RN => rst_BAR, 
                           Q => n18214, QN => n14138);
   clk_r_REG7772_S3 : DFFR_X1 port map( D => n16406, CK => clk, RN => rst_BAR, 
                           Q => n18217, QN => n14137);
   clk_r_REG7751_S3 : DFFR_X1 port map( D => n16405, CK => clk, RN => rst_BAR, 
                           Q => n18209, QN => n14136);
   clk_r_REG7750_S3 : DFFS_X1 port map( D => n16405, CK => clk, SN => rst_BAR, 
                           Q => n18222, QN => n14135);
   clk_r_REG7777_S3 : DFFR_X1 port map( D => n1904, CK => clk, RN => rst_BAR, Q
                           => n_1288, QN => n14133);
   clk_r_REG6940_S4 : DFFS_X1 port map( D => n8900, CK => clk, SN => rst_BAR, Q
                           => n14132, QN => n_1289);
   clk_r_REG7775_S3 : DFFS_X1 port map( D => n1902, CK => clk, SN => rst_BAR, Q
                           => n_1290, QN => n14131);
   clk_r_REG7822_S3 : DFFR_X1 port map( D => n1893, CK => clk, RN => rst_BAR, Q
                           => n18196, QN => n14130);
   clk_r_REG7758_S3 : DFFS_X1 port map( D => n1901, CK => clk, SN => rst_BAR, Q
                           => n18183, QN => n14129);
   clk_r_REG8186_S4 : DFFR_X1 port map( D => n8793, CK => clk, RN => rst_BAR, Q
                           => n14128, QN => n_1291);
   clk_r_REG8187_S5 : DFFR_X1 port map( D => n14128, CK => clk, RN => rst_BAR, 
                           Q => n14127, QN => n_1292);
   clk_r_REG8188_S6 : DFFR_X1 port map( D => n14127, CK => clk, RN => rst_BAR, 
                           Q => n14126, QN => n_1293);
   clk_r_REG8189_S7 : DFFR_X1 port map( D => n14126, CK => clk, RN => rst_BAR, 
                           Q => n14125, QN => n_1294);
   clk_r_REG8190_S8 : DFFR_X1 port map( D => n14125, CK => clk, RN => rst_BAR, 
                           Q => n14124, QN => n_1295);
   clk_r_REG8191_S9 : DFFR_X1 port map( D => n14124, CK => clk, RN => rst_BAR, 
                           Q => n14123, QN => n_1296);
   clk_r_REG7941_S8 : DFFR_X1 port map( D => n8792, CK => clk, RN => rst_BAR, Q
                           => n14122, QN => n_1297);
   clk_r_REG7656_S5 : DFFR_X1 port map( D => n8791, CK => clk, RN => rst_BAR, Q
                           => n14121, QN => n_1298);
   clk_r_REG7564_S5 : DFFR_X1 port map( D => n8790, CK => clk, RN => rst_BAR, Q
                           => n14120, QN => n_1299);
   clk_r_REG7390_S4 : DFFR_X1 port map( D => n8789, CK => clk, RN => rst_BAR, Q
                           => n14119, QN => n_1300);
   clk_r_REG7320_S4 : DFFR_X1 port map( D => n8788, CK => clk, RN => rst_BAR, Q
                           => n14118, QN => n_1301);
   clk_r_REG7319_S4 : DFFR_X1 port map( D => n8787, CK => clk, RN => rst_BAR, Q
                           => n14117, QN => n_1302);
   clk_r_REG7318_S4 : DFFR_X1 port map( D => n8786, CK => clk, RN => rst_BAR, Q
                           => n14116, QN => n_1303);
   clk_r_REG7316_S4 : DFFR_X1 port map( D => n8785, CK => clk, RN => rst_BAR, Q
                           => n14115, QN => n_1304);
   clk_r_REG7314_S4 : DFFR_X1 port map( D => n8784, CK => clk, RN => rst_BAR, Q
                           => n14114, QN => n_1305);
   clk_r_REG7286_S5 : DFFR_X1 port map( D => n8783, CK => clk, RN => rst_BAR, Q
                           => n14113, QN => n_1306);
   clk_r_REG7271_S5 : DFFR_X1 port map( D => n8782, CK => clk, RN => rst_BAR, Q
                           => n14112, QN => n_1307);
   clk_r_REG7280_S5 : DFFR_X1 port map( D => n8781, CK => clk, RN => rst_BAR, Q
                           => n14111, QN => n_1308);
   clk_r_REG7281_S5 : DFFR_X1 port map( D => n8780, CK => clk, RN => rst_BAR, Q
                           => n14110, QN => n_1309);
   clk_r_REG7282_S5 : DFFR_X1 port map( D => n8779, CK => clk, RN => rst_BAR, Q
                           => n14109, QN => n_1310);
   clk_r_REG7283_S6 : DFFR_X1 port map( D => n14109, CK => clk, RN => rst_BAR, 
                           Q => n14108, QN => n_1311);
   clk_r_REG7727_S5 : DFFR_X1 port map( D => n8773, CK => clk, RN => rst_BAR, Q
                           => n14107, QN => n_1312);
   clk_r_REG7728_S6 : DFFR_X1 port map( D => n14107, CK => clk, RN => rst_BAR, 
                           Q => n14106, QN => n_1313);
   clk_r_REG7729_S7 : DFFR_X1 port map( D => n14106, CK => clk, RN => rst_BAR, 
                           Q => n14105, QN => n_1314);
   clk_r_REG7730_S8 : DFFR_X1 port map( D => n14105, CK => clk, RN => rst_BAR, 
                           Q => n14104, QN => n_1315);
   clk_r_REG7731_S9 : DFFR_X1 port map( D => n14104, CK => clk, RN => rst_BAR, 
                           Q => n14103, QN => n_1316);
   clk_r_REG7277_S6 : DFFR_X1 port map( D => n8772, CK => clk, RN => rst_BAR, Q
                           => n14102, QN => n_1317);
   clk_r_REG7278_S6 : DFFR_X1 port map( D => n8771, CK => clk, RN => rst_BAR, Q
                           => n14101, QN => n_1318);
   clk_r_REG7279_S6 : DFFR_X1 port map( D => n8770, CK => clk, RN => rst_BAR, Q
                           => n14100, QN => n_1319);
   clk_r_REG7540_S5 : DFFR_X1 port map( D => n8765, CK => clk, RN => rst_BAR, Q
                           => n14099, QN => n_1320);
   clk_r_REG7541_S6 : DFFR_X1 port map( D => n14099, CK => clk, RN => rst_BAR, 
                           Q => n14098, QN => n_1321);
   clk_r_REG7542_S7 : DFFR_X1 port map( D => n14098, CK => clk, RN => rst_BAR, 
                           Q => n14097, QN => n_1322);
   clk_r_REG7543_S8 : DFFR_X1 port map( D => n14097, CK => clk, RN => rst_BAR, 
                           Q => n14096, QN => n_1323);
   clk_r_REG7544_S9 : DFFR_X1 port map( D => n14096, CK => clk, RN => rst_BAR, 
                           Q => n14095, QN => n_1324);
   clk_r_REG7275_S6 : DFFR_X1 port map( D => n8763, CK => clk, RN => rst_BAR, Q
                           => n14094, QN => n_1325);
   clk_r_REG7276_S6 : DFFR_X1 port map( D => n8762, CK => clk, RN => rst_BAR, Q
                           => n14093, QN => n_1326);
   clk_r_REG7321_S5 : DFFR_X1 port map( D => n8757, CK => clk, RN => rst_BAR, Q
                           => n14092, QN => n_1327);
   clk_r_REG7322_S6 : DFFR_X1 port map( D => n14092, CK => clk, RN => rst_BAR, 
                           Q => n14091, QN => n_1328);
   clk_r_REG7323_S7 : DFFR_X1 port map( D => n14091, CK => clk, RN => rst_BAR, 
                           Q => n14090, QN => n_1329);
   clk_r_REG7324_S8 : DFFR_X1 port map( D => n14090, CK => clk, RN => rst_BAR, 
                           Q => n14089, QN => n_1330);
   clk_r_REG7325_S9 : DFFR_X1 port map( D => n14089, CK => clk, RN => rst_BAR, 
                           Q => n14088, QN => n_1331);
   clk_r_REG7272_S6 : DFFR_X1 port map( D => n8750, CK => clk, RN => rst_BAR, Q
                           => n14087, QN => n_1332);
   clk_r_REG7273_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CK => clk, RN => rst_BAR, Q => n14086, QN => n_1333)
                           ;
   clk_r_REG7274_S6 : DFFR_X1 port map( D => n3996, CK => clk, RN => rst_BAR, Q
                           => n14085, QN => n_1334);
   clk_r_REG7057_S6 : DFFR_X1 port map( D => n8744, CK => clk, RN => rst_BAR, Q
                           => n14084, QN => n_1335);
   clk_r_REG7058_S7 : DFFR_X1 port map( D => n14084, CK => clk, RN => rst_BAR, 
                           Q => n14083, QN => n_1336);
   clk_r_REG7059_S8 : DFFR_X1 port map( D => n14083, CK => clk, RN => rst_BAR, 
                           Q => n14082, QN => n_1337);
   clk_r_REG7060_S9 : DFFR_X1 port map( D => n14082, CK => clk, RN => rst_BAR, 
                           Q => n14081, QN => n_1338);
   clk_r_REG7061_S10 : DFFR_X1 port map( D => n14081, CK => clk, RN => rst_BAR,
                           Q => n14080, QN => n_1339);
   clk_r_REG7317_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, CK => clk, 
                           RN => rst_BAR, Q => n_1340, QN => n16398);
   clk_r_REG7315_S5 : DFFR_X1 port map( D => n8742, CK => clk, RN => rst_BAR, Q
                           => n14078, QN => n_1341);
   clk_r_REG7287_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CK => clk, RN => rst_BAR, Q => n14077, QN => n_1342)
                           ;
   clk_r_REG7288_S6 : DFFR_X1 port map( D => n8741, CK => clk, RN => rst_BAR, Q
                           => n14076, QN => n_1343);
   clk_r_REG7092_S7 : DFFR_X1 port map( D => n8731, CK => clk, RN => rst_BAR, Q
                           => n14075, QN => n_1344);
   clk_r_REG7072_S7 : DFFR_X1 port map( D => n8730, CK => clk, RN => rst_BAR, Q
                           => n14074, QN => n_1345);
   clk_r_REG7179_S6 : DFFR_X1 port map( D => n8727, CK => clk, RN => rst_BAR, Q
                           => n14073, QN => n_1346);
   clk_r_REG7180_S7 : DFFR_X1 port map( D => n14073, CK => clk, RN => rst_BAR, 
                           Q => n14072, QN => n_1347);
   clk_r_REG7181_S8 : DFFR_X1 port map( D => n14072, CK => clk, RN => rst_BAR, 
                           Q => n14071, QN => n_1348);
   clk_r_REG7182_S9 : DFFR_X1 port map( D => n14071, CK => clk, RN => rst_BAR, 
                           Q => n14070, QN => n_1349);
   clk_r_REG7289_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, CK => clk, 
                           RN => rst_BAR, Q => n_1350, QN => n16397);
   clk_r_REG7230_S6 : DFFR_X1 port map( D => n8725, CK => clk, RN => rst_BAR, Q
                           => n14068, QN => n_1351);
   clk_r_REG7225_S6 : DFFR_X1 port map( D => n8724, CK => clk, RN => rst_BAR, Q
                           => n14067, QN => n_1352);
   clk_r_REG7220_S6 : DFFR_X1 port map( D => n8723, CK => clk, RN => rst_BAR, Q
                           => n14066, QN => n_1353);
   clk_r_REG7216_S6 : DFFR_X1 port map( D => n8722, CK => clk, RN => rst_BAR, Q
                           => n14065, QN => n_1354);
   clk_r_REG7211_S6 : DFFR_X1 port map( D => n8721, CK => clk, RN => rst_BAR, Q
                           => n14064, QN => n_1355);
   clk_r_REG6944_S6 : DFFR_X1 port map( D => n8720, CK => clk, RN => rst_BAR, Q
                           => n14063, QN => n_1356);
   clk_r_REG7207_S6 : DFFR_X1 port map( D => n8719, CK => clk, RN => rst_BAR, Q
                           => n14062, QN => n_1357);
   clk_r_REG7202_S6 : DFFR_X1 port map( D => n8718, CK => clk, RN => rst_BAR, Q
                           => n14061, QN => n_1358);
   clk_r_REG7197_S6 : DFFR_X1 port map( D => n8717, CK => clk, RN => rst_BAR, Q
                           => n14060, QN => n_1359);
   clk_r_REG7098_S7 : DFFR_X1 port map( D => n8716, CK => clk, RN => rst_BAR, Q
                           => n14059, QN => n_1360);
   clk_r_REG7099_S7 : DFFR_X1 port map( D => n8715, CK => clk, RN => rst_BAR, Q
                           => n14058, QN => n_1361);
   clk_r_REG7089_S8 : DFFR_X1 port map( D => n8714, CK => clk, RN => rst_BAR, Q
                           => n14057, QN => n_1362);
   clk_r_REG7090_S8 : DFFR_X1 port map( D => n8713, CK => clk, RN => rst_BAR, Q
                           => n14056, QN => n_1363);
   clk_r_REG7231_S7 : DFFR_X1 port map( D => n8710, CK => clk, RN => rst_BAR, Q
                           => n14055, QN => n_1364);
   clk_r_REG7232_S8 : DFFR_X1 port map( D => n14055, CK => clk, RN => rst_BAR, 
                           Q => n14054, QN => n_1365);
   clk_r_REG7233_S9 : DFFR_X1 port map( D => n14054, CK => clk, RN => rst_BAR, 
                           Q => n14053, QN => n_1366);
   clk_r_REG7226_S7 : DFFR_X1 port map( D => n8708, CK => clk, RN => rst_BAR, Q
                           => n14052, QN => n_1367);
   clk_r_REG7227_S8 : DFFR_X1 port map( D => n14052, CK => clk, RN => rst_BAR, 
                           Q => n14051, QN => n_1368);
   clk_r_REG7228_S9 : DFFR_X1 port map( D => n14051, CK => clk, RN => rst_BAR, 
                           Q => n14050, QN => n_1369);
   clk_r_REG7221_S7 : DFFR_X1 port map( D => n8706, CK => clk, RN => rst_BAR, Q
                           => n14049, QN => n_1370);
   clk_r_REG7222_S8 : DFFR_X1 port map( D => n14049, CK => clk, RN => rst_BAR, 
                           Q => n14048, QN => n_1371);
   clk_r_REG7223_S9 : DFFR_X1 port map( D => n14048, CK => clk, RN => rst_BAR, 
                           Q => n14047, QN => n_1372);
   clk_r_REG7217_S7 : DFFR_X1 port map( D => n8704, CK => clk, RN => rst_BAR, Q
                           => n14046, QN => n_1373);
   clk_r_REG7218_S8 : DFFR_X1 port map( D => n14046, CK => clk, RN => rst_BAR, 
                           Q => n14045, QN => n_1374);
   clk_r_REG7219_S9 : DFFR_X1 port map( D => n14045, CK => clk, RN => rst_BAR, 
                           Q => n14044, QN => n_1375);
   clk_r_REG7212_S7 : DFFR_X1 port map( D => n8702, CK => clk, RN => rst_BAR, Q
                           => n14043, QN => n_1376);
   clk_r_REG7213_S8 : DFFR_X1 port map( D => n14043, CK => clk, RN => rst_BAR, 
                           Q => n14042, QN => n_1377);
   clk_r_REG7214_S9 : DFFR_X1 port map( D => n14042, CK => clk, RN => rst_BAR, 
                           Q => n14041, QN => n_1378);
   clk_r_REG6945_S7 : DFFR_X1 port map( D => n8700, CK => clk, RN => rst_BAR, Q
                           => n14040, QN => n_1379);
   clk_r_REG6946_S8 : DFFR_X1 port map( D => n14040, CK => clk, RN => rst_BAR, 
                           Q => n14039, QN => n_1380);
   clk_r_REG6947_S9 : DFFR_X1 port map( D => n14039, CK => clk, RN => rst_BAR, 
                           Q => n14038, QN => n_1381);
   clk_r_REG7208_S7 : DFFR_X1 port map( D => n8698, CK => clk, RN => rst_BAR, Q
                           => n14037, QN => n_1382);
   clk_r_REG7209_S8 : DFFR_X1 port map( D => n14037, CK => clk, RN => rst_BAR, 
                           Q => n14036, QN => n_1383);
   clk_r_REG7210_S9 : DFFR_X1 port map( D => n14036, CK => clk, RN => rst_BAR, 
                           Q => n14035, QN => n_1384);
   clk_r_REG7203_S7 : DFFR_X1 port map( D => n8696, CK => clk, RN => rst_BAR, Q
                           => n14034, QN => n_1385);
   clk_r_REG7204_S8 : DFFR_X1 port map( D => n14034, CK => clk, RN => rst_BAR, 
                           Q => n14033, QN => n_1386);
   clk_r_REG7205_S9 : DFFR_X1 port map( D => n14033, CK => clk, RN => rst_BAR, 
                           Q => n14032, QN => n_1387);
   clk_r_REG7198_S7 : DFFR_X1 port map( D => n8694, CK => clk, RN => rst_BAR, Q
                           => n14031, QN => n_1388);
   clk_r_REG7199_S8 : DFFR_X1 port map( D => n14031, CK => clk, RN => rst_BAR, 
                           Q => n14030, QN => n_1389);
   clk_r_REG7200_S9 : DFFR_X1 port map( D => n14030, CK => clk, RN => rst_BAR, 
                           Q => n14029, QN => n_1390);
   clk_r_REG7100_S8 : DFFR_X1 port map( D => n8692, CK => clk, RN => rst_BAR, Q
                           => n14028, QN => n_1391);
   clk_r_REG7101_S9 : DFFR_X1 port map( D => n14028, CK => clk, RN => rst_BAR, 
                           Q => n14027, QN => n_1392);
   clk_r_REG7102_S10 : DFFR_X1 port map( D => n14027, CK => clk, RN => rst_BAR,
                           Q => n14026, QN => n_1393);
   clk_r_REG7093_S8 : DFFR_X1 port map( D => n8690, CK => clk, RN => rst_BAR, Q
                           => n14025, QN => n_1394);
   clk_r_REG7094_S9 : DFFR_X1 port map( D => n14025, CK => clk, RN => rst_BAR, 
                           Q => n14024, QN => n_1395);
   clk_r_REG7095_S10 : DFFR_X1 port map( D => n14024, CK => clk, RN => rst_BAR,
                           Q => n14023, QN => n_1396);
   clk_r_REG7073_S8 : DFFR_X1 port map( D => n8689, CK => clk, RN => rst_BAR, Q
                           => n14022, QN => n_1397);
   clk_r_REG7074_S8 : DFFR_X1 port map( D => n8686, CK => clk, RN => rst_BAR, Q
                           => n14021, QN => n_1398);
   clk_r_REG7075_S9 : DFFR_X1 port map( D => n14021, CK => clk, RN => rst_BAR, 
                           Q => n14020, QN => n_1399);
   clk_r_REG7076_S10 : DFFR_X1 port map( D => n14020, CK => clk, RN => rst_BAR,
                           Q => n14019, QN => n_1400);
   clk_r_REG7077_S9 : DFFR_X1 port map( D => n8685, CK => clk, RN => rst_BAR, Q
                           => n14018, QN => n_1401);
   clk_r_REG7078_S10 : DFFR_X1 port map( D => n14018, CK => clk, RN => rst_BAR,
                           Q => n14017, QN => n_1402);
   clk_r_REG7079_S9 : DFFR_X1 port map( D => n8683, CK => clk, RN => rst_BAR, Q
                           => n14016, QN => n_1403);
   clk_r_REG7080_S10 : DFFR_X1 port map( D => n14016, CK => clk, RN => rst_BAR,
                           Q => n14015, QN => n_1404);
   clk_r_REG7081_S9 : DFFR_X1 port map( D => n8682, CK => clk, RN => rst_BAR, Q
                           => n14014, QN => n_1405);
   clk_r_REG7082_S10 : DFFR_X1 port map( D => n14014, CK => clk, RN => rst_BAR,
                           Q => n14013, QN => n_1406);
   clk_r_REG7084_S9 : DFFR_X1 port map( D => n8681, CK => clk, RN => rst_BAR, Q
                           => n14012, QN => n_1407);
   clk_r_REG7085_S10 : DFFR_X1 port map( D => n14012, CK => clk, RN => rst_BAR,
                           Q => n14011, QN => n_1408);
   clk_r_REG7087_S9 : DFFR_X1 port map( D => n8679, CK => clk, RN => rst_BAR, Q
                           => n14010, QN => n_1409);
   clk_r_REG7088_S10 : DFFR_X1 port map( D => n14010, CK => clk, RN => rst_BAR,
                           Q => n14009, QN => n_1410);
   clk_r_REG7252_S3 : DFFR_X1 port map( D => n6095, CK => clk, RN => rst_BAR, Q
                           => n14008, QN => n_1411);
   clk_r_REG7649_S4 : DFFR_X1 port map( D => n11526, CK => clk, RN => rst_BAR, 
                           Q => n14007, QN => n_1412);
   clk_r_REG7042_S4 : DFFR_X1 port map( D => n1880, CK => clk, RN => rst_BAR, Q
                           => n_1413, QN => n14006);
   clk_r_REG7836_S3 : DFFS_X1 port map( D => n1886, CK => clk, SN => rst_BAR, Q
                           => n_1414, QN => n14005);
   clk_r_REG7841_S3 : DFFR_X1 port map( D => n11473, CK => clk, RN => rst_BAR, 
                           Q => n14004, QN => n_1415);
   clk_r_REG7842_S4 : DFFR_X1 port map( D => n11457, CK => clk, RN => rst_BAR, 
                           Q => n14003, QN => n_1416);
   clk_r_REG7839_S3 : DFFR_X1 port map( D => n1883, CK => clk, RN => rst_BAR, Q
                           => n_1417, QN => n14002);
   clk_r_REG7835_S4 : DFFS_X1 port map( D => n11449, CK => clk, SN => rst_BAR, 
                           Q => n14001, QN => n_1418);
   clk_r_REG7814_S3 : DFFS_X1 port map( D => n11436, CK => clk, SN => rst_BAR, 
                           Q => n14000, QN => n_1419);
   clk_r_REG7806_S3 : DFFS_X1 port map( D => n11435, CK => clk, SN => rst_BAR, 
                           Q => n13999, QN => n_1420);
   clk_r_REG7164_S4 : DFFR_X1 port map( D => n1877, CK => clk, RN => rst_BAR, Q
                           => n_1421, QN => n13998);
   clk_r_REG7801_S4 : DFFR_X1 port map( D => n11437, CK => clk, RN => rst_BAR, 
                           Q => n13997, QN => n_1422);
   clk_r_REG7845_S4 : DFFS_X1 port map( D => n1874, CK => clk, SN => rst_BAR, Q
                           => n_1423, QN => n13996);
   clk_r_REG7832_S4 : DFFR_X1 port map( D => n11444, CK => clk, RN => rst_BAR, 
                           Q => n13995, QN => n_1424);
   clk_r_REG7843_S4 : DFFR_X1 port map( D => n1876, CK => clk, RN => rst_BAR, Q
                           => n_1425, QN => n13994);
   clk_r_REG7114_S4 : DFFS_X1 port map( D => n1872, CK => clk, SN => rst_BAR, Q
                           => n18223, QN => n13993);
   clk_r_REG7043_S4 : DFFR_X1 port map( D => n11447, CK => clk, RN => rst_BAR, 
                           Q => n13992, QN => n_1426);
   clk_r_REG7165_S4 : DFFR_X1 port map( D => n11453, CK => clk, RN => rst_BAR, 
                           Q => n13991, QN => n_1427);
   clk_r_REG7817_S3 : DFFS_X1 port map( D => n11459, CK => clk, SN => rst_BAR, 
                           Q => n13990, QN => n_1428);
   clk_r_REG7804_S3 : DFFS_X1 port map( D => n11458, CK => clk, SN => rst_BAR, 
                           Q => n13989, QN => n_1429);
   clk_r_REG7833_S4 : DFFR_X1 port map( D => n11469, CK => clk, RN => rst_BAR, 
                           Q => n13988, QN => n_1430);
   clk_r_REG7520_S4 : DFFR_X1 port map( D => n11485, CK => clk, RN => rst_BAR, 
                           Q => n13987, QN => n_1431);
   clk_r_REG7847_S3 : DFFS_X1 port map( D => n1871, CK => clk, SN => rst_BAR, Q
                           => n_1432, QN => n13986);
   clk_r_REG7849_S3 : DFFS_X1 port map( D => n12392, CK => clk, SN => rst_BAR, 
                           Q => n13985, QN => n_1433);
   clk_r_REG7530_S8 : DFFR_X1 port map( D => n11540, CK => clk, RN => rst_BAR, 
                           Q => n13984, QN => n_1434);
   clk_r_REG7326_S3 : DFFS_X1 port map( D => n8675, CK => clk, SN => rst_BAR, Q
                           => n13983, QN => n_1435);
   clk_r_REG7355_S5 : DFFR_X1 port map( D => n8674, CK => clk, RN => rst_BAR, Q
                           => n13982, QN => n_1436);
   clk_r_REG7354_S5 : DFFR_X1 port map( D => n8673, CK => clk, RN => rst_BAR, Q
                           => n13981, QN => n_1437);
   clk_r_REG7396_S3 : DFFS_X1 port map( D => n8649, CK => clk, SN => rst_BAR, Q
                           => n13980, QN => n_1438);
   clk_r_REG7519_S4 : DFFR_X1 port map( D => n8647, CK => clk, RN => rst_BAR, Q
                           => n13979, QN => n_1439);
   clk_r_REG7405_S5 : DFFS_X1 port map( D => n11729, CK => clk, SN => rst_BAR, 
                           Q => n13978, QN => n_1440);
   clk_r_REG7559_S4 : DFFS_X1 port map( D => n8646, CK => clk, SN => rst_BAR, Q
                           => n13977, QN => n_1441);
   clk_r_REG7545_S3 : DFFS_X1 port map( D => n11754, CK => clk, SN => rst_BAR, 
                           Q => n13976, QN => n_1442);
   clk_r_REG7650_S3 : DFFR_X1 port map( D => n8642, CK => clk, RN => rst_BAR, Q
                           => n13975, QN => n_1443);
   clk_r_REG7531_S9 : DFFS_X1 port map( D => n8640, CK => clk, SN => rst_BAR, Q
                           => n13974, QN => n_1444);
   clk_r_REG7732_S3 : DFFS_X1 port map( D => n8639, CK => clk, SN => rst_BAR, Q
                           => n13973, QN => n_1445);
   clk_r_REG7736_S4 : DFFS_X1 port map( D => n8638, CK => clk, SN => rst_BAR, Q
                           => n13972, QN => n_1446);
   clk_r_REG7434_S4 : DFFS_X1 port map( D => n11789, CK => clk, SN => rst_BAR, 
                           Q => n13971, QN => n_1447);
   clk_r_REG8202_S4 : DFFS_X1 port map( D => n8636, CK => clk, SN => rst_BAR, Q
                           => n13970, QN => n_1448);
   clk_r_REG7749_S3 : DFFS_X1 port map( D => n8635, CK => clk, SN => rst_BAR, Q
                           => n13969, QN => n_1449);
   clk_r_REG8201_S4 : DFFR_X1 port map( D => n8634, CK => clk, RN => rst_BAR, Q
                           => n13968, QN => n_1450);
   clk_r_REG7412_S4 : DFFS_X1 port map( D => n11811, CK => clk, SN => rst_BAR, 
                           Q => n13967, QN => n_1451);
   clk_r_REG7862_S3 : DFFS_X1 port map( D => n8632, CK => clk, SN => rst_BAR, Q
                           => n13966, QN => n_1452);
   clk_r_REG8192_S3 : DFFS_X1 port map( D => n8631, CK => clk, SN => rst_BAR, Q
                           => n13965, QN => n_1453);
   clk_r_REG7414_S4 : DFFR_X1 port map( D => n11849, CK => clk, RN => rst_BAR, 
                           Q => n13964, QN => n_1454);
   clk_r_REG7305_S4 : DFFS_X1 port map( D => n8612, CK => clk, SN => rst_BAR, Q
                           => n13963, QN => n_1455);
   clk_r_REG7435_S4 : DFFR_X1 port map( D => n1855, CK => clk, RN => rst_BAR, Q
                           => n_1456, QN => n13962);
   clk_r_REG7425_S4 : DFFS_X1 port map( D => n1856, CK => clk, SN => rst_BAR, Q
                           => n_1457, QN => n13961);
   clk_r_REG7421_S4 : DFFS_X1 port map( D => n8604, CK => clk, SN => rst_BAR, Q
                           => n13960, QN => n_1458);
   clk_r_REG7040_S4 : DFFS_X1 port map( D => n1875, CK => clk, SN => rst_BAR, Q
                           => n_1459, QN => n13959);
   clk_r_REG7154_S4 : DFFR_X1 port map( D => n1879, CK => clk, RN => rst_BAR, Q
                           => n_1460, QN => n13958);
   clk_r_REG7159_S4 : DFFR_X1 port map( D => n11966, CK => clk, RN => rst_BAR, 
                           Q => n13957, QN => n_1461);
   clk_r_REG7158_S4 : DFFS_X1 port map( D => n11952, CK => clk, SN => rst_BAR, 
                           Q => n13956, QN => n_1462);
   clk_r_REG7157_S4 : DFFS_X1 port map( D => n11955, CK => clk, SN => rst_BAR, 
                           Q => n13955, QN => n_1463);
   clk_r_REG7156_S4 : DFFS_X1 port map( D => n11960, CK => clk, SN => rst_BAR, 
                           Q => n13954, QN => n_1464);
   clk_r_REG7039_S4 : DFFS_X1 port map( D => n11959, CK => clk, SN => rst_BAR, 
                           Q => n13953, QN => n_1465);
   clk_r_REG7304_S4 : DFFR_X1 port map( D => n11979, CK => clk, RN => rst_BAR, 
                           Q => n13952, QN => n_1466);
   clk_r_REG7302_S4 : DFFR_X1 port map( D => n1885, CK => clk, RN => rst_BAR, Q
                           => n_1467, QN => n13951);
   clk_r_REG7301_S4 : DFFR_X1 port map( D => n11981, CK => clk, RN => rst_BAR, 
                           Q => n13950, QN => n_1468);
   clk_r_REG7036_S4 : DFFS_X1 port map( D => n11996, CK => clk, SN => rst_BAR, 
                           Q => n13949, QN => n_1469);
   clk_r_REG7035_S4 : DFFS_X1 port map( D => n12004, CK => clk, SN => rst_BAR, 
                           Q => n13948, QN => n_1470);
   clk_r_REG7430_S4 : DFFS_X1 port map( D => n12032, CK => clk, SN => rst_BAR, 
                           Q => n13947, QN => n_1471);
   clk_r_REG7306_S4 : DFFR_X1 port map( D => n12031, CK => clk, RN => rst_BAR, 
                           Q => n13946, QN => n_1472);
   clk_r_REG7429_S4 : DFFR_X1 port map( D => n12042, CK => clk, RN => rst_BAR, 
                           Q => n13945, QN => n_1473);
   clk_r_REG7423_S4 : DFFR_X1 port map( D => n12045, CK => clk, RN => rst_BAR, 
                           Q => n13944, QN => n_1474);
   clk_r_REG7415_S4 : DFFR_X1 port map( D => n12047, CK => clk, RN => rst_BAR, 
                           Q => n13943, QN => n_1475);
   clk_r_REG7014_S4 : DFFR_X1 port map( D => n12088, CK => clk, RN => rst_BAR, 
                           Q => n13942, QN => n_1476);
   clk_r_REG7037_S4 : DFFR_X1 port map( D => n12087, CK => clk, RN => rst_BAR, 
                           Q => n13941, QN => n_1477);
   clk_r_REG7034_S4 : DFFS_X1 port map( D => n12086, CK => clk, SN => rst_BAR, 
                           Q => n13940, QN => n_1478);
   clk_r_REG7417_S4 : DFFS_X1 port map( D => n12526, CK => clk, SN => rst_BAR, 
                           Q => n13939, QN => n_1479);
   clk_r_REG7086_S11 : DFFR_X1 port map( D => n8601, CK => clk, RN => rst_BAR, 
                           Q => n13938, QN => n_1480);
   clk_r_REG6993_S5 : DFFS_X1 port map( D => n12162, CK => clk, SN => rst_BAR, 
                           Q => n13937, QN => n_1481);
   clk_r_REG7863_S3 : DFFS_X1 port map( D => n8600, CK => clk, SN => rst_BAR, Q
                           => n13936, QN => n_1482);
   clk_r_REG8199_S3 : DFFS_X1 port map( D => n8599, CK => clk, SN => rst_BAR, Q
                           => n13935, QN => n_1483);
   clk_r_REG7410_S4 : DFFS_X1 port map( D => n1861, CK => clk, SN => rst_BAR, Q
                           => n_1484, QN => n13934);
   clk_r_REG7413_S4 : DFFR_X1 port map( D => n12189, CK => clk, RN => rst_BAR, 
                           Q => n13933, QN => n_1485);
   clk_r_REG7083_S11 : DFFS_X1 port map( D => n8596, CK => clk, SN => rst_BAR, 
                           Q => n13932, QN => n_1486);
   clk_r_REG7740_S4 : DFFS_X1 port map( D => n8595, CK => clk, SN => rst_BAR, Q
                           => n13931, QN => n_1487);
   clk_r_REG6984_S4 : DFFR_X1 port map( D => n12213, CK => clk, RN => rst_BAR, 
                           Q => n13930, QN => n_1488);
   clk_r_REG6977_S5 : DFFS_X1 port map( D => n12229, CK => clk, SN => rst_BAR, 
                           Q => n13929, QN => n_1489);
   clk_r_REG6970_S4 : DFFS_X1 port map( D => n12246, CK => clk, SN => rst_BAR, 
                           Q => n13928, QN => n_1490);
   clk_r_REG6963_S5 : DFFS_X1 port map( D => n12254, CK => clk, SN => rst_BAR, 
                           Q => n13927, QN => n_1491);
   clk_r_REG6955_S4 : DFFR_X1 port map( D => n8591, CK => clk, RN => rst_BAR, Q
                           => n13926, QN => n_1492);
   clk_r_REG7103_S11 : DFFS_X1 port map( D => n12273, CK => clk, SN => rst_BAR,
                           Q => n13925, QN => n_1493);
   clk_r_REG7206_S10 : DFFS_X1 port map( D => n8588, CK => clk, SN => rst_BAR, 
                           Q => n13924, QN => n_1494);
   clk_r_REG7143_S4 : DFFR_X1 port map( D => n8584, CK => clk, RN => rst_BAR, Q
                           => n13923, QN => n_1495);
   clk_r_REG8344_S3 : DFFS_X1 port map( D => n8581, CK => clk, SN => rst_BAR, Q
                           => n13922, QN => n_1496);
   clk_r_REG7409_S4 : DFFS_X1 port map( D => n12722, CK => clk, SN => rst_BAR, 
                           Q => n13921, QN => n_1497);
   clk_r_REG7215_S10 : DFFS_X1 port map( D => n8579, CK => clk, SN => rst_BAR, 
                           Q => n13920, QN => n_1498);
   clk_r_REG7136_S4 : DFFR_X1 port map( D => n8578, CK => clk, RN => rst_BAR, Q
                           => n13919, QN => n_1499);
   clk_r_REG7224_S10 : DFFS_X1 port map( D => n8574, CK => clk, SN => rst_BAR, 
                           Q => n13918, QN => n_1500);
   clk_r_REG7122_S4 : DFFR_X1 port map( D => n8573, CK => clk, RN => rst_BAR, Q
                           => n13917, QN => n_1501);
   clk_r_REG7248_S4 : DFFR_X1 port map( D => n8572, CK => clk, RN => rst_BAR, Q
                           => n13916, QN => n_1502);
   clk_r_REG7229_S10 : DFFS_X1 port map( D => n8571, CK => clk, SN => rst_BAR, 
                           Q => n13915, QN => n_1503);
   clk_r_REG7234_S10 : DFFS_X1 port map( D => n12446, CK => clk, SN => rst_BAR,
                           Q => n13914, QN => n_1504);
   clk_r_REG7253_S3 : DFFR_X1 port map( D => n8942, CK => clk, RN => rst_BAR, Q
                           => n13913, QN => n_1505);
   clk_r_REG7360_S5 : DFFS_X1 port map( D => n8823, CK => clk, SN => rst_BAR, Q
                           => n13912, QN => n_1506);
   clk_r_REG7420_S4 : DFFR_X1 port map( D => n12473, CK => clk, RN => rst_BAR, 
                           Q => n13911, QN => n_1507);
   clk_r_REG7062_S11 : DFFS_X1 port map( D => n8567, CK => clk, SN => rst_BAR, 
                           Q => n13910, QN => n_1508);
   clk_r_REG7358_S5 : DFFS_X1 port map( D => n12509, CK => clk, SN => rst_BAR, 
                           Q => n13909, QN => n_1509);
   clk_r_REG6920_S10 : DFFS_X1 port map( D => n8565, CK => clk, SN => rst_BAR, 
                           Q => n13908, QN => n_1510);
   clk_r_REG7010_S4 : DFFR_X1 port map( D => n12751, CK => clk, RN => rst_BAR, 
                           Q => n13907, QN => n_1511);
   clk_r_REG7009_S4 : DFFS_X1 port map( D => n12750, CK => clk, SN => rst_BAR, 
                           Q => n13906, QN => n_1512);
   clk_r_REG7408_S4 : DFFS_X1 port map( D => n12721, CK => clk, SN => rst_BAR, 
                           Q => n13905, QN => n_1513);
   clk_r_REG7336_S6 : DFFR_X1 port map( D => n8927, CK => clk, RN => rst_BAR, Q
                           => n13904, QN => n_1514);
   clk_r_REG7337_S6 : DFFR_X1 port map( D => n8926, CK => clk, RN => rst_BAR, Q
                           => n13903, QN => n_1515);
   clk_r_REG7338_S6 : DFFR_X1 port map( D => n8925, CK => clk, RN => rst_BAR, Q
                           => n13902, QN => n_1516);
   clk_r_REG7339_S6 : DFFR_X1 port map( D => n8924, CK => clk, RN => rst_BAR, Q
                           => n13901, QN => n_1517);
   clk_r_REG7340_S6 : DFFR_X1 port map( D => n8923, CK => clk, RN => rst_BAR, Q
                           => n13900, QN => n_1518);
   clk_r_REG7285_S5 : DFFR_X1 port map( D => n8922, CK => clk, RN => rst_BAR, Q
                           => n13899, QN => n_1519);
   clk_r_REG7284_S5 : DFFR_X1 port map( D => n8921, CK => clk, RN => rst_BAR, Q
                           => n13898, QN => n_1520);
   clk_r_REG7091_S6 : DFFR_X1 port map( D => n8918, CK => clk, RN => rst_BAR, Q
                           => n13897, QN => n_1521);
   clk_r_REG7194_S6 : DFFR_X1 port map( D => n8915, CK => clk, RN => rst_BAR, Q
                           => n13896, QN => n_1522);
   clk_r_REG7766_S3 : DFFR_X1 port map( D => n16401, CK => clk, RN => rst_BAR, 
                           Q => n18221, QN => n13895);
   clk_r_REG7765_S3 : DFFS_X1 port map( D => n16401, CK => clk, SN => rst_BAR, 
                           Q => n_1523, QN => n13894);
   clk_r_REG7760_S3 : DFFS_X1 port map( D => n16400, CK => clk, SN => rst_BAR, 
                           Q => n18182, QN => n13893);
   clk_r_REG7411_S4 : DFFR_X1 port map( D => n1862, CK => clk, RN => rst_BAR, Q
                           => n_1524, QN => n13892);
   clk_r_REG7428_S4 : DFFS_X1 port map( D => n1852, CK => clk, SN => rst_BAR, Q
                           => n_1525, QN => n13891);
   clk_r_REG7382_S4 : DFFS_X1 port map( D => n1863, CK => clk, SN => rst_BAR, Q
                           => n_1526, QN => n13890);
   clk_r_REG7300_S4 : DFFS_X1 port map( D => n13186, CK => clk, SN => rst_BAR, 
                           Q => n18188, QN => n16399);
   clk_r_REG8020_S11 : DFFR_X1 port map( D => n8555, CK => clk, RN => rst_BAR, 
                           Q => n13888, QN => n_1527);
   clk_r_REG8021_S12 : DFFR_X1 port map( D => n13888, CK => clk, RN => rst_BAR,
                           Q => n13887, QN => n_1528);
   clk_r_REG8022_S13 : DFFR_X1 port map( D => n13887, CK => clk, RN => rst_BAR,
                           Q => n13886, QN => n_1529);
   clk_r_REG8023_S14 : DFFR_X1 port map( D => n13886, CK => clk, RN => rst_BAR,
                           Q => n13885, QN => n_1530);
   clk_r_REG8024_S15 : DFFR_X1 port map( D => n13885, CK => clk, RN => rst_BAR,
                           Q => n13884, QN => n_1531);
   clk_r_REG7635_S5 : DFFR_X1 port map( D => n8880, CK => clk, RN => rst_BAR, Q
                           => n13883, QN => n_1532);
   clk_r_REG7636_S6 : DFFR_X1 port map( D => n13883, CK => clk, RN => rst_BAR, 
                           Q => n13882, QN => n_1533);
   clk_r_REG7637_S7 : DFFR_X1 port map( D => n13882, CK => clk, RN => rst_BAR, 
                           Q => n13881, QN => n_1534);
   clk_r_REG7638_S8 : DFFR_X1 port map( D => n13881, CK => clk, RN => rst_BAR, 
                           Q => n13880, QN => n_1535);
   clk_r_REG7639_S9 : DFFR_X1 port map( D => n13880, CK => clk, RN => rst_BAR, 
                           Q => n13879, QN => n_1536);
   clk_r_REG7640_S10 : DFFS_X1 port map( D => n13879, CK => clk, SN => rst_BAR,
                           Q => n13878, QN => n_1537);
   clk_r_REG7051_S6 : DFFR_X1 port map( D => n8871, CK => clk, RN => rst_BAR, Q
                           => n13877, QN => n_1538);
   clk_r_REG7052_S7 : DFFR_X1 port map( D => n13877, CK => clk, RN => rst_BAR, 
                           Q => n13876, QN => n_1539);
   clk_r_REG7053_S8 : DFFR_X1 port map( D => n13876, CK => clk, RN => rst_BAR, 
                           Q => n13875, QN => n_1540);
   clk_r_REG7054_S9 : DFFR_X1 port map( D => n13875, CK => clk, RN => rst_BAR, 
                           Q => n13874, QN => n_1541);
   clk_r_REG7055_S10 : DFFR_X1 port map( D => n13874, CK => clk, RN => rst_BAR,
                           Q => n13873, QN => n_1542);
   clk_r_REG7174_S6 : DFFR_X1 port map( D => n8867, CK => clk, RN => rst_BAR, Q
                           => n13872, QN => n_1543);
   clk_r_REG7175_S7 : DFFR_X1 port map( D => n13872, CK => clk, RN => rst_BAR, 
                           Q => n13871, QN => n_1544);
   clk_r_REG7176_S8 : DFFR_X1 port map( D => n13871, CK => clk, RN => rst_BAR, 
                           Q => n13870, QN => n_1545);
   clk_r_REG7177_S9 : DFFR_X1 port map( D => n13870, CK => clk, RN => rst_BAR, 
                           Q => n13869, QN => n_1546);
   clk_r_REG7178_S10 : DFFS_X1 port map( D => n13869, CK => clk, SN => rst_BAR,
                           Q => n13868, QN => n_1547);
   clk_r_REG8345_S4 : DFFS_X1 port map( D => n8553, CK => clk, SN => rst_BAR, Q
                           => n13867, QN => n_1548);
   clk_r_REG7263_S7 : DFFR_X1 port map( D => n8824, CK => clk, RN => rst_BAR, Q
                           => n13866, QN => n_1549);
   clk_r_REG7264_S8 : DFFR_X1 port map( D => n13866, CK => clk, RN => rst_BAR, 
                           Q => n13865, QN => n_1550);
   clk_r_REG7265_S9 : DFFR_X1 port map( D => n13865, CK => clk, RN => rst_BAR, 
                           Q => n13864, QN => n_1551);
   clk_r_REG7364_S5 : DFFS_X1 port map( D => n8551, CK => clk, SN => rst_BAR, Q
                           => n13863, QN => n_1552);
   clk_r_REG7363_S5 : DFFR_X1 port map( D => n8550, CK => clk, RN => rst_BAR, Q
                           => n13862, QN => n_1553);
   clk_r_REG7294_S5 : DFFR_X1 port map( D => n8549, CK => clk, RN => rst_BAR, Q
                           => n13861, QN => n_1554);
   clk_r_REG7071_S6 : DFFR_X1 port map( D => n8548, CK => clk, RN => rst_BAR, Q
                           => n13860, QN => n_1555);
   clk_r_REG7193_S6 : DFFR_X1 port map( D => n8547, CK => clk, RN => rst_BAR, Q
                           => n13859, QN => n_1556);
   clk_r_REG7419_S4 : DFFR_X1 port map( D => n12487, CK => clk, RN => rst_BAR, 
                           Q => n13858, QN => n_1557);
   clk_r_REG7362_S5 : DFFR_X1 port map( D => n8819, CK => clk, RN => rst_BAR, Q
                           => n13857, QN => n_1558);
   clk_r_REG7864_S3 : DFFS_X1 port map( D => n8818, CK => clk, SN => rst_BAR, Q
                           => n13856, QN => n_1559);
   clk_r_REG6943_S5 : DFFR_X1 port map( D => n8535, CK => clk, RN => rst_BAR, Q
                           => n13855, QN => n_1560);
   clk_r_REG7295_S5 : DFFR_X1 port map( D => n8534, CK => clk, RN => rst_BAR, Q
                           => n13854, QN => n_1561);
   clk_r_REG8338_S4 : DFFR_X1 port map( D => n8528, CK => clk, RN => rst_BAR, Q
                           => n13853, QN => n_1562);
   clk_r_REG8339_S5 : DFFR_X1 port map( D => n13853, CK => clk, RN => rst_BAR, 
                           Q => n13852, QN => n_1563);
   clk_r_REG8340_S6 : DFFR_X1 port map( D => n13852, CK => clk, RN => rst_BAR, 
                           Q => n13851, QN => n_1564);
   clk_r_REG8341_S7 : DFFR_X1 port map( D => n13851, CK => clk, RN => rst_BAR, 
                           Q => n13850, QN => n_1565);
   clk_r_REG8342_S8 : DFFR_X1 port map( D => n13850, CK => clk, RN => rst_BAR, 
                           Q => n13849, QN => n_1566);
   clk_r_REG8343_S9 : DFFR_X1 port map( D => n13849, CK => clk, RN => rst_BAR, 
                           Q => n13848, QN => n_1567);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n554, Q => 
                           DATA2_I_28_port);
   clk_r_REG7851_S3 : DFFR_X1 port map( D => n1897, CK => clk, RN => rst_BAR, Q
                           => n18187, QN => n14231);
   clk_r_REG7826_S3 : DFFR_X1 port map( D => n16404, CK => clk, RN => rst_BAR, 
                           Q => n18181, QN => n14134);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port);
   clk_r_REG7341_S5 : DFFS_X1 port map( D => n12927, CK => clk, SN => rst_BAR, 
                           Q => n14141, QN => n_1568);
   clk_r_REG7344_S5 : DFFR_X1 port map( D => n12924, CK => clk, RN => rst_BAR, 
                           Q => n14285, QN => n_1569);
   clk_r_REG7342_S5 : DFFS_X1 port map( D => n16416, CK => clk, SN => rst_BAR, 
                           Q => n_1570, QN => n14284);
   clk_r_REG7557_S5 : DFFR_X1 port map( D => n1847, CK => clk, RN => rst_BAR, Q
                           => n_1571, QN => n14283);
   clk_r_REG7553_S5 : DFFR_X1 port map( D => n16419, CK => clk, RN => rst_BAR, 
                           Q => n14419, QN => n_1572);
   clk_r_REG7794_S3 : DFFR_X1 port map( D => n16408, CK => clk, RN => rst_BAR, 
                           Q => n_1573, QN => n14228);
   clk_r_REG6941_S4 : DFFS_X1 port map( D => n16417, CK => clk, SN => rst_BAR, 
                           Q => n_1574, QN => n14223);
   clk_r_REG7554_S5 : DFFS_X1 port map( D => n8931, CK => clk, SN => rst_BAR, Q
                           => n14251, QN => n_1575);
   U3 : NOR2_X2 port map( A1 => n14290, A2 => n17970, ZN => n17999);
   U4 : NOR2_X2 port map( A1 => n16389, A2 => n18008, ZN => n18042);
   U5 : NOR2_X2 port map( A1 => n18199, A2 => n18008, ZN => n18041);
   U6 : INV_X2 port map( A => n17192, ZN => n17279);
   U7 : AOI21_X2 port map( B1 => n18060, B2 => DATA2(3), A => n16653, ZN => 
                           n1897);
   U8 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_2_3_port,
                           A2 => n17802, ZN => n17833);
   U9 : NOR2_X2 port map( A1 => n17970, A2 => n16390, ZN => n18003);
   U10 : NOR2_X2 port map( A1 => n14287, A2 => n17932, ZN => n17965);
   U11 : NOR3_X4 port map( A1 => n16389, A2 => n14292, A3 => n16394, ZN => 
                           n18043);
   U12 : NOR2_X2 port map( A1 => n16978, A2 => n18069, ZN => n17339);
   U13 : INV_X1 port map( A => n18150, ZN => n18116);
   U14 : INV_X2 port map( A => n18137, ZN => n18159);
   U15 : INV_X1 port map( A => n18152, ZN => n18144);
   U16 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n16440);
   U17 : INV_X1 port map( A => n554, ZN => n17769);
   U18 : INV_X1 port map( A => n9078, ZN => n1839);
   U19 : INV_X1 port map( A => data1_mul_0_port, ZN => n1844);
   U20 : INV_X1 port map( A => n7769, ZN => n18075);
   U21 : NAND3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4295, A3 => n18075, ZN => n8814);
   U22 : NOR2_X1 port map( A1 => n7769, A2 => n8978, ZN => n18072);
   U23 : AOI21_X1 port map( B1 => n8978, B2 => n7769, A => n18072, ZN => n1846)
                           ;
   U24 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_2_4_port, ZN => 
                           n1835);
   U25 : NOR2_X1 port map( A1 => n4295, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n17871);
   U26 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, B2 
                           => n4295, A => n17871, ZN => n1848);
   U27 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n17841);
   U28 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n17841, ZN => n8900);
   U29 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_5_port, 
                           ZN => n18073);
   U30 : OR2_X1 port map( A1 => n18073, A2 => n8900, ZN => n16417);
   U31 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n1821);
   U32 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n1819);
   U33 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n1817);
   U34 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n1815);
   U35 : INV_X1 port map( A => data1_mul_15_port, ZN => n1814);
   U36 : XOR2_X1 port map( A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, B 
                           => n1814, Z => n18051);
   U37 : INV_X1 port map( A => n18051, ZN => n1812);
   U38 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n1813);
   U39 : NAND2_X1 port map( A1 => DATA2(4), A2 => DATA2(3), ZN => n18077);
   U40 : INV_X1 port map( A => DATA2(1), ZN => n18059);
   U41 : NAND2_X1 port map( A1 => n18059, A2 => DATA2(0), ZN => n18069);
   U42 : OR3_X1 port map( A1 => n18077, A2 => n18069, A3 => DATA2(2), ZN => 
                           n16402);
   U43 : NOR2_X2 port map( A1 => DATA2(5), A2 => DATA2(4), ZN => n13099);
   U44 : INV_X1 port map( A => DATA2(3), ZN => n18082);
   U45 : NOR2_X1 port map( A1 => n13099, A2 => n18082, ZN => n13096);
   U46 : INV_X1 port map( A => DATA2(0), ZN => n18062);
   U47 : NOR2_X1 port map( A1 => n18059, A2 => n18062, ZN => n18060);
   U48 : INV_X1 port map( A => n18060, ZN => n18078);
   U49 : NOR2_X1 port map( A1 => n18078, A2 => DATA2(2), ZN => n18063);
   U50 : AND3_X1 port map( A1 => n18082, A2 => DATA2(4), A3 => n18063, ZN => 
                           n16412);
   U51 : NOR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n18081);
   U52 : INV_X1 port map( A => n18081, ZN => n18066);
   U53 : NOR2_X1 port map( A1 => n18066, A2 => DATA2(2), ZN => n18083);
   U54 : OR2_X1 port map( A1 => n18077, A2 => n18083, ZN => n1904);
   U55 : INV_X1 port map( A => DATA2(2), ZN => n18079);
   U56 : OAI21_X1 port map( B1 => n18082, B2 => n18079, A => n13099, ZN => 
                           n16653);
   U57 : INV_X1 port map( A => n16653, ZN => n16652);
   U58 : AOI21_X1 port map( B1 => n13099, B2 => n18078, A => n16652, ZN => 
                           n1899);
   U59 : INV_X1 port map( A => n1899, ZN => n9011);
   U60 : INV_X1 port map( A => FUNC(2), ZN => n16436);
   U61 : NAND2_X1 port map( A1 => n16440, A2 => n16436, ZN => n554);
   U62 : INV_X1 port map( A => n17769, ZN => n18230);
   U63 : NAND2_X1 port map( A1 => n14464, A2 => DATA2_I_4_port, ZN => n16727);
   U64 : OAI21_X1 port map( B1 => n14464, B2 => DATA2_I_4_port, A => n16727, ZN
                           => n1429);
   U65 : INV_X1 port map( A => DATA1(21), ZN => n16606);
   U66 : XNOR2_X1 port map( A => DATA2_I_21_port, B => n16606, ZN => n1809);
   U67 : INV_X1 port map( A => FUNC(3), ZN => n1870);
   U68 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n16435);
   U69 : INV_X1 port map( A => DATA1(20), ZN => n16566);
   U70 : XOR2_X1 port map( A => DATA2_I_20_port, B => n16566, Z => n16452);
   U71 : INV_X1 port map( A => n16452, ZN => n17326);
   U72 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => n16434
                           );
   U73 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n17393);
   U74 : XOR2_X1 port map( A => DATA1(17), B => DATA2_I_17_port, Z => n17408);
   U75 : NAND3_X1 port map( A1 => DATA1(16), A2 => n17408, A3 => 
                           DATA2_I_16_port, ZN => n17412);
   U76 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n16433);
   U77 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => n16433
                           , ZN => n17392);
   U78 : AOI21_X1 port map( B1 => n17393, B2 => n17412, A => n17392, ZN => 
                           n17394);
   U79 : AOI21_X1 port map( B1 => DATA2_I_18_port, B2 => DATA1(18), A => n17394
                           , ZN => n17380);
   U80 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n16451);
   U81 : OAI21_X1 port map( B1 => n16434, B2 => n17380, A => n16451, ZN => 
                           n17323);
   U82 : NAND2_X1 port map( A1 => n17326, A2 => n17323, ZN => n17322);
   U83 : NAND2_X1 port map( A1 => n16435, A2 => n17322, ZN => n18172);
   U84 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n16430);
   U85 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => n16430
                           , ZN => n17444);
   U86 : INV_X1 port map( A => DATA1(14), ZN => n17655);
   U87 : XOR2_X1 port map( A => DATA2_I_14_port, B => n17655, Z => n17459);
   U88 : INV_X1 port map( A => n17459, ZN => n17467);
   U89 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n17456);
   U90 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => n17456
                           , ZN => n17476);
   U91 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n17475);
   U92 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => n17475
                           , ZN => n18165);
   U93 : NOR2_X1 port map( A1 => n17476, A2 => n18165, ZN => n17438);
   U94 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => n16421
                           );
   U95 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n17512)
                           ;
   U96 : XNOR2_X1 port map( A => DATA1(9), B => DATA2_I_9_port, ZN => n16761);
   U97 : INV_X1 port map( A => n16761, ZN => n16420);
   U98 : NAND3_X1 port map( A1 => n14469, A2 => n16420, A3 => DATA2_I_8_port, 
                           ZN => n17523);
   U99 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n17435);
   U100 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n17435, ZN => n17513);
   U101 : AOI21_X1 port map( B1 => n17512, B2 => n17523, A => n17513, ZN => 
                           n17509);
   U102 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => DATA1(10), A => 
                           n17509, ZN => n17496);
   U103 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n17436);
   U104 : OAI21_X1 port map( B1 => n16421, B2 => n17496, A => n17436, ZN => 
                           n17483);
   U105 : NOR2_X1 port map( A1 => n17476, A2 => n17475, ZN => n17437);
   U106 : AOI21_X1 port map( B1 => n17438, B2 => n17483, A => n17437, ZN => 
                           n17458);
   U107 : NAND2_X1 port map( A1 => n17458, A2 => n17456, ZN => n17462);
   U108 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n17467, B2 => n17462, ZN => n17445);
   U109 : NOR2_X1 port map( A1 => n14469, A2 => DATA2_I_8_port, ZN => n16758);
   U110 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => n14469, A => n16758, 
                           ZN => n16806);
   U111 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n17436, ZN => n17501);
   U112 : NOR4_X1 port map( A1 => n17513, A2 => n16761, A3 => n17459, A4 => 
                           n17501, ZN => n16429);
   U113 : NAND2_X1 port map( A1 => DATA2_I_7_port, A2 => n14467, ZN => n16427);
   U114 : OAI21_X1 port map( B1 => DATA2_I_7_port, B2 => n14467, A => n16427, 
                           ZN => n16818);
   U115 : NAND2_X1 port map( A1 => n14466, A2 => DATA2_I_6_port, ZN => n16819);
   U116 : XOR2_X1 port map( A => n14326, B => DATA2_I_3_port, Z => n16723);
   U117 : NAND2_X1 port map( A1 => n14327, A2 => DATA2_I_2_port, ZN => n16721);
   U118 : OAI21_X1 port map( B1 => n14327, B2 => DATA2_I_2_port, A => n16721, 
                           ZN => n17150);
   U119 : NAND2_X1 port map( A1 => n14463, A2 => DATA2_I_1_port, ZN => n16724);
   U120 : NAND2_X1 port map( A1 => n14461, A2 => DATA2_I_0_port, ZN => n17341);
   U121 : INV_X1 port map( A => n17341, ZN => n17532);
   U122 : NOR2_X1 port map( A1 => n14461, A2 => DATA2_I_0_port, ZN => n17531);
   U123 : OAI21_X1 port map( B1 => n14463, B2 => DATA2_I_1_port, A => n16724, 
                           ZN => n17340);
   U124 : NOR2_X1 port map( A1 => n17531, A2 => n17340, ZN => n17336);
   U125 : OAI21_X1 port map( B1 => n14460, B2 => n17532, A => n17336, ZN => 
                           n16422);
   U126 : OAI221_X1 port map( B1 => n17150, B2 => n16724, C1 => n17150, C2 => 
                           n16422, A => n16721, ZN => n16423);
   U127 : AND2_X1 port map( A1 => n14326, A2 => DATA2_I_3_port, ZN => n16726);
   U128 : AOI21_X1 port map( B1 => n16723, B2 => n16423, A => n16726, ZN => 
                           n16424);
   U129 : XOR2_X1 port map( A => n14453, B => DATA2_I_5_port, Z => n16855);
   U130 : AOI221_X1 port map( B1 => n16424, B2 => n16727, C1 => n1429, C2 => 
                           n16727, A => n16855, ZN => n16426);
   U131 : AND2_X1 port map( A1 => n14465, A2 => DATA2_I_5_port, ZN => n16728);
   U132 : XNOR2_X1 port map( A => DATA2_I_6_port, B => n14466, ZN => n16845);
   U133 : INV_X1 port map( A => n16845, ZN => n16425);
   U134 : OAI21_X1 port map( B1 => n16426, B2 => n16728, A => n16425, ZN => 
                           n16428);
   U135 : OAI221_X1 port map( B1 => n16818, B2 => n16819, C1 => n16818, C2 => 
                           n16428, A => n16427, ZN => n17473);
   U136 : NAND4_X1 port map( A1 => n17438, A2 => n16806, A3 => n16429, A4 => 
                           n17473, ZN => n16431);
   U137 : OAI221_X1 port map( B1 => n17444, B2 => n17445, C1 => n17444, C2 => 
                           n16431, A => n16430, ZN => n16453);
   U138 : NOR2_X1 port map( A1 => n18230, A2 => n16453, ZN => n18173);
   U139 : INV_X1 port map( A => n18173, ZN => n17413);
   U140 : NAND2_X1 port map( A1 => n17769, A2 => n16453, ZN => n17409);
   U141 : OAI21_X1 port map( B1 => DATA1(16), B2 => DATA2_I_16_port, A => 
                           n17408, ZN => n17396);
   U142 : AOI21_X1 port map( B1 => n17393, B2 => n17396, A => n17392, ZN => 
                           n16432);
   U143 : INV_X1 port map( A => n16432, ZN => n17397);
   U144 : AND2_X1 port map( A1 => n16433, A2 => n17397, ZN => n17382);
   U145 : OAI21_X1 port map( B1 => n16434, B2 => n17382, A => n16451, ZN => 
                           n17325);
   U146 : NAND2_X1 port map( A1 => n17326, A2 => n17325, ZN => n17324);
   U147 : NAND2_X1 port map( A1 => n16435, A2 => n17324, ZN => n18174);
   U148 : OAI22_X1 port map( A1 => n18172, A2 => n17413, B1 => n17409, B2 => 
                           n18174, ZN => n16438);
   U149 : NAND3_X1 port map( A1 => FUNC(2), A2 => FUNC(3), A3 => n16440, ZN => 
                           n17530);
   U150 : INV_X1 port map( A => DATA2(21), ZN => n17780);
   U151 : INV_X1 port map( A => FUNC(0), ZN => n17572);
   U152 : NAND3_X1 port map( A1 => n16436, A2 => n17572, A3 => FUNC(1), ZN => 
                           n17521);
   U153 : INV_X1 port map( A => n17521, ZN => n18171);
   U154 : NAND2_X1 port map( A1 => n18171, A2 => n1870, ZN => n17424);
   U155 : OAI21_X1 port map( B1 => n17530, B2 => n17780, A => n17424, ZN => 
                           n16437);
   U156 : AOI22_X1 port map( A1 => n16438, A2 => n1809, B1 => n16437, B2 => 
                           DATA1(21), ZN => n16439);
   U157 : INV_X1 port map( A => n16439, ZN => n8584);
   U158 : NAND3_X1 port map( A1 => FUNC(2), A2 => n16440, A3 => n1870, ZN => 
                           n7822);
   U159 : NOR4_X1 port map( A1 => DATA2(12), A2 => DATA2(8), A3 => DATA2(7), A4
                           => DATA2(15), ZN => n16447);
   U160 : NAND2_X1 port map( A1 => n13099, A2 => n18082, ZN => n16488);
   U161 : OR2_X1 port map( A1 => DATA2(2), A2 => n16488, ZN => n16978);
   U162 : INV_X1 port map( A => n16978, ZN => n17264);
   U163 : NAND2_X1 port map( A1 => n18081, A2 => n17264, ZN => n17000);
   U164 : INV_X1 port map( A => DATA2(14), ZN => n17787);
   U165 : INV_X1 port map( A => DATA2(13), ZN => n17788);
   U166 : INV_X1 port map( A => DATA2(10), ZN => n17790);
   U167 : INV_X1 port map( A => DATA2(9), ZN => n17791);
   U168 : NAND4_X1 port map( A1 => n17787, A2 => n17788, A3 => n17790, A4 => 
                           n17791, ZN => n16441);
   U169 : NOR4_X1 port map( A1 => DATA2(11), A2 => DATA2(6), A3 => n17000, A4 
                           => n16441, ZN => n16446);
   U170 : INV_X1 port map( A => DATA1(13), ZN => n16493);
   U171 : INV_X1 port map( A => DATA1(12), ZN => n18161);
   U172 : INV_X1 port map( A => DATA1(9), ZN => n16514);
   U173 : NAND4_X1 port map( A1 => n17655, A2 => n16493, A3 => n18161, A4 => 
                           n16514, ZN => n16444);
   U174 : NOR4_X1 port map( A1 => DATA1(11), A2 => n14469, A3 => n14327, A4 => 
                           n14467, ZN => n16442);
   U175 : INV_X1 port map( A => DATA1(10), ZN => n17520);
   U176 : INV_X1 port map( A => DATA1(15), ZN => n17441);
   U177 : NAND4_X1 port map( A1 => n14328, A2 => n16442, A3 => n17520, A4 => 
                           n17441, ZN => n16443);
   U178 : NOR4_X1 port map( A1 => n13984, A2 => n18202, A3 => n16444, A4 => 
                           n16443, ZN => n16445);
   U179 : AOI211_X1 port map( C1 => n16447, C2 => n16446, A => n16445, B => 
                           n7822, ZN => n6095);
   U180 : NOR2_X1 port map( A1 => DATA1(13), A2 => n17788, ZN => n17593);
   U181 : INV_X1 port map( A => n17593, ZN => n17652);
   U182 : NAND2_X1 port map( A1 => DATA1(13), A2 => n17788, ZN => n17649);
   U183 : NAND2_X1 port map( A1 => n17652, A2 => n17649, ZN => n17542);
   U184 : AOI22_X1 port map( A1 => n6095, A2 => n14070, B1 => n18171, B2 => 
                           n17542, ZN => n16448);
   U185 : INV_X1 port map( A => n16448, ZN => n1851);
   U186 : NOR2_X1 port map( A1 => DATA2(21), A2 => n16606, ZN => n17674);
   U187 : INV_X1 port map( A => n17674, ZN => n16449);
   U188 : NAND2_X1 port map( A1 => DATA2(21), A2 => n16606, ZN => n17672);
   U189 : NAND2_X1 port map( A1 => n16449, A2 => n17672, ZN => n17544);
   U190 : AOI22_X1 port map( A1 => n6095, A2 => n14035, B1 => n18171, B2 => 
                           n17544, ZN => n16450);
   U191 : INV_X1 port map( A => n16450, ZN => n1849);
   U192 : INV_X1 port map( A => DATA1(23), ZN => n1882);
   U193 : INV_X1 port map( A => DATA1(25), ZN => n17275);
   U194 : XNOR2_X1 port map( A => DATA2_I_25_port, B => n17275, ZN => n17243);
   U195 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n17259);
   U196 : INV_X1 port map( A => n17259, ZN => n17256);
   U197 : XNOR2_X1 port map( A => DATA2_I_23_port, B => n1882, ZN => n17288);
   U198 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n17283);
   U199 : OAI21_X1 port map( B1 => DATA1(22), B2 => DATA2_I_22_port, A => 
                           n17283, ZN => n17300);
   U200 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, B1 => 
                           n1809, B2 => n18172, ZN => n17286);
   U201 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n17415);
   U202 : OAI21_X1 port map( B1 => DATA1(16), B2 => DATA2_I_16_port, A => 
                           n17415, ZN => n16720);
   U203 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => 
                           n16451, ZN => n17381);
   U204 : NOR4_X1 port map( A1 => n17392, A2 => n16452, A3 => n16720, A4 => 
                           n17381, ZN => n16454);
   U205 : NAND4_X1 port map( A1 => n17408, A2 => n1809, A3 => n16454, A4 => 
                           n16453, ZN => n16455);
   U206 : OAI221_X1 port map( B1 => n17300, B2 => n17286, C1 => n17300, C2 => 
                           n16455, A => n17283, ZN => n16456);
   U207 : AOI22_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, B1 => 
                           n17288, B2 => n16456, ZN => n16460);
   U208 : NOR2_X1 port map( A1 => n18230, A2 => n16460, ZN => n17260);
   U209 : NAND2_X1 port map( A1 => n17243, A2 => n17256, ZN => n16462);
   U210 : OAI211_X1 port map( C1 => n17243, C2 => n17256, A => n17260, B => 
                           n16462, ZN => n16457);
   U211 : INV_X1 port map( A => n16457, ZN => n8591);
   U212 : NOR2_X1 port map( A1 => n18230, A2 => n14460, ZN => n17537);
   U213 : INV_X1 port map( A => n17537, ZN => n1866);
   U214 : CLKBUF_X1 port map( A => n6095, Z => n17538);
   U215 : NOR2_X1 port map( A1 => DATA2(25), A2 => n17275, ZN => n17685);
   U216 : INV_X1 port map( A => n17685, ZN => n16458);
   U217 : NAND2_X1 port map( A1 => DATA2(25), A2 => n17275, ZN => n17686);
   U218 : NAND2_X1 port map( A1 => n16458, A2 => n17686, ZN => n17543);
   U219 : AOI22_X1 port map( A1 => n17538, A2 => n14023, B1 => n18171, B2 => 
                           n17543, ZN => n16459);
   U220 : INV_X1 port map( A => n16459, ZN => n1850);
   U221 : INV_X1 port map( A => DATA1(28), ZN => n17695);
   U222 : XNOR2_X1 port map( A => DATA2_I_28_port, B => n17695, ZN => n16467);
   U223 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n16465);
   U224 : INV_X1 port map( A => DATA1(27), ZN => n17209);
   U225 : XOR2_X1 port map( A => DATA2_I_27_port, B => n17209, Z => n17216);
   U226 : INV_X1 port map( A => n17216, ZN => n17214);
   U227 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n16464);
   U228 : INV_X1 port map( A => DATA1(26), ZN => n17689);
   U229 : XNOR2_X1 port map( A => DATA2_I_26_port, B => n17689, ZN => n17234);
   U230 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n16463);
   U231 : NAND3_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, A3 => 
                           n17243, ZN => n17242);
   U232 : NAND2_X1 port map( A1 => n16463, A2 => n17242, ZN => n17231);
   U233 : NAND2_X1 port map( A1 => n17234, A2 => n17231, ZN => n17230);
   U234 : NAND2_X1 port map( A1 => n16464, A2 => n17230, ZN => n17213);
   U235 : NAND2_X1 port map( A1 => n17214, A2 => n17213, ZN => n17211);
   U236 : NAND2_X1 port map( A1 => n16465, A2 => n17211, ZN => n16461);
   U237 : NAND2_X1 port map( A1 => n17769, A2 => n16460, ZN => n17182);
   U238 : INV_X1 port map( A => n17182, ZN => n17258);
   U239 : NAND2_X1 port map( A1 => n16467, A2 => n16461, ZN => n17181);
   U240 : OAI211_X1 port map( C1 => n16467, C2 => n16461, A => n17258, B => 
                           n17181, ZN => n16469);
   U241 : NAND2_X1 port map( A1 => n16463, A2 => n16462, ZN => n17233);
   U242 : NAND2_X1 port map( A1 => n17234, A2 => n17233, ZN => n17232);
   U243 : NAND2_X1 port map( A1 => n16464, A2 => n17232, ZN => n17220);
   U244 : NAND2_X1 port map( A1 => n17214, A2 => n17220, ZN => n17200);
   U245 : NAND2_X1 port map( A1 => n16465, A2 => n17200, ZN => n16466);
   U246 : NAND2_X1 port map( A1 => n16467, A2 => n16466, ZN => n17179);
   U247 : OAI211_X1 port map( C1 => n16467, C2 => n16466, A => n17260, B => 
                           n17179, ZN => n16468);
   U248 : AND2_X1 port map( A1 => n16469, A2 => n16468, ZN => n12229);
   U249 : INV_X1 port map( A => DATA1(1), ZN => n1891);
   U250 : INV_X1 port map( A => DATA1(0), ZN => n1892);
   U251 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN =>
                           n1823);
   U252 : INV_X1 port map( A => DATA1(4), ZN => n1890);
   U253 : INV_X1 port map( A => n9048, ZN => n1818);
   U254 : INV_X1 port map( A => n9045, ZN => n1816);
   U255 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN =>
                           n1842);
   U256 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN =>
                           n1840);
   U257 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN =>
                           n1838);
   U258 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN =>
                           n1836);
   U259 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN =>
                           n1833);
   U260 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN =>
                           n1831);
   U261 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN =>
                           n1829);
   U262 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN =>
                           n1827);
   U263 : INV_X1 port map( A => n9051, ZN => n1820);
   U264 : INV_X1 port map( A => n9054, ZN => n1822);
   U265 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN =>
                           n1825);
   U266 : INV_X1 port map( A => n9057, ZN => n1824);
   U267 : INV_X1 port map( A => n9060, ZN => n1826);
   U268 : INV_X1 port map( A => n9063, ZN => n1828);
   U269 : INV_X1 port map( A => n9075, ZN => n1837);
   U270 : INV_X1 port map( A => n9072, ZN => n1834);
   U271 : INV_X1 port map( A => n9069, ZN => n1832);
   U272 : INV_X1 port map( A => n9066, ZN => n1830);
   U273 : NAND2_X1 port map( A1 => DATA1(29), A2 => n4395, ZN => n17137);
   U274 : OAI21_X1 port map( B1 => DATA1(29), B2 => n4395, A => n17137, ZN => 
                           n8847);
   U275 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n17185);
   U276 : AOI21_X1 port map( B1 => n17185, B2 => n17181, A => n8847, ZN => 
                           n16999);
   U277 : AOI21_X1 port map( B1 => n17185, B2 => n17179, A => n8847, ZN => 
                           n16998);
   U278 : AOI22_X1 port map( A1 => n17258, A2 => n16999, B1 => n17260, B2 => 
                           n16998, ZN => n12162);
   U279 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n17002);
   U280 : OAI21_X1 port map( B1 => DATA1(30), B2 => DATA2_I_30_port, A => 
                           n17002, ZN => n11946);
   U281 : INV_X1 port map( A => DATA1(6), ZN => n1888);
   U282 : INV_X1 port map( A => n16488, ZN => n16470);
   U283 : OAI21_X1 port map( B1 => n18059, B2 => n18079, A => n16470, ZN => 
                           n16475);
   U284 : CLKBUF_X1 port map( A => n16475, Z => n16945);
   U285 : NAND3_X1 port map( A1 => DATA2(1), A2 => n17264, A3 => n18062, ZN => 
                           n17276);
   U286 : NOR2_X1 port map( A1 => n18161, A2 => n17000, ZN => n16471);
   U287 : OR2_X1 port map( A1 => n16978, A2 => n18078, ZN => n17192);
   U288 : NOR2_X1 port map( A1 => n17441, A2 => n17192, ZN => n16924);
   U289 : AOI211_X1 port map( C1 => DATA1(16), C2 => n16978, A => n16471, B => 
                           n16924, ZN => n16472);
   U290 : NAND2_X1 port map( A1 => DATA1(13), A2 => n17339, ZN => n16504);
   U291 : OAI211_X1 port map( C1 => n17276, C2 => n17655, A => n16472, B => 
                           n16504, ZN => n16600);
   U292 : NOR2_X1 port map( A1 => n16493, A2 => n17192, ZN => n16592);
   U293 : INV_X1 port map( A => n17000, ZN => n17713);
   U294 : CLKBUF_X1 port map( A => n17713, Z => n17345);
   U295 : NAND2_X1 port map( A1 => DATA1(10), A2 => n17345, ZN => n16473);
   U296 : INV_X1 port map( A => n17276, ZN => n17144);
   U297 : NAND2_X1 port map( A1 => DATA1(12), A2 => n17144, ZN => n16502);
   U298 : OAI211_X1 port map( C1 => n17264, C2 => n17655, A => n16473, B => 
                           n16502, ZN => n16474);
   U299 : AOI211_X1 port map( C1 => n17339, C2 => DATA1(11), A => n16592, B => 
                           n16474, ZN => n16489);
   U300 : INV_X1 port map( A => n16475, ZN => n17716);
   U301 : CLKBUF_X1 port map( A => n17716, Z => n17315);
   U302 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(0), ZN => n16687);
   U303 : AND2_X1 port map( A1 => n17315, A2 => n16687, ZN => n17352);
   U304 : CLKBUF_X1 port map( A => n17352, Z => n17305);
   U305 : INV_X1 port map( A => n17305, ZN => n17318);
   U306 : INV_X1 port map( A => n17339, ZN => n17348);
   U307 : NOR2_X1 port map( A1 => n18161, A2 => n17348, ZN => n16507);
   U308 : NAND2_X1 port map( A1 => DATA1(11), A2 => n17345, ZN => n16476);
   U309 : NAND2_X1 port map( A1 => DATA1(15), A2 => n16978, ZN => n16614);
   U310 : OAI211_X1 port map( C1 => n17276, C2 => n16493, A => n16476, B => 
                           n16614, ZN => n16477);
   U311 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(14), A => n16507, B => 
                           n16477, ZN => n16491);
   U312 : NOR3_X1 port map( A1 => n18079, A2 => n16488, A3 => n18069, ZN => 
                           n16492);
   U313 : INV_X1 port map( A => n16492, ZN => n17718);
   U314 : CLKBUF_X1 port map( A => n17718, Z => n17349);
   U315 : OAI22_X1 port map( A1 => n16489, A2 => n17318, B1 => n16491, B2 => 
                           n17349, ZN => n16478);
   U316 : AOI21_X1 port map( B1 => n16945, B2 => n16600, A => n16478, ZN => 
                           n18140);
   U317 : AOI21_X1 port map( B1 => DATA2(3), B2 => DATA2(1), A => n16653, ZN =>
                           n16479);
   U318 : INV_X1 port map( A => n16479, ZN => n18123);
   U319 : NAND3_X1 port map( A1 => n16479, A2 => n18066, A3 => n16488, ZN => 
                           n18152);
   U320 : NAND3_X1 port map( A1 => DATA2(3), A2 => n13099, A3 => n18083, ZN => 
                           n18150);
   U321 : CLKBUF_X1 port map( A => n18116, Z => n18114);
   U322 : INV_X1 port map( A => n17305, ZN => n17720);
   U323 : NOR2_X1 port map( A1 => n16514, A2 => n17000, ZN => n16482);
   U324 : NAND2_X1 port map( A1 => DATA1(10), A2 => n17339, ZN => n16480);
   U325 : NAND2_X1 port map( A1 => DATA1(11), A2 => n17144, ZN => n16508);
   U326 : OAI211_X1 port map( C1 => n17264, C2 => n16493, A => n16480, B => 
                           n16508, ZN => n16481);
   U327 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(12), A => n16482, B => 
                           n16481, ZN => n16490);
   U328 : OAI222_X1 port map( A1 => n17720, A2 => n16490, B1 => n17718, B2 => 
                           n16489, C1 => n17716, C2 => n16491, ZN => n18143);
   U329 : OAI21_X1 port map( B1 => DATA2(0), B2 => n16488, A => n16945, ZN => 
                           n16483);
   U330 : INV_X1 port map( A => n16483, ZN => n18137);
   U331 : AOI22_X1 port map( A1 => DATA1(10), A2 => n17279, B1 => n14469, B2 =>
                           n17339, ZN => n16484);
   U332 : NAND2_X1 port map( A1 => n17345, A2 => n14467, ZN => n16525);
   U333 : NAND2_X1 port map( A1 => DATA1(9), A2 => n17144, ZN => n16511);
   U334 : NAND2_X1 port map( A1 => DATA1(11), A2 => n16978, ZN => n16584);
   U335 : AND4_X1 port map( A1 => n16484, A2 => n16525, A3 => n16511, A4 => 
                           n16584, ZN => n16682);
   U336 : NOR2_X1 port map( A1 => n16514, A2 => n17348, ZN => n16485);
   U337 : NOR2_X1 port map( A1 => n17264, A2 => n18161, ZN => n16593);
   U338 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(11), A => n16485, B => 
                           n16593, ZN => n16486);
   U339 : NAND2_X1 port map( A1 => n14469, A2 => n17345, ZN => n16515);
   U340 : OAI211_X1 port map( C1 => n17276, C2 => n17520, A => n16486, B => 
                           n16515, ZN => n16487);
   U341 : INV_X1 port map( A => n16487, ZN => n16659);
   U342 : OAI222_X1 port map( A1 => n17720, A2 => n16682, B1 => n17718, B2 => 
                           n16659, C1 => n17716, C2 => n16490, ZN => n16905);
   U343 : AOI22_X1 port map( A1 => n18114, A2 => n18143, B1 => n18159, B2 => 
                           n16905, ZN => n16497);
   U344 : NOR2_X1 port map( A1 => n16488, A2 => n18159, ZN => n16531);
   U345 : CLKBUF_X1 port map( A => n16531, Z => n18118);
   U346 : OAI222_X1 port map( A1 => n17318, A2 => n16659, B1 => n17718, B2 => 
                           n16490, C1 => n17716, C2 => n16489, ZN => n16692);
   U347 : INV_X1 port map( A => n16491, ZN => n16495);
   U348 : CLKBUF_X1 port map( A => n16492, Z => n16942);
   U349 : INV_X1 port map( A => DATA1(16), ZN => n17423);
   U350 : NOR2_X1 port map( A1 => n17441, A2 => n17276, ZN => n16939);
   U351 : NOR2_X1 port map( A1 => n16493, A2 => n17000, ZN => n16506);
   U352 : AOI211_X1 port map( C1 => DATA1(17), C2 => n16978, A => n16939, B => 
                           n16506, ZN => n16494);
   U353 : NAND2_X1 port map( A1 => DATA1(14), A2 => n17339, ZN => n16582);
   U354 : OAI211_X1 port map( C1 => n17192, C2 => n17423, A => n16494, B => 
                           n16582, ZN => n16599);
   U355 : AOI222_X1 port map( A1 => n17305, A2 => n16495, B1 => n16942, B2 => 
                           n16600, C1 => n16945, C2 => n16599, ZN => n18084);
   U356 : INV_X1 port map( A => n18084, ZN => n16731);
   U357 : AOI22_X1 port map( A1 => n18118, A2 => n16692, B1 => n18123, B2 => 
                           n16731, ZN => n16496);
   U358 : OAI211_X1 port map( C1 => n18140, C2 => n18152, A => n16497, B => 
                           n16496, ZN => n1865);
   U359 : INV_X1 port map( A => DATA1(5), ZN => n1889);
   U360 : INV_X1 port map( A => DATA2(5), ZN => n17797);
   U361 : NAND4_X1 port map( A1 => n17572, A2 => n17797, A3 => FUNC(2), A4 => 
                           FUNC(1), ZN => n17540);
   U362 : INV_X1 port map( A => n17540, ZN => n16498);
   U363 : NOR2_X1 port map( A1 => n18079, A2 => n18077, ZN => n18068);
   U364 : NAND2_X1 port map( A1 => n18060, A2 => n18068, ZN => n17539);
   U365 : NAND2_X1 port map( A1 => n16498, A2 => n17539, ZN => n16538);
   U366 : NOR2_X1 port map( A1 => n1870, A2 => n16538, ZN => n1869);
   U367 : NOR2_X1 port map( A1 => n16514, A2 => n17192, ZN => n16501);
   U368 : NAND2_X1 port map( A1 => n14469, A2 => n16978, ZN => n16660);
   U369 : NAND2_X1 port map( A1 => DATA1(10), A2 => n17144, ZN => n16499);
   U370 : OAI211_X1 port map( C1 => n17000, C2 => n18161, A => n16660, B => 
                           n16499, ZN => n16500);
   U371 : AOI211_X1 port map( C1 => n17339, C2 => DATA1(11), A => n16501, B => 
                           n16500, ZN => n16522);
   U372 : INV_X1 port map( A => n16522, ZN => n16518);
   U373 : NOR2_X1 port map( A1 => n17264, A2 => n17520, ZN => n16654);
   U374 : INV_X1 port map( A => n16502, ZN => n16503);
   U375 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(11), A => n16654, B => 
                           n16503, ZN => n16505);
   U376 : OAI211_X1 port map( C1 => n17000, C2 => n17655, A => n16505, B => 
                           n16504, ZN => n16594);
   U377 : NOR2_X1 port map( A1 => n17264, A2 => n16514, ZN => n16668);
   U378 : NOR3_X1 port map( A1 => n16668, A2 => n16507, A3 => n16506, ZN => 
                           n16509);
   U379 : OAI211_X1 port map( C1 => n17192, C2 => n17520, A => n16509, B => 
                           n16508, ZN => n16586);
   U380 : AOI222_X1 port map( A1 => n16518, A2 => n16945, B1 => n16594, B2 => 
                           n17352, C1 => n16586, C2 => n16942, ZN => n16967);
   U381 : NOR2_X1 port map( A1 => n16393, A2 => n17276, ZN => n16670);
   U382 : NOR2_X1 port map( A1 => n14453, A2 => n17264, ZN => n17344);
   U383 : AOI211_X1 port map( C1 => n17339, C2 => n14469, A => n16670, B => 
                           n17344, ZN => n16510);
   U384 : NAND2_X1 port map( A1 => n14466, A2 => n17279, ZN => n16678);
   U385 : OAI211_X1 port map( C1 => n17000, C2 => n16514, A => n16510, B => 
                           n16678, ZN => n16530);
   U386 : NOR2_X1 port map( A1 => n18193, A2 => n17192, ZN => n16669);
   U387 : NOR2_X1 port map( A1 => n16393, A2 => n17264, ZN => n16676);
   U388 : AOI211_X1 port map( C1 => n17713, C2 => DATA1(11), A => n16669, B => 
                           n16676, ZN => n16512);
   U389 : OAI211_X1 port map( C1 => n17348, C2 => n17520, A => n16512, B => 
                           n16511, ZN => n16519);
   U390 : NOR2_X1 port map( A1 => n18193, A2 => n17276, ZN => n16655);
   U391 : NOR2_X1 port map( A1 => n14437, A2 => n17264, ZN => n16671);
   U392 : AOI211_X1 port map( C1 => n17713, C2 => DATA1(10), A => n16655, B => 
                           n16671, ZN => n16513);
   U393 : NAND2_X1 port map( A1 => n17279, A2 => n14467, ZN => n16661);
   U394 : OAI211_X1 port map( C1 => n17348, C2 => n16514, A => n16513, B => 
                           n16661, ZN => n16520);
   U395 : AOI222_X1 port map( A1 => n16530, A2 => n16945, B1 => n16519, B2 => 
                           n17352, C1 => n16520, C2 => n16942, ZN => n18151);
   U396 : INV_X1 port map( A => n18151, ZN => n16632);
   U397 : NOR2_X1 port map( A1 => n16393, A2 => n17348, ZN => n16656);
   U398 : INV_X1 port map( A => n16978, ZN => n17710);
   U399 : NAND2_X1 port map( A1 => n14465, A2 => n17279, ZN => n16673);
   U400 : OAI211_X1 port map( C1 => n14438, C2 => n17710, A => n16515, B => 
                           n16673, ZN => n16516);
   U401 : AOI211_X1 port map( C1 => n17144, C2 => n14466, A => n16656, B => 
                           n16516, ZN => n16528);
   U402 : INV_X1 port map( A => n16528, ZN => n16517);
   U403 : AOI222_X1 port map( A1 => n16517, A2 => n16945, B1 => n16520, B2 => 
                           n17352, C1 => n16530, C2 => n16942, ZN => n18153);
   U404 : INV_X1 port map( A => n18153, ZN => n16633);
   U405 : AOI22_X1 port map( A1 => n18144, A2 => n16632, B1 => n18123, B2 => 
                           n16633, ZN => n16524);
   U406 : AOI222_X1 port map( A1 => n16519, A2 => n16945, B1 => n16586, B2 => 
                           n17352, C1 => n16518, C2 => n16942, ZN => n16968);
   U407 : INV_X1 port map( A => n16968, ZN => n18158);
   U408 : AOI22_X1 port map( A1 => n16945, A2 => n16520, B1 => n16942, B2 => 
                           n16519, ZN => n16521);
   U409 : OAI21_X1 port map( B1 => n16522, B2 => n17720, A => n16521, ZN => 
                           n18147);
   U410 : AOI22_X1 port map( A1 => n18118, A2 => n18158, B1 => n18116, B2 => 
                           n18147, ZN => n16523);
   U411 : OAI211_X1 port map( C1 => n18137, C2 => n16967, A => n16524, B => 
                           n16523, ZN => n1853);
   U412 : NOR2_X1 port map( A1 => n14438, A2 => n17192, ZN => n17343);
   U413 : NAND2_X1 port map( A1 => n14466, A2 => n17339, ZN => n16665);
   U414 : OAI211_X1 port map( C1 => n14449, C2 => n17264, A => n16525, B => 
                           n16665, ZN => n16526);
   U415 : AOI211_X1 port map( C1 => n17144, C2 => n18213, A => n17343, B => 
                           n16526, ZN => n16533);
   U416 : NOR2_X1 port map( A1 => n14437, A2 => n17000, ZN => n16657);
   U417 : NAND2_X1 port map( A1 => n17279, A2 => n18206, ZN => n17708);
   U418 : NAND2_X1 port map( A1 => n17339, A2 => n18213, ZN => n16663);
   U419 : OAI211_X1 port map( C1 => n14438, C2 => n17276, A => n17708, B => 
                           n16663, ZN => n16527);
   U420 : AOI211_X1 port map( C1 => n14336, C2 => n16978, A => n16657, B => 
                           n16527, ZN => n16535);
   U421 : OAI222_X1 port map( A1 => n17318, A2 => n16528, B1 => n17718, B2 => 
                           n16533, C1 => n17716, C2 => n16535, ZN => n16802);
   U422 : OAI22_X1 port map( A1 => n16533, A2 => n17315, B1 => n16528, B2 => 
                           n17349, ZN => n16529);
   U423 : AOI21_X1 port map( B1 => n17352, B2 => n16530, A => n16529, ZN => 
                           n18154);
   U424 : INV_X1 port map( A => n16531, ZN => n18148);
   U425 : CLKBUF_X1 port map( A => n18148, Z => n18138);
   U426 : OAI22_X1 port map( A1 => n18137, A2 => n18153, B1 => n18154, B2 => 
                           n18138, ZN => n16537);
   U427 : NOR2_X1 port map( A1 => n14438, A2 => n17348, ZN => n16680);
   U428 : NAND2_X1 port map( A1 => n14465, A2 => n17345, ZN => n16666);
   U429 : NAND2_X1 port map( A1 => n17144, A2 => n18206, ZN => n17346);
   U430 : OAI211_X1 port map( C1 => n14328, C2 => n17710, A => n16666, B => 
                           n17346, ZN => n16532);
   U431 : AOI211_X1 port map( C1 => n17279, C2 => n14327, A => n16680, B => 
                           n16532, ZN => n16846);
   U432 : OAI222_X1 port map( A1 => n17720, A2 => n16533, B1 => n17718, B2 => 
                           n16535, C1 => n17716, C2 => n16846, ZN => n16800);
   U433 : INV_X1 port map( A => n16800, ZN => n16825);
   U434 : NOR2_X1 port map( A1 => n14451, A2 => n17276, ZN => n17712);
   U435 : NAND2_X1 port map( A1 => n14464, A2 => n17345, ZN => n16662);
   U436 : NAND2_X1 port map( A1 => n17339, A2 => n18206, ZN => n16674);
   U437 : OAI211_X1 port map( C1 => n14329, C2 => n17710, A => n16662, B => 
                           n16674, ZN => n16534);
   U438 : AOI211_X1 port map( C1 => n17279, C2 => n14463, A => n17712, B => 
                           n16534, ZN => n16879);
   U439 : OAI222_X1 port map( A1 => n17318, A2 => n16535, B1 => n17349, B2 => 
                           n16846, C1 => n17315, C2 => n16879, ZN => n16801);
   U440 : INV_X1 port map( A => n16801, ZN => n16824);
   U441 : OAI22_X1 port map( A1 => n16825, A2 => n18152, B1 => n16824, B2 => 
                           n18155, ZN => n16536);
   U442 : AOI211_X1 port map( C1 => n18114, C2 => n16802, A => n16537, B => 
                           n16536, ZN => n12526);
   U443 : NOR2_X1 port map( A1 => FUNC(3), A2 => n16538, ZN => n1868);
   U444 : INV_X1 port map( A => n1868, ZN => n16878);
   U445 : INV_X1 port map( A => n1897, ZN => n17499);
   U446 : OR3_X1 port map( A1 => n16878, A2 => n17499, A3 => n12526, ZN => 
                           n12527);
   U447 : NOR2_X1 port map( A1 => n17689, A2 => n17348, ZN => n17249);
   U448 : NOR2_X1 port map( A1 => n17275, A2 => n17276, ZN => n16540);
   U449 : NOR2_X1 port map( A1 => n17264, A2 => n1882, ZN => n16563);
   U450 : INV_X1 port map( A => DATA1(24), ZN => n17683);
   U451 : NAND2_X1 port map( A1 => DATA1(27), A2 => n17713, ZN => n17204);
   U452 : OAI21_X1 port map( B1 => n17192, B2 => n17683, A => n17204, ZN => 
                           n16539);
   U453 : NOR4_X1 port map( A1 => n17249, A2 => n16540, A3 => n16563, A4 => 
                           n16539, ZN => n16955);
   U454 : NOR2_X1 port map( A1 => n17275, A2 => n17348, ZN => n17266);
   U455 : NAND2_X1 port map( A1 => DATA1(26), A2 => n17345, ZN => n17225);
   U456 : NAND2_X1 port map( A1 => DATA1(22), A2 => n16978, ZN => n16541);
   U457 : NAND2_X1 port map( A1 => DATA1(23), A2 => n17279, ZN => n16559);
   U458 : NAND2_X1 port map( A1 => DATA1(24), A2 => n17144, ZN => n16642);
   U459 : NAND4_X1 port map( A1 => n17225, A2 => n16541, A3 => n16559, A4 => 
                           n16642, ZN => n16542);
   U460 : NOR2_X1 port map( A1 => n17266, A2 => n16542, ZN => n16550);
   U461 : INV_X1 port map( A => DATA1(22), ZN => n17675);
   U462 : NOR2_X1 port map( A1 => n17683, A2 => n17348, ZN => n17278);
   U463 : NOR2_X1 port map( A1 => n1882, A2 => n17276, ZN => n16637);
   U464 : AOI211_X1 port map( C1 => DATA1(21), C2 => n16978, A => n17278, B => 
                           n16637, ZN => n16543);
   U465 : NAND2_X1 port map( A1 => DATA1(25), A2 => n17345, ZN => n17245);
   U466 : OAI211_X1 port map( C1 => n17192, C2 => n17675, A => n16543, B => 
                           n17245, ZN => n16555);
   U467 : INV_X1 port map( A => n16555, ZN => n16549);
   U468 : OAI222_X1 port map( A1 => n17720, A2 => n16955, B1 => n17718, B2 => 
                           n16550, C1 => n17315, C2 => n16549, ZN => n16989);
   U469 : NOR2_X1 port map( A1 => n17209, A2 => n17348, ZN => n17228);
   U470 : NOR2_X1 port map( A1 => n17264, A2 => n17683, ZN => n16544);
   U471 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(25), A => n17228, B => 
                           n16544, ZN => n16545);
   U472 : NAND2_X1 port map( A1 => DATA1(26), A2 => n17144, ZN => n17263);
   U473 : OAI211_X1 port map( C1 => n17000, C2 => n17695, A => n16545, B => 
                           n17263, ZN => n16546);
   U474 : INV_X1 port map( A => n16546, ZN => n16963);
   U475 : OAI222_X1 port map( A1 => n16550, A2 => n17716, B1 => n16963, B2 => 
                           n17318, C1 => n16955, C2 => n17349, ZN => n16976);
   U476 : INV_X1 port map( A => n16976, ZN => n16960);
   U477 : NOR2_X1 port map( A1 => n17264, A2 => n16566, ZN => n16548);
   U478 : NOR2_X1 port map( A1 => n16606, A2 => n17192, ZN => n16561);
   U479 : NOR2_X1 port map( A1 => n1882, A2 => n17348, ZN => n16644);
   U480 : NAND2_X1 port map( A1 => DATA1(24), A2 => n17345, ZN => n17262);
   U481 : OAI21_X1 port map( B1 => n17276, B2 => n17675, A => n17262, ZN => 
                           n16547);
   U482 : NOR4_X1 port map( A1 => n16548, A2 => n16561, A3 => n16644, A4 => 
                           n16547, ZN => n16553);
   U483 : OAI222_X1 port map( A1 => n17720, A2 => n16550, B1 => n17718, B2 => 
                           n16549, C1 => n17315, C2 => n16553, ZN => n16957);
   U484 : INV_X1 port map( A => n16957, ZN => n16994);
   U485 : OAI22_X1 port map( A1 => n18137, A2 => n16960, B1 => n16994, B2 => 
                           n18150, ZN => n16557);
   U486 : INV_X1 port map( A => n18123, ZN => n18155);
   U487 : NAND2_X1 port map( A1 => DATA1(23), A2 => n17345, ZN => n17274);
   U488 : NAND2_X1 port map( A1 => DATA1(19), A2 => n16978, ZN => n16572);
   U489 : NAND2_X1 port map( A1 => DATA1(20), A2 => n17279, ZN => n16568);
   U490 : NAND2_X1 port map( A1 => DATA1(22), A2 => n17339, ZN => n16638);
   U491 : NAND4_X1 port map( A1 => n17274, A2 => n16572, A3 => n16568, A4 => 
                           n16638, ZN => n16551);
   U492 : AOI21_X1 port map( B1 => DATA1(21), B2 => n17144, A => n16551, ZN => 
                           n16610);
   U493 : NOR2_X1 port map( A1 => n16606, A2 => n17348, ZN => n16558);
   U494 : INV_X1 port map( A => DATA1(18), ZN => n17600);
   U495 : NAND2_X1 port map( A1 => DATA1(19), A2 => n17279, ZN => n16565);
   U496 : NAND2_X1 port map( A1 => DATA1(22), A2 => n17345, ZN => n16641);
   U497 : OAI211_X1 port map( C1 => n17264, C2 => n17600, A => n16565, B => 
                           n16641, ZN => n16552);
   U498 : AOI211_X1 port map( C1 => n17144, C2 => DATA1(20), A => n16558, B => 
                           n16552, ZN => n16626);
   U499 : OAI222_X1 port map( A1 => n17720, A2 => n16553, B1 => n17718, B2 => 
                           n16610, C1 => n17716, C2 => n16626, ZN => n16991);
   U500 : INV_X1 port map( A => n16991, ZN => n16623);
   U501 : OAI22_X1 port map( A1 => n16610, A2 => n17716, B1 => n16553, B2 => 
                           n17349, ZN => n16554);
   U502 : AOI21_X1 port map( B1 => n17352, B2 => n16555, A => n16554, ZN => 
                           n16956);
   U503 : OAI22_X1 port map( A1 => n18155, A2 => n16623, B1 => n16956, B2 => 
                           n18152, ZN => n16556);
   U504 : AOI211_X1 port map( C1 => n18118, C2 => n16989, A => n16557, B => 
                           n16556, ZN => n1873);
   U505 : NOR2_X1 port map( A1 => n16566, A2 => n17000, ZN => n16616);
   U506 : AOI211_X1 port map( C1 => DATA1(24), C2 => n16978, A => n16616, B => 
                           n16558, ZN => n16560);
   U507 : OAI211_X1 port map( C1 => n17276, C2 => n17675, A => n16560, B => 
                           n16559, ZN => n16645);
   U508 : NOR2_X1 port map( A1 => n17600, A2 => n17000, ZN => n16922);
   U509 : AOI211_X1 port map( C1 => DATA1(22), C2 => n16978, A => n16922, B => 
                           n16561, ZN => n16562);
   U510 : NAND2_X1 port map( A1 => DATA1(19), A2 => n17339, ZN => n16618);
   U511 : OAI211_X1 port map( C1 => n17276, C2 => n16566, A => n16562, B => 
                           n16618, ZN => n16570);
   U512 : INV_X1 port map( A => DATA1(19), ZN => n17379);
   U513 : NOR2_X1 port map( A1 => n17379, A2 => n17000, ZN => n16611);
   U514 : AOI211_X1 port map( C1 => n17144, C2 => DATA1(21), A => n16611, B => 
                           n16563, ZN => n16564);
   U515 : NAND2_X1 port map( A1 => DATA1(20), A2 => n17339, ZN => n16608);
   U516 : OAI211_X1 port map( C1 => n17192, C2 => n17675, A => n16564, B => 
                           n16608, ZN => n16640);
   U517 : AOI222_X1 port map( A1 => n16645, A2 => n16945, B1 => n16570, B2 => 
                           n17352, C1 => n16640, C2 => n16942, ZN => n18111);
   U518 : NOR2_X1 port map( A1 => n17600, A2 => n17276, ZN => n16617);
   U519 : NAND2_X1 port map( A1 => DATA1(16), A2 => n17345, ZN => n16589);
   U520 : OAI211_X1 port map( C1 => n17264, C2 => n16566, A => n16589, B => 
                           n16565, ZN => n16567);
   U521 : AOI211_X1 port map( C1 => n17339, C2 => DATA1(17), A => n16617, B => 
                           n16567, ZN => n16575);
   U522 : INV_X1 port map( A => n16575, ZN => n16578);
   U523 : NOR2_X1 port map( A1 => n17379, A2 => n17276, ZN => n16607);
   U524 : NAND2_X1 port map( A1 => DATA1(17), A2 => n17345, ZN => n16935);
   U525 : OAI211_X1 port map( C1 => n17264, C2 => n16606, A => n16935, B => 
                           n16568, ZN => n16569);
   U526 : AOI211_X1 port map( C1 => n17339, C2 => DATA1(18), A => n16607, B => 
                           n16569, ZN => n16574);
   U527 : INV_X1 port map( A => n16574, ZN => n16571);
   U528 : AOI222_X1 port map( A1 => n17352, A2 => n16578, B1 => n16942, B2 => 
                           n16571, C1 => n16945, C2 => n16570, ZN => n16739);
   U529 : INV_X1 port map( A => n16739, ZN => n16735);
   U530 : AOI222_X1 port map( A1 => n17352, A2 => n16571, B1 => n16942, B2 => 
                           n16570, C1 => n16945, C2 => n16640, ZN => n18107);
   U531 : INV_X1 port map( A => n18107, ZN => n16743);
   U532 : AOI22_X1 port map( A1 => n18114, A2 => n16735, B1 => n18144, B2 => 
                           n16743, ZN => n16581);
   U533 : NOR2_X1 port map( A1 => n17423, A2 => n17348, ZN => n16938);
   U534 : NAND2_X1 port map( A1 => DATA1(17), A2 => n17144, ZN => n16612);
   U535 : OAI211_X1 port map( C1 => n17000, C2 => n17441, A => n16572, B => 
                           n16612, ZN => n16573);
   U536 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(18), A => n16938, B => 
                           n16573, ZN => n16577);
   U537 : OAI222_X1 port map( A1 => n17720, A2 => n16577, B1 => n17718, B2 => 
                           n16575, C1 => n17716, C2 => n16574, ZN => n16736);
   U538 : NOR2_X1 port map( A1 => n17441, A2 => n17348, ZN => n16591);
   U539 : NOR2_X1 port map( A1 => n17423, A2 => n17276, ZN => n16923);
   U540 : AOI211_X1 port map( C1 => DATA1(18), C2 => n16978, A => n16591, B => 
                           n16923, ZN => n16576);
   U541 : NAND2_X1 port map( A1 => DATA1(17), A2 => n17279, ZN => n16619);
   U542 : OAI211_X1 port map( C1 => n17000, C2 => n17655, A => n16576, B => 
                           n16619, ZN => n16601);
   U543 : INV_X1 port map( A => n16577, ZN => n16598);
   U544 : AOI222_X1 port map( A1 => n17352, A2 => n16601, B1 => n16942, B2 => 
                           n16598, C1 => n16945, C2 => n16578, ZN => n16579);
   U545 : INV_X1 port map( A => n16579, ZN => n18089);
   U546 : AOI22_X1 port map( A1 => n18118, A2 => n16736, B1 => n18159, B2 => 
                           n18089, ZN => n16580);
   U547 : OAI211_X1 port map( C1 => n18155, C2 => n18111, A => n16581, B => 
                           n16580, ZN => n1880);
   U548 : AOI22_X1 port map( A1 => n18116, A2 => n18158, B1 => n18144, B2 => 
                           n18147, ZN => n16588);
   U549 : AOI22_X1 port map( A1 => DATA1(13), A2 => n17144, B1 => DATA1(15), B2
                           => n17713, ZN => n16585);
   U550 : NAND2_X1 port map( A1 => DATA1(12), A2 => n17279, ZN => n16583);
   U551 : NAND4_X1 port map( A1 => n16585, A2 => n16584, A3 => n16583, A4 => 
                           n16582, ZN => n16941);
   U552 : AOI222_X1 port map( A1 => n16586, A2 => n16945, B1 => n16941, B2 => 
                           n17352, C1 => n16594, C2 => n16942, ZN => n16970);
   U553 : INV_X1 port map( A => n16970, ZN => n16595);
   U554 : AOI22_X1 port map( A1 => n18159, A2 => n16595, B1 => n18123, B2 => 
                           n16632, ZN => n16587);
   U555 : OAI211_X1 port map( C1 => n16967, C2 => n18148, A => n16588, B => 
                           n16587, ZN => n1852);
   U556 : OAI21_X1 port map( B1 => n17276, B2 => n17655, A => n16589, ZN => 
                           n16590);
   U557 : OR4_X1 port map( A1 => n16593, A2 => n16592, A3 => n16591, A4 => 
                           n16590, ZN => n16940);
   U558 : AOI222_X1 port map( A1 => n16594, A2 => n16945, B1 => n16940, B2 => 
                           n17352, C1 => n16941, C2 => n16942, ZN => n16969);
   U559 : INV_X1 port map( A => n16969, ZN => n18090);
   U560 : AOI22_X1 port map( A1 => n18159, A2 => n18090, B1 => n18123, B2 => 
                           n18147, ZN => n16597);
   U561 : AOI22_X1 port map( A1 => n18118, A2 => n16595, B1 => n18144, B2 => 
                           n18158, ZN => n16596);
   U562 : OAI211_X1 port map( C1 => n16967, C2 => n18150, A => n16597, B => 
                           n16596, ZN => n1854);
   U563 : AOI222_X1 port map( A1 => n17352, A2 => n16599, B1 => n16942, B2 => 
                           n16601, C1 => n16945, C2 => n16598, ZN => n18085);
   U564 : OAI22_X1 port map( A1 => n18155, A2 => n16739, B1 => n18085, B2 => 
                           n18148, ZN => n16603);
   U565 : AOI222_X1 port map( A1 => n16601, A2 => n16945, B1 => n16600, B2 => 
                           n17352, C1 => n16599, C2 => n16942, ZN => n18086);
   U566 : INV_X1 port map( A => n16736, ZN => n16740);
   U567 : OAI22_X1 port map( A1 => n18137, A2 => n18086, B1 => n16740, B2 => 
                           n18152, ZN => n16602);
   U568 : AOI211_X1 port map( C1 => n18114, C2 => n18089, A => n16603, B => 
                           n16602, ZN => n1883);
   U569 : INV_X1 port map( A => n18143, ZN => n16629);
   U570 : OAI22_X1 port map( A1 => n18137, A2 => n16629, B1 => n18086, B2 => 
                           n18152, ZN => n16605);
   U571 : OAI22_X1 port map( A1 => n18155, A2 => n18085, B1 => n18140, B2 => 
                           n18148, ZN => n16604);
   U572 : AOI211_X1 port map( C1 => n18114, C2 => n16731, A => n16605, B => 
                           n16604, ZN => n1887);
   U573 : OR4_X1 port map( A1 => DATA1(5), A2 => DATA1(4), A3 => DATA1(0), A4 
                           => DATA1(3), ZN => n11540);
   U574 : NOR2_X1 port map( A1 => n16606, A2 => n17000, ZN => n16636);
   U575 : AOI211_X1 port map( C1 => DATA1(17), C2 => n16978, A => n16607, B => 
                           n16636, ZN => n16609);
   U576 : OAI211_X1 port map( C1 => n17192, C2 => n17600, A => n16609, B => 
                           n16608, ZN => n16622);
   U577 : INV_X1 port map( A => n16622, ZN => n16625);
   U578 : OAI222_X1 port map( A1 => n17720, A2 => n16610, B1 => n17718, B2 => 
                           n16626, C1 => n17716, C2 => n16625, ZN => n18102);
   U579 : AOI21_X1 port map( B1 => n17339, B2 => DATA1(18), A => n16611, ZN => 
                           n16615);
   U580 : NAND2_X1 port map( A1 => DATA1(16), A2 => n17279, ZN => n16613);
   U581 : NAND4_X1 port map( A1 => n16615, A2 => n16614, A3 => n16613, A4 => 
                           n16612, ZN => n16944);
   U582 : NOR2_X1 port map( A1 => n16617, A2 => n16616, ZN => n16621);
   U583 : NAND2_X1 port map( A1 => DATA1(16), A2 => n16978, ZN => n16620);
   U584 : NAND4_X1 port map( A1 => n16621, A2 => n16620, A3 => n16619, A4 => 
                           n16618, ZN => n16928);
   U585 : AOI222_X1 port map( A1 => n16944, A2 => n16945, B1 => n16622, B2 => 
                           n17352, C1 => n16928, C2 => n16942, ZN => n18099);
   U586 : OAI22_X1 port map( A1 => n18155, A2 => n18099, B1 => n16623, B2 => 
                           n18138, ZN => n16628);
   U587 : INV_X1 port map( A => n16928, ZN => n16624);
   U588 : OAI222_X1 port map( A1 => n17720, A2 => n16626, B1 => n17349, B2 => 
                           n16625, C1 => n17716, C2 => n16624, ZN => n18101);
   U589 : INV_X1 port map( A => n18101, ZN => n18096);
   U590 : OAI22_X1 port map( A1 => n18137, A2 => n16956, B1 => n18096, B2 => 
                           n18152, ZN => n16627);
   U591 : AOI211_X1 port map( C1 => n18114, C2 => n18102, A => n16628, B => 
                           n16627, ZN => n1879);
   U592 : INV_X1 port map( A => n16692, ZN => n18135);
   U593 : OAI22_X1 port map( A1 => n18137, A2 => n18135, B1 => n16629, B2 => 
                           n18138, ZN => n16631);
   U594 : OAI22_X1 port map( A1 => n18155, A2 => n18086, B1 => n18140, B2 => 
                           n18150, ZN => n16630);
   U595 : AOI211_X1 port map( C1 => n18144, C2 => n16731, A => n16631, B => 
                           n16630, ZN => n8647);
   U596 : AOI22_X1 port map( A1 => n18118, A2 => n16632, B1 => n18159, B2 => 
                           n18147, ZN => n16635);
   U597 : AOI22_X1 port map( A1 => n18116, A2 => n16633, B1 => n16802, B2 => 
                           n18123, ZN => n16634);
   U598 : OAI211_X1 port map( C1 => n18154, C2 => n18152, A => n16635, B => 
                           n16634, ZN => n1857);
   U599 : AOI211_X1 port map( C1 => DATA1(25), C2 => n16978, A => n16637, B => 
                           n16636, ZN => n16639);
   U600 : OAI211_X1 port map( C1 => n17192, C2 => n17683, A => n16639, B => 
                           n16638, ZN => n17313);
   U601 : AOI222_X1 port map( A1 => n17313, A2 => n16945, B1 => n16640, B2 => 
                           n17352, C1 => n16645, C2 => n16942, ZN => n18110);
   U602 : INV_X1 port map( A => n18110, ZN => n18117);
   U603 : OAI211_X1 port map( C1 => n17264, C2 => n17689, A => n16642, B => 
                           n16641, ZN => n16643);
   U604 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(25), A => n16644, B => 
                           n16643, ZN => n17316);
   U605 : AOI22_X1 port map( A1 => n17305, A2 => n16645, B1 => n16942, B2 => 
                           n17313, ZN => n16646);
   U606 : OAI21_X1 port map( B1 => n17316, B2 => n17716, A => n16646, ZN => 
                           n18125);
   U607 : AOI22_X1 port map( A1 => n18159, A2 => n16735, B1 => n18123, B2 => 
                           n18125, ZN => n16647);
   U608 : INV_X1 port map( A => n16647, ZN => n16649);
   U609 : OAI22_X1 port map( A1 => n18138, A2 => n18107, B1 => n18150, B2 => 
                           n18111, ZN => n16648);
   U610 : AOI211_X1 port map( C1 => n18117, C2 => n18144, A => n16649, B => 
                           n16648, ZN => n16745);
   U611 : INV_X1 port map( A => n16745, ZN => n1877);
   U612 : OAI22_X1 port map( A1 => n18137, A2 => n18151, B1 => n18153, B2 => 
                           n18138, ZN => n16651);
   U613 : OAI22_X1 port map( A1 => n16825, A2 => n18155, B1 => n18154, B2 => 
                           n18150, ZN => n16650);
   U614 : AOI211_X1 port map( C1 => n18144, C2 => n16802, A => n16651, B => 
                           n16650, ZN => n8604);
   U615 : AOI21_X1 port map( B1 => n13099, B2 => n18059, A => n16652, ZN => 
                           n13151);
   U616 : INV_X1 port map( A => n13151, ZN => n1895);
   U617 : NAND3_X1 port map( A1 => n16687, A2 => n1895, A3 => n16653, ZN => 
                           n1896);
   U618 : INV_X1 port map( A => n1896, ZN => n11927);
   U619 : OR4_X1 port map( A1 => n16657, A2 => n16656, A3 => n16655, A4 => 
                           n16654, ZN => n16658);
   U620 : AOI21_X1 port map( B1 => DATA1(9), B2 => n17279, A => n16658, ZN => 
                           n16683);
   U621 : OAI222_X1 port map( A1 => n16659, A2 => n17716, B1 => n16683, B2 => 
                           n17318, C1 => n16682, C2 => n17349, ZN => n16688);
   U622 : INV_X1 port map( A => n16688, ZN => n18136);
   U623 : NAND4_X1 port map( A1 => n16663, A2 => n16662, A3 => n16661, A4 => 
                           n16660, ZN => n16664);
   U624 : AOI21_X1 port map( B1 => n14466, B2 => n17144, A => n16664, ZN => 
                           n16681);
   U625 : NAND2_X1 port map( A1 => n16666, A2 => n16665, ZN => n16667);
   U626 : NOR4_X1 port map( A1 => n16670, A2 => n16669, A3 => n16668, A4 => 
                           n16667, ZN => n16684);
   U627 : OAI222_X1 port map( A1 => n17720, A2 => n16681, B1 => n17718, B2 => 
                           n16684, C1 => n17716, C2 => n16683, ZN => n17723);
   U628 : NOR2_X1 port map( A1 => n14451, A2 => n17000, ZN => n17143);
   U629 : INV_X1 port map( A => n16671, ZN => n16672);
   U630 : NAND3_X1 port map( A1 => n16674, A2 => n16673, A3 => n16672, ZN => 
                           n16675);
   U631 : AOI211_X1 port map( C1 => n17144, C2 => n14464, A => n17143, B => 
                           n16675, ZN => n17715);
   U632 : INV_X1 port map( A => n16676, ZN => n16677);
   U633 : OAI211_X1 port map( C1 => n17276, C2 => n18219, A => n16678, B => 
                           n16677, ZN => n16679);
   U634 : AOI211_X1 port map( C1 => n17713, C2 => n14326, A => n16680, B => 
                           n16679, ZN => n17350);
   U635 : OAI222_X1 port map( A1 => n17318, A2 => n17715, B1 => n17349, B2 => 
                           n17350, C1 => n17315, C2 => n16681, ZN => n17722);
   U636 : AOI22_X1 port map( A1 => n18114, A2 => n17723, B1 => n18159, B2 => 
                           n17722, ZN => n16686);
   U637 : OAI222_X1 port map( A1 => n17720, A2 => n17350, B1 => n17718, B2 => 
                           n16681, C1 => n17716, C2 => n16684, ZN => n17724);
   U638 : OAI222_X1 port map( A1 => n17720, A2 => n16684, B1 => n17718, B2 => 
                           n16683, C1 => n17315, C2 => n16682, ZN => n16691);
   U639 : AOI22_X1 port map( A1 => n18118, A2 => n17724, B1 => n18144, B2 => 
                           n16691, ZN => n16685);
   U640 : OAI211_X1 port map( C1 => n18155, C2 => n18136, A => n16686, B => 
                           n16685, ZN => n1861);
   U641 : NOR3_X2 port map( A1 => n13151, A2 => n16687, A3 => n18082, ZN => 
                           n1894);
   U642 : INV_X1 port map( A => n1894, ZN => n9020);
   U643 : INV_X1 port map( A => n16691, ZN => n17355);
   U644 : AOI22_X1 port map( A1 => n18114, A2 => n16688, B1 => n18159, B2 => 
                           n17723, ZN => n16690);
   U645 : AOI22_X1 port map( A1 => n18144, A2 => n16905, B1 => n18123, B2 => 
                           n16692, ZN => n16689);
   U646 : OAI211_X1 port map( C1 => n17355, C2 => n18148, A => n16690, B => 
                           n16689, ZN => n1862);
   U647 : AOI22_X1 port map( A1 => n18114, A2 => n16905, B1 => n18159, B2 => 
                           n16691, ZN => n16694);
   U648 : AOI22_X1 port map( A1 => n18144, A2 => n16692, B1 => n18123, B2 => 
                           n18143, ZN => n16693);
   U649 : OAI211_X1 port map( C1 => n18136, C2 => n18148, A => n16694, B => 
                           n16693, ZN => n1859);
   U650 : NAND3_X1 port map( A1 => DATA2(3), A2 => n13099, A3 => n18063, ZN => 
                           n17728);
   U651 : INV_X1 port map( A => n17728, ZN => n1898);
   U652 : AOI211_X1 port map( C1 => n14365, C2 => n14337, A => n13947, B => 
                           n13946, ZN => n16707);
   U653 : AOI22_X1 port map( A1 => n16399, A2 => n14383, B1 => n13962, B2 => 
                           n14186, ZN => n16696);
   U654 : AOI22_X1 port map( A1 => n14187, A2 => n14411, B1 => n14430, B2 => 
                           n14434, ZN => n16695);
   U655 : OAI211_X1 port map( C1 => n13963, C2 => n14226, A => n16696, B => 
                           n16695, ZN => n16697);
   U656 : INV_X1 port map( A => n16697, ZN => n16710);
   U657 : AOI22_X1 port map( A1 => n14334, A2 => n14410, B1 => n16399, B2 => 
                           n18185, ZN => n16700);
   U658 : OAI22_X1 port map( A1 => n14454, A2 => n13963, B1 => n14231, B2 => 
                           n13951, ZN => n16698);
   U659 : INV_X1 port map( A => n16698, ZN => n16699);
   U660 : OAI211_X1 port map( C1 => n14274, C2 => n14409, A => n16700, B => 
                           n16699, ZN => n16701);
   U661 : INV_X1 port map( A => n16701, ZN => n17013);
   U662 : OAI222_X1 port map( A1 => n14374, A2 => n16707, B1 => n16710, B2 => 
                           n14228, C1 => n14455, C2 => n17013, ZN => n17051);
   U663 : INV_X1 port map( A => n17051, ZN => n17059);
   U664 : OAI22_X1 port map( A1 => n14409, A2 => n14231, B1 => n14436, B2 => 
                           n14412, ZN => n16702);
   U665 : AOI211_X1 port map( C1 => n14337, C2 => n14364, A => n13945, B => 
                           n16702, ZN => n16708);
   U666 : OAI22_X1 port map( A1 => n14228, A2 => n16707, B1 => n14374, B2 => 
                           n16708, ZN => n16703);
   U667 : INV_X1 port map( A => n16703, ZN => n16704);
   U668 : OAI21_X1 port map( B1 => n14455, B2 => n16710, A => n16704, ZN => 
                           n17385);
   U669 : OAI22_X1 port map( A1 => n14226, A2 => n13891, B1 => n14349, B2 => 
                           n14412, ZN => n16705);
   U670 : AOI211_X1 port map( C1 => n14337, C2 => n14363, A => n13944, B => 
                           n16705, ZN => n16714);
   U671 : OAI22_X1 port map( A1 => n14454, A2 => n14412, B1 => n14231, B2 => 
                           n13891, ZN => n16706);
   U672 : AOI211_X1 port map( C1 => n14364, C2 => n14392, A => n13943, B => 
                           n16706, ZN => n17450);
   U673 : OAI222_X1 port map( A1 => n14228, A2 => n16714, B1 => n14455, B2 => 
                           n16708, C1 => n14374, C2 => n17450, ZN => n17417);
   U674 : AOI22_X1 port map( A1 => n13893, A2 => n17385, B1 => n14220, B2 => 
                           n17417, ZN => n16712);
   U675 : OAI222_X1 port map( A1 => n14228, A2 => n16708, B1 => n14455, B2 => 
                           n16707, C1 => n14374, C2 => n16714, ZN => n17403);
   U676 : OAI22_X1 port map( A1 => n14231, A2 => n13952, B1 => n13951, B2 => 
                           n14226, ZN => n16709);
   U677 : AOI211_X1 port map( C1 => n14187, C2 => n13962, A => n13950, B => 
                           n16709, ZN => n17024);
   U678 : OAI222_X1 port map( A1 => n14374, A2 => n16710, B1 => n17013, B2 => 
                           n14228, C1 => n17024, C2 => n14455, ZN => n17055);
   U679 : AOI22_X1 port map( A1 => n14395, A2 => n17403, B1 => n14130, B2 => 
                           n17055, ZN => n16711);
   U680 : OAI211_X1 port map( C1 => n14134, C2 => n17059, A => n16712, B => 
                           n16711, ZN => n17121);
   U681 : AOI22_X1 port map( A1 => n14340, A2 => n14337, B1 => n14393, B2 => 
                           n13961, ZN => n16713);
   U682 : OAI211_X1 port map( C1 => n14436, C2 => n13939, A => n14423, B => 
                           n16713, ZN => n17452);
   U683 : INV_X1 port map( A => n17452, ZN => n17470);
   U684 : OAI222_X1 port map( A1 => n14228, A2 => n17450, B1 => n14455, B2 => 
                           n16714, C1 => n14374, C2 => n17470, ZN => n17429);
   U685 : AOI22_X1 port map( A1 => n14220, A2 => n17429, B1 => n14395, B2 => 
                           n17417, ZN => n16716);
   U686 : AOI22_X1 port map( A1 => n13893, A2 => n17403, B1 => n18181, B2 => 
                           n17385, ZN => n16715);
   U687 : OAI211_X1 port map( C1 => n17059, C2 => n14389, A => n16716, B => 
                           n16715, ZN => n17332);
   U688 : AOI22_X1 port map( A1 => n18189, A2 => n17121, B1 => n18209, B2 => 
                           n17332, ZN => n16717);
   U689 : OAI22_X1 port map( A1 => n14378, A2 => n14452, B1 => n16717, B2 => 
                           n18212, ZN => n16718);
   U690 : OR4_X1 port map( A1 => n13923, A2 => n14414, A3 => n18229, A4 => 
                           n16718, ZN => OUTALU(21));
   U691 : INV_X1 port map( A => n4302, ZN => n1845);
   U692 : INV_X1 port map( A => n9084, ZN => n1843);
   U693 : INV_X1 port map( A => n9081, ZN => n1841);
   U694 : INV_X1 port map( A => n1846, ZN => n18071);
   U695 : NOR2_X1 port map( A1 => n1845, A2 => n18071, ZN => n12924);
   U696 : INV_X1 port map( A => n1848, ZN => n18074);
   U697 : NOR2_X1 port map( A1 => n7769, A2 => n18074, ZN => n1847);
   U698 : INV_X1 port map( A => n8814, ZN => n16719);
   U699 : NOR2_X1 port map( A1 => n16719, A2 => n1847, ZN => n8929);
   U700 : INV_X1 port map( A => n16720, ZN => n17425);
   U701 : NOR2_X1 port map( A1 => n17425, A2 => n17409, ZN => n8943);
   U702 : NAND2_X1 port map( A1 => n17769, A2 => n14460, ZN => n17335);
   U703 : INV_X1 port map( A => n17335, ZN => n17533);
   U704 : INV_X1 port map( A => n16855, ZN => n16852);
   U705 : INV_X1 port map( A => n16721, ZN => n16725);
   U706 : INV_X1 port map( A => n17336, ZN => n16722);
   U707 : AOI21_X1 port map( B1 => n16724, B2 => n16722, A => n17150, ZN => 
                           n17148);
   U708 : NOR2_X1 port map( A1 => n16725, A2 => n17148, ZN => n16903);
   U709 : INV_X1 port map( A => n16723, ZN => n18056);
   U710 : NOR2_X1 port map( A1 => n16903, A2 => n18056, ZN => n16902);
   U711 : NOR2_X1 port map( A1 => n16726, A2 => n16902, ZN => n16885);
   U712 : OAI21_X1 port map( B1 => n16885, B2 => n1429, A => n16727, ZN => 
                           n16851);
   U713 : AOI21_X1 port map( B1 => n16852, B2 => n16851, A => n16728, ZN => 
                           n16843);
   U714 : INV_X1 port map( A => n17340, ZN => n17342);
   U715 : INV_X1 port map( A => n16724, ZN => n17147);
   U716 : AOI21_X1 port map( B1 => n17532, B2 => n17342, A => n17147, ZN => 
                           n17146);
   U717 : NOR2_X1 port map( A1 => n17146, A2 => n17150, ZN => n17145);
   U718 : NOR2_X1 port map( A1 => n16725, A2 => n17145, ZN => n18057);
   U719 : NOR2_X1 port map( A1 => n18057, A2 => n18056, ZN => n18055);
   U720 : NOR2_X1 port map( A1 => n16726, A2 => n18055, ZN => n16884);
   U721 : OAI21_X1 port map( B1 => n16884, B2 => n1429, A => n16727, ZN => 
                           n16850);
   U722 : AOI21_X1 port map( B1 => n16852, B2 => n16850, A => n16728, ZN => 
                           n16842);
   U723 : AOI22_X1 port map( A1 => n17533, A2 => n16843, B1 => n17537, B2 => 
                           n16842, ZN => n16730);
   U724 : NAND3_X1 port map( A1 => n1868, A2 => n18159, A3 => n16801, ZN => 
                           n16729);
   U725 : OAI21_X1 port map( B1 => n16730, B2 => n16845, A => n16729, ZN => 
                           n11526);
   U726 : AOI22_X1 port map( A1 => n18144, A2 => n18089, B1 => n18159, B2 => 
                           n16731, ZN => n16734);
   U727 : INV_X1 port map( A => n18085, ZN => n16732);
   U728 : AOI22_X1 port map( A1 => n18116, A2 => n16732, B1 => n18123, B2 => 
                           n16736, ZN => n16733);
   U729 : OAI211_X1 port map( C1 => n18086, C2 => n18148, A => n16734, B => 
                           n16733, ZN => n11473);
   U730 : AOI22_X1 port map( A1 => n1897, A2 => n11473, B1 => n1894, B2 => 
                           n1880, ZN => n11436);
   U731 : AOI22_X1 port map( A1 => n18118, A2 => n18089, B1 => n18144, B2 => 
                           n16735, ZN => n16738);
   U732 : AOI22_X1 port map( A1 => n18114, A2 => n16736, B1 => n18123, B2 => 
                           n16743, ZN => n16737);
   U733 : OAI211_X1 port map( C1 => n18137, C2 => n18085, A => n16738, B => 
                           n16737, ZN => n11457);
   U734 : INV_X1 port map( A => n1883, ZN => n16746);
   U735 : AOI22_X1 port map( A1 => n1898, A2 => n16746, B1 => n11927, B2 => 
                           n11457, ZN => n11435);
   U736 : OAI22_X1 port map( A1 => n18155, A2 => n18110, B1 => n18111, B2 => 
                           n18152, ZN => n16742);
   U737 : OAI22_X1 port map( A1 => n18137, A2 => n16740, B1 => n16739, B2 => 
                           n18148, ZN => n16741);
   U738 : AOI211_X1 port map( C1 => n18114, C2 => n16743, A => n16742, B => 
                           n16741, ZN => n11449);
   U739 : INV_X1 port map( A => n1880, ZN => n16744);
   U740 : OAI22_X1 port map( A1 => n16744, A2 => n1896, B1 => n11449, B2 => 
                           n9020, ZN => n11437);
   U741 : OAI22_X1 port map( A1 => n11449, A2 => n17499, B1 => n16745, B2 => 
                           n17728, ZN => n11444);
   U742 : OAI22_X1 port map( A1 => n16744, A2 => n17728, B1 => n11449, B2 => 
                           n1896, ZN => n11447);
   U743 : OAI22_X1 port map( A1 => n11449, A2 => n17728, B1 => n16745, B2 => 
                           n1896, ZN => n11453);
   U744 : INV_X1 port map( A => n1887, ZN => n16856);
   U745 : AOI22_X1 port map( A1 => n1897, A2 => n16856, B1 => n1894, B2 => 
                           n16746, ZN => n11459);
   U746 : AOI22_X1 port map( A1 => n13151, A2 => n11457, B1 => n11927, B2 => 
                           n11473, ZN => n11458);
   U747 : INV_X1 port map( A => n1865, ZN => n16747);
   U748 : OAI22_X1 port map( A1 => n8647, A2 => n17728, B1 => n16747, B2 => 
                           n17499, ZN => n11469);
   U749 : OAI22_X1 port map( A1 => n8647, A2 => n1896, B1 => n16747, B2 => 
                           n17728, ZN => n11485);
   U750 : INV_X1 port map( A => n17530, ZN => n17518);
   U751 : INV_X1 port map( A => n17424, ZN => n17517);
   U752 : NOR2_X1 port map( A1 => n17518, A2 => n17517, ZN => n18162);
   U753 : INV_X1 port map( A => DATA2(22), ZN => n17779);
   U754 : NOR3_X1 port map( A1 => n18162, A2 => n17779, A3 => n17675, ZN => 
                           n8892);
   U755 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n18073, ZN => n2808);
   U756 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n2808, ZN => n8887);
   U757 : NOR3_X1 port map( A1 => n14459, A2 => n14132, A3 => n1844, ZN => 
                           n3026);
   U758 : AOI221_X1 port map( B1 => n14132, B2 => n14459, C1 => n1844, C2 => 
                           n14459, A => n3026, ZN => n8555);
   U759 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, ZN => 
                           n16748);
   U760 : NOR3_X1 port map( A1 => n14189, A2 => n1844, A3 => n16748, ZN => 
                           n3030);
   U761 : AOI221_X1 port map( B1 => n14189, B2 => n16748, C1 => n1844, C2 => 
                           n16748, A => n3030, ZN => n8880);
   U762 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_4_8_port, ZN => 
                           n16749);
   U763 : NOR3_X1 port map( A1 => n14181, A2 => n1844, A3 => n16749, ZN => 
                           n3029);
   U764 : AOI21_X1 port map( B1 => n14433, B2 => data1_mul_0_port, A => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, ZN => n16750
                           );
   U765 : NOR2_X1 port map( A1 => n3029, A2 => n16750, ZN => n8875);
   U766 : NAND2_X1 port map( A1 => n16410, A2 => n14286, ZN => n16751);
   U767 : OAI21_X1 port map( B1 => n16410, B2 => n14286, A => n16751, ZN => 
                           n17932);
   U768 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_5_10_port, ZN => 
                           n16752);
   U769 : NOR3_X1 port map( A1 => n1844, A2 => n17932, A3 => n16752, ZN => 
                           n3028);
   U770 : OR2_X1 port map( A1 => n1844, A2 => n17932, ZN => n16753);
   U771 : AOI21_X1 port map( B1 => n16753, B2 => n16752, A => n3028, ZN => 
                           n8871);
   U772 : NAND2_X1 port map( A1 => n16396, A2 => n14288, ZN => n16754);
   U773 : OAI21_X1 port map( B1 => n16396, B2 => n14288, A => n16754, ZN => 
                           n17970);
   U774 : NOR3_X1 port map( A1 => n14353, A2 => n16398, A3 => n17970, ZN => 
                           n3027);
   U775 : AOI221_X1 port map( B1 => n14353, B2 => n16398, C1 => n17970, C2 => 
                           n16398, A => n3027, ZN => n8867);
   U776 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n18048);
   U777 : INV_X1 port map( A => n18048, ZN => n18052);
   U778 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN 
                           => n17800);
   U779 : NAND2_X1 port map( A1 => n17800, A2 => data2_mul_1_port, ZN => n18047
                           );
   U780 : INV_X1 port map( A => n18047, ZN => n18050);
   U781 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => n17800, ZN => n18046)
                           ;
   U782 : AOI222_X1 port map( A1 => n18052, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           n18050, B2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C1 => 
                           n18046, C2 => n9081, ZN => n16756);
   U783 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n17836);
   U784 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n17836, ZN => n17803);
   U785 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n17803, ZN => n16755
                           );
   U786 : NOR2_X1 port map( A1 => n16756, A2 => n16755, ZN => n3036);
   U787 : AOI21_X1 port map( B1 => n16756, B2 => n16755, A => n3036, ZN => 
                           n8861);
   U788 : NAND2_X1 port map( A1 => DATA1(9), A2 => n17791, ZN => n17641);
   U789 : NOR2_X1 port map( A1 => DATA1(9), A2 => n17791, ZN => n17587);
   U790 : INV_X1 port map( A => n17587, ZN => n17640);
   U791 : NAND2_X1 port map( A1 => n17641, A2 => n17640, ZN => n16757);
   U792 : AOI22_X1 port map( A1 => n17538, A2 => n14088, B1 => n18171, B2 => 
                           n16757, ZN => n8675);
   U793 : NOR2_X1 port map( A1 => n16758, A2 => n16761, ZN => n17514);
   U794 : NAND2_X1 port map( A1 => n17473, A2 => n17769, ZN => n18163);
   U795 : AOI211_X1 port map( C1 => n16758, C2 => n16761, A => n17514, B => 
                           n18163, ZN => n8674);
   U796 : NAND2_X1 port map( A1 => n14469, A2 => DATA2_I_8_port, ZN => n16760);
   U797 : INV_X1 port map( A => n17523, ZN => n16759);
   U798 : NOR2_X1 port map( A1 => n18230, A2 => n17473, ZN => n17481);
   U799 : INV_X1 port map( A => n17481, ZN => n17508);
   U800 : AOI211_X1 port map( C1 => n16761, C2 => n16760, A => n16759, B => 
                           n17508, ZN => n8673);
   U801 : INV_X1 port map( A => n18162, ZN => n17493);
   U802 : NAND3_X1 port map( A1 => DATA2(9), A2 => DATA1(9), A3 => n17493, ZN 
                           => n8859);
   U803 : INV_X1 port map( A => n16802, ZN => n16762);
   U804 : OAI22_X1 port map( A1 => n16825, A2 => n18150, B1 => n16762, B2 => 
                           n18138, ZN => n16764);
   U805 : OAI22_X1 port map( A1 => n16824, A2 => n18152, B1 => n18137, B2 => 
                           n18154, ZN => n16763);
   U806 : OAI21_X1 port map( B1 => n16764, B2 => n16763, A => n1868, ZN => 
                           n11714);
   U807 : AOI22_X1 port map( A1 => n14383, A2 => n13994, B1 => n14396, B2 => 
                           n14440, ZN => n16766);
   U808 : AOI22_X1 port map( A1 => n14334, A2 => n13985, B1 => n14393, B2 => 
                           n13996, ZN => n16765);
   U809 : OAI211_X1 port map( C1 => n14274, C2 => n14441, A => n16766, B => 
                           n16765, ZN => n17420);
   U810 : INV_X1 port map( A => n17420, ZN => n17427);
   U811 : AOI22_X1 port map( A1 => n14383, A2 => n14445, B1 => n13996, B2 => 
                           n14396, ZN => n16768);
   U812 : AOI22_X1 port map( A1 => n14187, A2 => n13986, B1 => n14393, B2 => 
                           n13994, ZN => n16767);
   U813 : OAI211_X1 port map( C1 => n14349, C2 => n13993, A => n16768, B => 
                           n16767, ZN => n16769);
   U814 : INV_X1 port map( A => n16769, ZN => n17428);
   U815 : OAI22_X1 port map( A1 => n14454, A2 => n14446, B1 => n14391, B2 => 
                           n13993, ZN => n16770);
   U816 : AOI211_X1 port map( C1 => n14333, C2 => n13996, A => n13995, B => 
                           n16770, ZN => n16775);
   U817 : OAI222_X1 port map( A1 => n17427, A2 => n18186, B1 => n17428, B2 => 
                           n18177, C1 => n16775, C2 => n18198, ZN => n17453);
   U818 : INV_X1 port map( A => n17453, ZN => n17488);
   U819 : OAI22_X1 port map( A1 => n14274, A2 => n14446, B1 => n14436, B2 => 
                           n14444, ZN => n16771);
   U820 : AOI211_X1 port map( C1 => n14383, C2 => n14448, A => n13991, B => 
                           n16771, ZN => n16776);
   U821 : OAI222_X1 port map( A1 => n18177, A2 => n16775, B1 => n18198, B2 => 
                           n16776, C1 => n18186, C2 => n17428, ZN => n16791);
   U822 : AOI22_X1 port map( A1 => n14334, A2 => n13994, B1 => n14340, B2 => 
                           n14003, ZN => n16772);
   U823 : INV_X1 port map( A => n16772, ZN => n16773);
   U824 : AOI211_X1 port map( C1 => n14364, C2 => n14445, A => n13992, B => 
                           n16773, ZN => n16779);
   U825 : OAI22_X1 port map( A1 => n14231, A2 => n14447, B1 => n14391, B2 => 
                           n13998, ZN => n16774);
   U826 : AOI211_X1 port map( C1 => n14003, C2 => n14341, A => n13997, B => 
                           n16774, ZN => n16784);
   U827 : OAI222_X1 port map( A1 => n18180, A2 => n16776, B1 => n14228, B2 => 
                           n16779, C1 => n14390, C2 => n16784, ZN => n16792);
   U828 : AOI22_X1 port map( A1 => n18176, A2 => n16791, B1 => n18181, B2 => 
                           n16792, ZN => n16781);
   U829 : OAI22_X1 port map( A1 => n14228, A2 => n16776, B1 => n14373, B2 => 
                           n16775, ZN => n16777);
   U830 : INV_X1 port map( A => n16777, ZN => n16778);
   U831 : OAI21_X1 port map( B1 => n16779, B2 => n14390, A => n16778, ZN => 
                           n16795);
   U832 : OAI211_X1 port map( C1 => n14436, C2 => n14001, A => n14000, B => 
                           n13999, ZN => n16786);
   U833 : INV_X1 port map( A => n16786, ZN => n16785);
   U834 : OAI222_X1 port map( A1 => n18195, A2 => n16785, B1 => n14228, B2 => 
                           n16784, C1 => n16779, C2 => n14373, ZN => n16834);
   U835 : AOI22_X1 port map( A1 => n13893, A2 => n16795, B1 => n18184, B2 => 
                           n16834, ZN => n16780);
   U836 : OAI211_X1 port map( C1 => n14332, C2 => n17488, A => n16781, B => 
                           n16780, ZN => n17524);
   U837 : INV_X1 port map( A => n16834, ZN => n16811);
   U838 : AOI22_X1 port map( A1 => n14383, A2 => n14005, B1 => n14003, B2 => 
                           n14435, ZN => n16783);
   U839 : AOI22_X1 port map( A1 => n14363, A2 => n14002, B1 => n14393, B2 => 
                           n14004, ZN => n16782);
   U840 : OAI211_X1 port map( C1 => n14006, C2 => n14366, A => n16783, B => 
                           n16782, ZN => n16787);
   U841 : INV_X1 port map( A => n16787, ZN => n16810);
   U842 : OAI222_X1 port map( A1 => n16785, A2 => n18177, B1 => n16784, B2 => 
                           n18180, C1 => n16810, C2 => n18195, ZN => n16833);
   U843 : AOI22_X1 port map( A1 => n18176, A2 => n16792, B1 => n16833, B2 => 
                           n14348, ZN => n16790);
   U844 : OAI211_X1 port map( C1 => n14226, C2 => n14443, A => n13990, B => 
                           n13989, ZN => n16809);
   U845 : AOI222_X1 port map( A1 => n16787, A2 => n14420, B1 => n16786, B2 => 
                           n14456, C1 => n16809, C2 => n14188, ZN => n16867);
   U846 : INV_X1 port map( A => n16795, ZN => n17486);
   U847 : OAI22_X1 port map( A1 => n14389, A2 => n16867, B1 => n14350, B2 => 
                           n17486, ZN => n16788);
   U848 : INV_X1 port map( A => n16788, ZN => n16789);
   U849 : OAI211_X1 port map( C1 => n14417, C2 => n16811, A => n16790, B => 
                           n16789, ZN => n16814);
   U850 : INV_X1 port map( A => n16791, ZN => n17487);
   U851 : INV_X1 port map( A => n16833, ZN => n16868);
   U852 : OAI22_X1 port map( A1 => n14332, A2 => n17487, B1 => n14389, B2 => 
                           n16868, ZN => n16794);
   U853 : INV_X1 port map( A => n16792, ZN => n17485);
   U854 : OAI22_X1 port map( A1 => n14134, A2 => n16811, B1 => n14417, B2 => 
                           n17485, ZN => n16793);
   U855 : AOI211_X1 port map( C1 => n14395, C2 => n16795, A => n16794, B => 
                           n16793, ZN => n16837);
   U856 : INV_X1 port map( A => n16837, ZN => n17525);
   U857 : AOI222_X1 port map( A1 => n18178, A2 => n17524, B1 => n16814, B2 => 
                           n18189, C1 => n17525, C2 => n18209, ZN => n16798);
   U858 : NAND2_X1 port map( A1 => n13983, A2 => n14169, ZN => n16796);
   U859 : NOR3_X1 port map( A1 => n13982, A2 => n13981, A3 => n16796, ZN => 
                           n16797);
   U860 : OAI211_X1 port map( C1 => n16798, C2 => n18208, A => n14168, B => 
                           n16797, ZN => OUTALU(9));
   U861 : NOR2_X1 port map( A1 => n18193, A2 => DATA2(8), ZN => n17637);
   U862 : AOI21_X1 port map( B1 => n18193, B2 => DATA2(8), A => n17637, ZN => 
                           n16799);
   U863 : INV_X1 port map( A => n16799, ZN => n17557);
   U864 : AOI22_X1 port map( A1 => n14176, A2 => n17538, B1 => n18171, B2 => 
                           n17557, ZN => n8649);
   U865 : INV_X1 port map( A => DATA2(8), ZN => n17792);
   U866 : NOR3_X1 port map( A1 => n18162, A2 => n17792, A3 => n18193, ZN => 
                           n16805);
   U867 : AOI222_X1 port map( A1 => n16802, A2 => n18159, B1 => n16801, B2 => 
                           n18114, C1 => n16800, C2 => n18118, ZN => n16803);
   U868 : OAI22_X1 port map( A1 => n16806, A2 => n18163, B1 => n16803, B2 => 
                           n16878, ZN => n16804);
   U869 : AOI211_X1 port map( C1 => n17481, C2 => n16806, A => n16805, B => 
                           n16804, ZN => n11729);
   U870 : OAI22_X1 port map( A1 => n14134, A2 => n16867, B1 => n14332, B2 => 
                           n17485, ZN => n16813);
   U871 : OAI22_X1 port map( A1 => n14231, A2 => n13979, B1 => n14226, B2 => 
                           n14442, ZN => n16808);
   U872 : OAI22_X1 port map( A1 => n14454, A2 => n14443, B1 => n14436, B2 => 
                           n14447, ZN => n16807);
   U873 : AOI211_X1 port map( C1 => n14333, C2 => n14004, A => n16808, B => 
                           n16807, ZN => n16860);
   U874 : INV_X1 port map( A => n16809, ZN => n16832);
   U875 : OAI222_X1 port map( A1 => n14367, A2 => n16860, B1 => n16810, B2 => 
                           n18180, C1 => n16832, C2 => n18177, ZN => n16863);
   U876 : INV_X1 port map( A => n16863, ZN => n16890);
   U877 : OAI22_X1 port map( A1 => n14225, A2 => n16811, B1 => n14389, B2 => 
                           n16890, ZN => n16812);
   U878 : AOI211_X1 port map( C1 => n16833, C2 => n13893, A => n16813, B => 
                           n16812, ZN => n16874);
   U879 : INV_X1 port map( A => n16874, ZN => n16891);
   U880 : INV_X1 port map( A => n16814, ZN => n16873);
   U881 : AOI22_X1 port map( A1 => n18217, A2 => n17524, B1 => n18178, B2 => 
                           n17525, ZN => n16815);
   U882 : OAI21_X1 port map( B1 => n14136, B2 => n16873, A => n16815, ZN => 
                           n16816);
   U883 : AOI21_X1 port map( B1 => n18189, B2 => n16891, A => n16816, ZN => 
                           n16817);
   U884 : OAI211_X1 port map( C1 => n16817, C2 => n18208, A => n13980, B => 
                           n13978, ZN => OUTALU(8));
   U885 : OAI221_X1 port map( B1 => n16393, B2 => n17530, C1 => n14467, C2 => 
                           n17521, A => n17424, ZN => n16821);
   U886 : INV_X1 port map( A => n16818, ZN => n16829);
   U887 : OAI21_X1 port map( B1 => n16843, B2 => n16845, A => n16819, ZN => 
                           n16823);
   U888 : OAI21_X1 port map( B1 => n16842, B2 => n16845, A => n16819, ZN => 
                           n16822);
   U889 : OAI22_X1 port map( A1 => n17335, A2 => n16823, B1 => n1866, B2 => 
                           n16822, ZN => n16820);
   U890 : AOI22_X1 port map( A1 => DATA2(7), A2 => n16821, B1 => n16829, B2 => 
                           n16820, ZN => n8646);
   U891 : NAND2_X1 port map( A1 => n1869, A2 => n1904, ZN => n11755);
   U892 : NOR2_X1 port map( A1 => n16393, A2 => DATA2(7), ZN => n17636);
   U893 : AOI22_X1 port map( A1 => n17533, A2 => n16823, B1 => n17537, B2 => 
                           n16822, ZN => n16828);
   U894 : OAI22_X1 port map( A1 => n18137, A2 => n16825, B1 => n16824, B2 => 
                           n18148, ZN => n16826);
   U895 : AOI22_X1 port map( A1 => n17538, A2 => n14095, B1 => n1868, B2 => 
                           n16826, ZN => n16827);
   U896 : OAI21_X1 port map( B1 => n16829, B2 => n16828, A => n16827, ZN => 
                           n16830);
   U897 : AOI21_X1 port map( B1 => n17636, B2 => n18171, A => n16830, ZN => 
                           n11754);
   U898 : OAI22_X1 port map( A1 => n14274, A2 => n14443, B1 => n14454, B2 => 
                           n14442, ZN => n16831);
   U899 : AOI211_X1 port map( C1 => n14004, C2 => n14187, A => n13988, B => 
                           n16831, ZN => n16859);
   U900 : OAI222_X1 port map( A1 => n18180, A2 => n16832, B1 => n18177, B2 => 
                           n16860, C1 => n16859, C2 => n14367, ZN => n16912);
   U901 : AOI22_X1 port map( A1 => n18176, A2 => n16833, B1 => n18184, B2 => 
                           n16912, ZN => n16836);
   U902 : AOI22_X1 port map( A1 => n14221, A2 => n16834, B1 => n18181, B2 => 
                           n16863, ZN => n16835);
   U903 : OAI211_X1 port map( C1 => n16867, C2 => n14345, A => n16836, B => 
                           n16835, ZN => n16915);
   U904 : INV_X1 port map( A => n16915, ZN => n16894);
   U905 : OAI22_X1 port map( A1 => n14136, A2 => n16874, B1 => n16894, B2 => 
                           n18183, ZN => n16839);
   U906 : OAI22_X1 port map( A1 => n14137, A2 => n16837, B1 => n14403, B2 => 
                           n16873, ZN => n16838);
   U907 : AOI211_X1 port map( C1 => n18192, C2 => n17524, A => n16839, B => 
                           n16838, ZN => n18130);
   U908 : OAI211_X1 port map( C1 => n18130, C2 => n14273, A => n13977, B => 
                           n13976, ZN => OUTALU(7));
   U909 : INV_X1 port map( A => DATA2(6), ZN => n17796);
   U910 : NOR2_X1 port map( A1 => n17796, A2 => n18202, ZN => n16840);
   U911 : AOI21_X1 port map( B1 => n17796, B2 => n14466, A => n16840, ZN => 
                           n17635);
   U912 : AOI21_X1 port map( B1 => n17518, B2 => n14466, A => n17517, ZN => 
                           n16841);
   U913 : OAI22_X1 port map( A1 => n17635, A2 => n17521, B1 => n16841, B2 => 
                           n17796, ZN => n8642);
   U914 : OAI22_X1 port map( A1 => n16843, A2 => n17335, B1 => n16842, B2 => 
                           n1866, ZN => n16844);
   U915 : NAND2_X1 port map( A1 => n16845, A2 => n16844, ZN => n8957);
   U916 : OAI21_X1 port map( B1 => n14453, B2 => n17530, A => n17424, ZN => 
                           n16848);
   U917 : OAI22_X1 port map( A1 => n16879, A2 => n17349, B1 => n16846, B2 => 
                           n17318, ZN => n16847);
   U918 : AOI22_X1 port map( A1 => DATA2(5), A2 => n16848, B1 => n1868, B2 => 
                           n16847, ZN => n8640);
   U919 : AOI22_X1 port map( A1 => DATA2(5), A2 => n14465, B1 => n14453, B2 => 
                           n17797, ZN => n17555);
   U920 : AOI22_X1 port map( A1 => n17538, A2 => n14103, B1 => n18171, B2 => 
                           n17555, ZN => n8639);
   U921 : AOI22_X1 port map( A1 => n16851, A2 => n17533, B1 => n16850, B2 => 
                           n17537, ZN => n16849);
   U922 : INV_X1 port map( A => n16849, ZN => n16854);
   U923 : OAI22_X1 port map( A1 => n17335, A2 => n16851, B1 => n1866, B2 => 
                           n16850, ZN => n16853);
   U924 : AOI22_X1 port map( A1 => n16855, A2 => n16854, B1 => n16853, B2 => 
                           n16852, ZN => n8638);
   U925 : AOI22_X1 port map( A1 => n1897, A2 => n1859, B1 => n13151, B2 => 
                           n16856, ZN => n11789);
   U926 : OAI211_X1 port map( C1 => n14226, C2 => n14405, A => n14432, B => 
                           n13971, ZN => n16910);
   U927 : OAI22_X1 port map( A1 => n14274, A2 => n14442, B1 => n14436, B2 => 
                           n14443, ZN => n16857);
   U928 : AOI211_X1 port map( C1 => n14383, C2 => n13890, A => n13987, B => 
                           n16857, ZN => n16887);
   U929 : OAI22_X1 port map( A1 => n16859, A2 => n18180, B1 => n16887, B2 => 
                           n18177, ZN => n16858);
   U930 : AOI21_X1 port map( B1 => n14188, B2 => n16910, A => n16858, ZN => 
                           n17165);
   U931 : INV_X1 port map( A => n17165, ZN => n17362);
   U932 : AOI22_X1 port map( A1 => n18197, A2 => n16912, B1 => n18184, B2 => 
                           n17362, ZN => n16865);
   U933 : OAI22_X1 port map( A1 => n16860, A2 => n18180, B1 => n16859, B2 => 
                           n18177, ZN => n16861);
   U934 : INV_X1 port map( A => n16861, ZN => n16862);
   U935 : OAI21_X1 port map( B1 => n18195, B2 => n16887, A => n16862, ZN => 
                           n17162);
   U936 : AOI22_X1 port map( A1 => n18176, A2 => n16863, B1 => n18181, B2 => 
                           n17162, ZN => n16864);
   U937 : OAI211_X1 port map( C1 => n16867, C2 => n18200, A => n16865, B => 
                           n16864, ZN => n17166);
   U938 : INV_X1 port map( A => n17166, ZN => n17368);
   U939 : OAI22_X1 port map( A1 => n14137, A2 => n16874, B1 => n17368, B2 => 
                           n18183, ZN => n16872);
   U940 : INV_X1 port map( A => n17162, ZN => n16866);
   U941 : OAI22_X1 port map( A1 => n14225, A2 => n16867, B1 => n16866, B2 => 
                           n18196, ZN => n16870);
   U942 : OAI22_X1 port map( A1 => n16868, A2 => n18200, B1 => n16890, B2 => 
                           n18182, ZN => n16869);
   U943 : AOI211_X1 port map( C1 => n14348, C2 => n16912, A => n16870, B => 
                           n16869, ZN => n17169);
   U944 : OAI22_X1 port map( A1 => n14136, A2 => n17169, B1 => n14458, B2 => 
                           n16873, ZN => n16871);
   U945 : AOI211_X1 port map( C1 => n13894, C2 => n16915, A => n16872, B => 
                           n16871, ZN => n16908);
   U946 : OAI22_X1 port map( A1 => n14136, A2 => n16894, B1 => n16873, B2 => 
                           n18203, ZN => n16876);
   U947 : OAI22_X1 port map( A1 => n14401, A2 => n17169, B1 => n14403, B2 => 
                           n16874, ZN => n16875);
   U948 : AOI211_X1 port map( C1 => n18192, C2 => n17525, A => n16876, B => 
                           n16875, ZN => n18131);
   U949 : OAI222_X1 port map( A1 => n14133, A2 => n16908, B1 => n14330, B2 => 
                           n18130, C1 => n14382, C2 => n18131, ZN => n17374);
   U950 : NAND3_X1 port map( A1 => n18190, A2 => n17374, A3 => n18179, ZN => 
                           n16877);
   U951 : NAND4_X1 port map( A1 => n13973, A2 => n13972, A3 => n13974, A4 => 
                           n16877, ZN => OUTALU(5));
   U952 : AOI22_X1 port map( A1 => n17533, A2 => n16885, B1 => n17537, B2 => 
                           n16884, ZN => n8636);
   U953 : NOR3_X1 port map( A1 => n16879, A2 => n16878, A3 => n17318, ZN => 
                           n16883);
   U954 : INV_X1 port map( A => DATA2(4), ZN => n18058);
   U955 : NAND2_X1 port map( A1 => n18058, A2 => n14464, ZN => n17629);
   U956 : NAND2_X1 port map( A1 => DATA2(4), A2 => n14438, ZN => n17633);
   U957 : NAND2_X1 port map( A1 => n17629, A2 => n17633, ZN => n17549);
   U958 : INV_X1 port map( A => n17549, ZN => n16881);
   U959 : AOI21_X1 port map( B1 => n17518, B2 => n14464, A => n17517, ZN => 
                           n16880);
   U960 : OAI22_X1 port map( A1 => n16881, A2 => n17521, B1 => n16880, B2 => 
                           n18058, ZN => n16882);
   U961 : AOI211_X1 port map( C1 => n17538, C2 => n13884, A => n16883, B => 
                           n16882, ZN => n8635);
   U962 : OAI22_X1 port map( A1 => n16885, A2 => n17335, B1 => n16884, B2 => 
                           n1866, ZN => n8634);
   U963 : AOI22_X1 port map( A1 => n1897, A2 => n1862, B1 => n1894, B2 => n1865
                           , ZN => n11811);
   U964 : OAI211_X1 port map( C1 => n14454, C2 => n14405, A => n13967, B => 
                           n14431, ZN => n17159);
   U965 : AOI22_X1 port map( A1 => n14420, A2 => n16910, B1 => n14188, B2 => 
                           n17159, ZN => n16886);
   U966 : OAI21_X1 port map( B1 => n16887, B2 => n18180, A => n16886, ZN => 
                           n17739);
   U967 : AOI22_X1 port map( A1 => n18205, A2 => n17739, B1 => n18181, B2 => 
                           n17362, ZN => n16889);
   U968 : AOI22_X1 port map( A1 => n13893, A2 => n17162, B1 => n18176, B2 => 
                           n16912, ZN => n16888);
   U969 : OAI211_X1 port map( C1 => n14332, C2 => n16890, A => n16889, B => 
                           n16888, ZN => n17748);
   U970 : INV_X1 port map( A => n17169, ZN => n16916);
   U971 : AOI22_X1 port map( A1 => n14129, A2 => n17748, B1 => n18178, B2 => 
                           n16916, ZN => n16893);
   U972 : AOI22_X1 port map( A1 => n14387, A2 => n17166, B1 => n18192, B2 => 
                           n16891, ZN => n16892);
   U973 : OAI211_X1 port map( C1 => n14137, C2 => n16894, A => n16893, B => 
                           n16892, ZN => n17170);
   U974 : INV_X1 port map( A => n17170, ZN => n16895);
   U975 : OAI222_X1 port map( A1 => n14133, A2 => n16895, B1 => n14330, B2 => 
                           n18131, C1 => n14382, C2 => n16908, ZN => n17758);
   U976 : INV_X1 port map( A => n17758, ZN => n17157);
   U977 : INV_X1 port map( A => n17374, ZN => n17158);
   U978 : OAI22_X1 port map( A1 => n14400, A2 => n17157, B1 => n14397, B2 => 
                           n17158, ZN => n16896);
   U979 : AOI22_X1 port map( A1 => n14386, A2 => n16896, B1 => n13968, B2 => 
                           n14185, ZN => n16897);
   U980 : OAI211_X1 port map( C1 => n14185, C2 => n13970, A => n13969, B => 
                           n16897, ZN => OUTALU(4));
   U981 : NAND2_X1 port map( A1 => n14326, A2 => n18082, ZN => n17628);
   U982 : NAND2_X1 port map( A1 => DATA2(3), A2 => n14449, ZN => n17627);
   U983 : NAND2_X1 port map( A1 => n17628, A2 => n17627, ZN => n17560);
   U984 : AOI22_X1 port map( A1 => n17279, A2 => n14461, B1 => n17144, B2 => 
                           n18194, ZN => n16899);
   U985 : NAND2_X1 port map( A1 => n14326, A2 => n17345, ZN => n16898);
   U986 : OAI211_X1 port map( C1 => n14451, C2 => n17348, A => n16899, B => 
                           n16898, ZN => n16900);
   U987 : AOI22_X1 port map( A1 => n18171, A2 => n17560, B1 => n1868, B2 => 
                           n16900, ZN => n8632);
   U988 : OAI21_X1 port map( B1 => n14449, B2 => n17530, A => n17424, ZN => 
                           n16901);
   U989 : AOI22_X1 port map( A1 => DATA2(3), A2 => n16901, B1 => n17538, B2 => 
                           n14123, ZN => n8631);
   U990 : AOI21_X1 port map( B1 => n18056, B2 => n16903, A => n16902, ZN => 
                           n16904);
   U991 : NAND2_X1 port map( A1 => n17533, A2 => n16904, ZN => n8956);
   U992 : INV_X1 port map( A => n1859, ZN => n17358);
   U993 : OAI22_X1 port map( A1 => n17355, A2 => n18150, B1 => n18136, B2 => 
                           n18152, ZN => n16907);
   U994 : INV_X1 port map( A => n16905, ZN => n18139);
   U995 : INV_X1 port map( A => n17723, ZN => n17354);
   U996 : OAI22_X1 port map( A1 => n18155, A2 => n18139, B1 => n17354, B2 => 
                           n18138, ZN => n16906);
   U997 : AOI211_X1 port map( C1 => n18159, C2 => n17724, A => n16907, B => 
                           n16906, ZN => n17731);
   U998 : OAI22_X1 port map( A1 => n17358, A2 => n1896, B1 => n17731, B2 => 
                           n17499, ZN => n11849);
   U999 : INV_X1 port map( A => n16908, ZN => n16919);
   U1000 : INV_X1 port map( A => n17748, ZN => n17367);
   U1001 : OAI22_X1 port map( A1 => n14274, A2 => n14405, B1 => n14226, B2 => 
                           n13892, ZN => n16909);
   U1002 : AOI211_X1 port map( C1 => n14187, C2 => n14404, A => n13964, B => 
                           n16909, ZN => n17361);
   U1003 : AOI22_X1 port map( A1 => n14420, A2 => n17159, B1 => n14456, B2 => 
                           n16910, ZN => n16911);
   U1004 : OAI21_X1 port map( B1 => n17361, B2 => n18195, A => n16911, ZN => 
                           n17738);
   U1005 : AOI22_X1 port map( A1 => n14130, A2 => n17738, B1 => n14384, B2 => 
                           n17739, ZN => n16914);
   U1006 : AOI22_X1 port map( A1 => n14220, A2 => n16912, B1 => n14395, B2 => 
                           n17162, ZN => n16913);
   U1007 : OAI211_X1 port map( C1 => n14417, C2 => n17165, A => n16914, B => 
                           n16913, ZN => n17736);
   U1008 : AOI22_X1 port map( A1 => n14129, A2 => n17736, B1 => n13894, B2 => 
                           n17166, ZN => n16918);
   U1009 : AOI22_X1 port map( A1 => n14398, A2 => n16916, B1 => n14375, B2 => 
                           n16915, ZN => n16917);
   U1010 : OAI211_X1 port map( C1 => n14136, C2 => n17367, A => n16918, B => 
                           n16917, ZN => n17371);
   U1011 : AOI222_X1 port map( A1 => n14139, A2 => n17170, B1 => n14229, B2 => 
                           n16919, C1 => n14381, C2 => n17371, ZN => n17373);
   U1012 : OAI222_X1 port map( A1 => n14400, A2 => n17373, B1 => n14232, B2 => 
                           n17158, C1 => n14397, C2 => n17157, ZN => n16920);
   U1013 : AOI22_X1 port map( A1 => n14386, A2 => n16920, B1 => n14140, B2 => 
                           n14277, ZN => n16921);
   U1014 : NAND4_X1 port map( A1 => n13966, A2 => n13965, A3 => n14271, A4 => 
                           n16921, ZN => OUTALU(3));
   U1015 : NOR2_X1 port map( A1 => n17264, A2 => n17655, ZN => n16925);
   U1016 : OR4_X1 port map( A1 => n16925, A2 => n16924, A3 => n16923, A4 => 
                           n16922, ZN => n16926);
   U1017 : AOI21_X1 port map( B1 => DATA1(17), B2 => n17339, A => n16926, ZN =>
                           n16927);
   U1018 : INV_X1 port map( A => n16927, ZN => n16943);
   U1019 : AOI222_X1 port map( A1 => n17352, A2 => n16928, B1 => n16942, B2 => 
                           n16944, C1 => n16945, C2 => n16943, ZN => n16929);
   U1020 : INV_X1 port map( A => n16929, ZN => n18106);
   U1021 : AOI22_X1 port map( A1 => n18159, A2 => n16991, B1 => n18123, B2 => 
                           n18106, ZN => n16931);
   U1022 : AOI22_X1 port map( A1 => n18118, A2 => n18102, B1 => n18116, B2 => 
                           n18101, ZN => n16930);
   U1023 : OAI211_X1 port map( C1 => n18099, C2 => n18152, A => n16931, B => 
                           n16930, ZN => n11966);
   U1024 : INV_X1 port map( A => n1879, ZN => n16934);
   U1025 : AOI22_X1 port map( A1 => n1894, A2 => n11966, B1 => n11927, B2 => 
                           n16934, ZN => n11952);
   U1026 : AOI22_X1 port map( A1 => n1898, A2 => n16934, B1 => n11927, B2 => 
                           n11966, ZN => n11955);
   U1027 : AOI22_X1 port map( A1 => n18116, A2 => n16991, B1 => n18159, B2 => 
                           n16957, ZN => n16933);
   U1028 : AOI22_X1 port map( A1 => n18144, A2 => n18102, B1 => n18123, B2 => 
                           n18101, ZN => n16932);
   U1029 : OAI211_X1 port map( C1 => n16956, C2 => n18148, A => n16933, B => 
                           n16932, ZN => n1878);
   U1030 : AOI22_X1 port map( A1 => n1894, A2 => n16934, B1 => n11927, B2 => 
                           n1878, ZN => n11960);
   U1031 : INV_X1 port map( A => n1873, ZN => n16995);
   U1032 : AOI22_X1 port map( A1 => n1897, A2 => n16995, B1 => n13151, B2 => 
                           n11966, ZN => n11959);
   U1033 : NAND2_X1 port map( A1 => DATA1(13), A2 => n16978, ZN => n16936);
   U1034 : OAI211_X1 port map( C1 => n17192, C2 => n17655, A => n16936, B => 
                           n16935, ZN => n16937);
   U1035 : OR3_X1 port map( A1 => n16939, A2 => n16938, A3 => n16937, ZN => 
                           n16946);
   U1036 : AOI222_X1 port map( A1 => n17352, A2 => n16943, B1 => n16942, B2 => 
                           n16946, C1 => n16945, C2 => n16940, ZN => n18095);
   U1037 : OAI22_X1 port map( A1 => n18137, A2 => n18099, B1 => n18095, B2 => 
                           n18152, ZN => n16948);
   U1038 : AOI222_X1 port map( A1 => n16941, A2 => n16945, B1 => n16946, B2 => 
                           n17352, C1 => n16940, C2 => n16942, ZN => n16966);
   U1039 : AOI222_X1 port map( A1 => n16946, A2 => n16945, B1 => n16944, B2 => 
                           n17352, C1 => n16943, C2 => n16942, ZN => n18100);
   U1040 : OAI22_X1 port map( A1 => n18155, A2 => n16966, B1 => n18100, B2 => 
                           n18150, ZN => n16947);
   U1041 : AOI211_X1 port map( C1 => n18118, C2 => n18106, A => n16948, B => 
                           n16947, ZN => n11979);
   U1042 : INV_X1 port map( A => n18095, ZN => n18092);
   U1043 : OAI22_X1 port map( A1 => n18155, A2 => n16967, B1 => n16969, B2 => 
                           n18150, ZN => n16950);
   U1044 : OAI22_X1 port map( A1 => n16966, A2 => n18148, B1 => n16970, B2 => 
                           n18152, ZN => n16949);
   U1045 : AOI211_X1 port map( C1 => n18159, C2 => n18092, A => n16950, B => 
                           n16949, ZN => n8612);
   U1046 : OAI22_X1 port map( A1 => n16966, A2 => n18150, B1 => n16969, B2 => 
                           n18152, ZN => n16952);
   U1047 : OAI22_X1 port map( A1 => n18137, A2 => n18100, B1 => n18155, B2 => 
                           n16970, ZN => n16951);
   U1048 : AOI211_X1 port map( C1 => n18118, C2 => n18092, A => n16952, B => 
                           n16951, ZN => n13186);
   U1049 : OAI22_X1 port map( A1 => n8612, A2 => n9020, B1 => n13186, B2 => 
                           n1896, ZN => n11981);
   U1050 : NOR2_X1 port map( A1 => n17695, A2 => n17348, ZN => n17203);
   U1051 : NAND2_X1 port map( A1 => DATA1(27), A2 => n17144, ZN => n17246);
   U1052 : NAND2_X1 port map( A1 => DATA1(25), A2 => n16978, ZN => n16953);
   U1053 : OAI211_X1 port map( C1 => n17192, C2 => n17689, A => n17246, B => 
                           n16953, ZN => n16954);
   U1054 : AOI211_X1 port map( C1 => n17713, C2 => DATA1(29), A => n17203, B =>
                           n16954, ZN => n16981);
   U1055 : OAI222_X1 port map( A1 => n17720, A2 => n16981, B1 => n17718, B2 => 
                           n16963, C1 => n17315, C2 => n16955, ZN => n16988);
   U1056 : AOI22_X1 port map( A1 => n18116, A2 => n16989, B1 => n18159, B2 => 
                           n16988, ZN => n16959);
   U1057 : INV_X1 port map( A => n16956, ZN => n16990);
   U1058 : AOI22_X1 port map( A1 => n18144, A2 => n16957, B1 => n18123, B2 => 
                           n16990, ZN => n16958);
   U1059 : OAI211_X1 port map( C1 => n16960, C2 => n18148, A => n16959, B => 
                           n16958, ZN => n16996);
   U1060 : AOI22_X1 port map( A1 => n1898, A2 => n16995, B1 => n1897, B2 => 
                           n16996, ZN => n11996);
   U1061 : INV_X1 port map( A => DATA1(29), ZN => n17247);
   U1062 : NOR2_X1 port map( A1 => n17247, A2 => n17348, ZN => n17194);
   U1063 : NAND2_X1 port map( A1 => DATA1(28), A2 => n17144, ZN => n17226);
   U1064 : NAND2_X1 port map( A1 => DATA1(27), A2 => n17279, ZN => n16961);
   U1065 : OAI211_X1 port map( C1 => n17264, C2 => n17689, A => n17226, B => 
                           n16961, ZN => n16962);
   U1066 : AOI211_X1 port map( C1 => n17713, C2 => DATA1(30), A => n17194, B =>
                           n16962, ZN => n16982);
   U1067 : OAI222_X1 port map( A1 => n17720, A2 => n16982, B1 => n17718, B2 => 
                           n16981, C1 => n17315, C2 => n16963, ZN => n16977);
   U1068 : AOI22_X1 port map( A1 => n18116, A2 => n16976, B1 => n18159, B2 => 
                           n16977, ZN => n16965);
   U1069 : AOI22_X1 port map( A1 => n18118, A2 => n16988, B1 => n18144, B2 => 
                           n16989, ZN => n16964);
   U1070 : OAI211_X1 port map( C1 => n18155, C2 => n16994, A => n16965, B => 
                           n16964, ZN => n16997);
   U1071 : AOI22_X1 port map( A1 => n1898, A2 => n16996, B1 => n1897, B2 => 
                           n16997, ZN => n12004);
   U1072 : INV_X1 port map( A => n16966, ZN => n18091);
   U1073 : OAI22_X1 port map( A1 => n18155, A2 => n16968, B1 => n16967, B2 => 
                           n18152, ZN => n16972);
   U1074 : OAI22_X1 port map( A1 => n16970, A2 => n18150, B1 => n16969, B2 => 
                           n18138, ZN => n16971);
   U1075 : AOI211_X1 port map( C1 => n18159, C2 => n18091, A => n16972, B => 
                           n16971, ZN => n1855);
   U1076 : INV_X1 port map( A => n1852, ZN => n16973);
   U1077 : OAI22_X1 port map( A1 => n1855, A2 => n17728, B1 => n16973, B2 => 
                           n9020, ZN => n12032);
   U1078 : INV_X1 port map( A => n1854, ZN => n16974);
   U1079 : OAI22_X1 port map( A1 => n8612, A2 => n17499, B1 => n16974, B2 => 
                           n1896, ZN => n12031);
   U1080 : OAI22_X1 port map( A1 => n16973, A2 => n1896, B1 => n16974, B2 => 
                           n17728, ZN => n12042);
   U1081 : INV_X1 port map( A => n1857, ZN => n17484);
   U1082 : OAI22_X1 port map( A1 => n17484, A2 => n1895, B1 => n16974, B2 => 
                           n17499, ZN => n12045);
   U1083 : INV_X1 port map( A => n1853, ZN => n16975);
   U1084 : OAI22_X1 port map( A1 => n8604, A2 => n1895, B1 => n16975, B2 => 
                           n17728, ZN => n12047);
   U1085 : AOI22_X1 port map( A1 => n18118, A2 => n16977, B1 => n18144, B2 => 
                           n16976, ZN => n16986);
   U1086 : NOR2_X1 port map( A1 => n17247, A2 => n17276, ZN => n17202);
   U1087 : INV_X1 port map( A => DATA1(30), ZN => n17702);
   U1088 : NAND2_X1 port map( A1 => DATA1(28), A2 => n17279, ZN => n16979);
   U1089 : NAND2_X1 port map( A1 => DATA1(27), A2 => n16978, ZN => n17273);
   U1090 : OAI211_X1 port map( C1 => n17348, C2 => n17702, A => n16979, B => 
                           n17273, ZN => n16980);
   U1091 : AOI211_X1 port map( C1 => n17713, C2 => DATA1(31), A => n17202, B =>
                           n16980, ZN => n16983);
   U1092 : OAI222_X1 port map( A1 => n17720, A2 => n16983, B1 => n17718, B2 => 
                           n16982, C1 => n17315, C2 => n16981, ZN => n16984);
   U1093 : AOI22_X1 port map( A1 => n18159, A2 => n16984, B1 => n18123, B2 => 
                           n16989, ZN => n16985);
   U1094 : NAND2_X1 port map( A1 => n16986, A2 => n16985, ZN => n16987);
   U1095 : AOI21_X1 port map( B1 => n18116, B2 => n16988, A => n16987, ZN => 
                           n12088);
   U1096 : AOI22_X1 port map( A1 => n18116, A2 => n16990, B1 => n18159, B2 => 
                           n16989, ZN => n16993);
   U1097 : AOI22_X1 port map( A1 => n18144, A2 => n16991, B1 => n18123, B2 => 
                           n18102, ZN => n16992);
   U1098 : OAI211_X1 port map( C1 => n16994, C2 => n18148, A => n16993, B => 
                           n16992, ZN => n1875);
   U1099 : AOI22_X1 port map( A1 => n13151, A2 => n1875, B1 => n1894, B2 => 
                           n16995, ZN => n12087);
   U1100 : AOI22_X1 port map( A1 => n1898, A2 => n16997, B1 => n11927, B2 => 
                           n16996, ZN => n12086);
   U1101 : INV_X1 port map( A => n17260, ZN => n17180);
   U1102 : OAI22_X1 port map( A1 => n16999, A2 => n17182, B1 => n16998, B2 => 
                           n17180, ZN => n17183);
   U1103 : AOI22_X1 port map( A1 => n17769, A2 => n11946, B1 => n17137, B2 => 
                           n17183, ZN => n1808);
   U1104 : INV_X1 port map( A => DATA2(31), ZN => n17770);
   U1105 : INV_X1 port map( A => n1869, ZN => n17292);
   U1106 : OAI22_X1 port map( A1 => n17770, A2 => n17530, B1 => n17000, B2 => 
                           n17292, ZN => n17010);
   U1107 : NAND2_X1 port map( A1 => DATA1(31), A2 => n17770, ZN => n17707);
   U1108 : INV_X1 port map( A => DATA1(31), ZN => n17206);
   U1109 : NAND2_X1 port map( A1 => DATA2(31), A2 => n17206, ZN => n17621);
   U1110 : NAND2_X1 port map( A1 => n17707, A2 => n17621, ZN => n17561);
   U1111 : AOI22_X1 port map( A1 => n6095, A2 => n14009, B1 => n18171, B2 => 
                           n17561, ZN => n17001);
   U1112 : OAI21_X1 port map( B1 => n17770, B2 => n17424, A => n17001, ZN => 
                           n17009);
   U1113 : XNOR2_X1 port map( A => n4293, B => n17206, ZN => n17005);
   U1114 : NAND2_X1 port map( A1 => n17002, A2 => n17005, ZN => n17007);
   U1115 : OAI21_X1 port map( B1 => n11946, B2 => n17137, A => n17002, ZN => 
                           n17004);
   U1116 : INV_X1 port map( A => n11946, ZN => n17138);
   U1117 : INV_X1 port map( A => n12162, ZN => n17003);
   U1118 : AOI22_X1 port map( A1 => n17769, A2 => n17004, B1 => n17138, B2 => 
                           n17003, ZN => n17006);
   U1119 : OAI22_X1 port map( A1 => n1808, A2 => n17007, B1 => n17006, B2 => 
                           n17005, ZN => n17008);
   U1120 : AOI211_X1 port map( C1 => DATA1(31), C2 => n17010, A => n17009, B =>
                           n17008, ZN => n12151);
   U1121 : INV_X1 port map( A => n17055, ZN => n17054);
   U1122 : OAI22_X1 port map( A1 => n14231, A2 => n14407, B1 => n14226, B2 => 
                           n13952, ZN => n17012);
   U1123 : OAI22_X1 port map( A1 => n13963, A2 => n14391, B1 => n14274, B2 => 
                           n18188, ZN => n17011);
   U1124 : AOI211_X1 port map( C1 => n14344, C2 => n14427, A => n17012, B => 
                           n17011, ZN => n17022);
   U1125 : OAI222_X1 port map( A1 => n18228, A2 => n17024, B1 => n14455, B2 => 
                           n17022, C1 => n14374, C2 => n17013, ZN => n17056);
   U1126 : AOI22_X1 port map( A1 => n18185, A2 => n18201, B1 => n13957, B2 => 
                           n14340, ZN => n17016);
   U1127 : OAI22_X1 port map( A1 => n14274, A2 => n13952, B1 => n13951, B2 => 
                           n14436, ZN => n17014);
   U1128 : INV_X1 port map( A => n17014, ZN => n17015);
   U1129 : OAI211_X1 port map( C1 => n14454, C2 => n14407, A => n17016, B => 
                           n17015, ZN => n17032);
   U1130 : INV_X1 port map( A => n17032, ZN => n17021);
   U1131 : OAI22_X1 port map( A1 => n14231, A2 => n14428, B1 => n14407, B2 => 
                           n14376, ZN => n17018);
   U1132 : OAI22_X1 port map( A1 => n14454, A2 => n14408, B1 => n13952, B2 => 
                           n14391, ZN => n17017);
   U1133 : AOI211_X1 port map( C1 => n13957, C2 => n14341, A => n17018, B => 
                           n17017, ZN => n17027);
   U1134 : OAI22_X1 port map( A1 => n14454, A2 => n13952, B1 => n18188, B2 => 
                           n18204, ZN => n17020);
   U1135 : OAI22_X1 port map( A1 => n14274, A2 => n13951, B1 => n14226, B2 => 
                           n14407, ZN => n17019);
   U1136 : AOI211_X1 port map( C1 => n18187, C2 => n18201, A => n17020, B => 
                           n17019, ZN => n17023);
   U1137 : OAI222_X1 port map( A1 => n14228, A2 => n17021, B1 => n14455, B2 => 
                           n17027, C1 => n14374, C2 => n17023, ZN => n17037);
   U1138 : AOI22_X1 port map( A1 => n18176, A2 => n17056, B1 => n17037, B2 => 
                           n18211, ZN => n17026);
   U1139 : OAI222_X1 port map( A1 => n14228, A2 => n17023, B1 => n14455, B2 => 
                           n17021, C1 => n14374, C2 => n17022, ZN => n17047);
   U1140 : OAI222_X1 port map( A1 => n18186, A2 => n17024, B1 => n14455, B2 => 
                           n17023, C1 => n17022, C2 => n14228, ZN => n17050);
   U1141 : AOI22_X1 port map( A1 => n14348, A2 => n17047, B1 => n17050, B2 => 
                           n18197, ZN => n17025);
   U1142 : OAI211_X1 port map( C1 => n17054, C2 => n14360, A => n17026, B => 
                           n17025, ZN => n17110);
   U1143 : INV_X1 port map( A => n17027, ZN => n17033);
   U1144 : OAI22_X1 port map( A1 => n14407, A2 => n14436, B1 => n14408, B2 => 
                           n14349, ZN => n17028);
   U1145 : INV_X1 port map( A => n17028, ZN => n17029);
   U1146 : OAI211_X1 port map( C1 => n14231, C2 => n14166, A => n13955, B => 
                           n17029, ZN => n17034);
   U1147 : OAI22_X1 port map( A1 => n14231, A2 => n13959, B1 => n14436, B2 => 
                           n14408, ZN => n17030);
   U1148 : INV_X1 port map( A => n17030, ZN => n17031);
   U1149 : OAI211_X1 port map( C1 => n14226, C2 => n14166, A => n13956, B => 
                           n17031, ZN => n17071);
   U1150 : AOI222_X1 port map( A1 => n17033, A2 => n14457, B1 => n17034, B2 => 
                           n14420, C1 => n17071, C2 => n14357, ZN => n17067);
   U1151 : OAI211_X1 port map( C1 => n14226, C2 => n13959, A => n13954, B => 
                           n13953, ZN => n17079);
   U1152 : AOI222_X1 port map( A1 => n17034, A2 => n14457, B1 => n17079, B2 => 
                           n14331, C1 => n17071, C2 => n14420, ZN => n17092);
   U1153 : OAI22_X1 port map( A1 => n14134, A2 => n17067, B1 => n17092, B2 => 
                           n18196, ZN => n17036);
   U1154 : INV_X1 port map( A => n17047, ZN => n17040);
   U1155 : AOI222_X1 port map( A1 => n17034, A2 => n14357, B1 => n17033, B2 => 
                           n14358, C1 => n17032, C2 => n14457, ZN => n17080);
   U1156 : OAI22_X1 port map( A1 => n17040, A2 => n14360, B1 => n17080, B2 => 
                           n14417, ZN => n17035);
   U1157 : AOI211_X1 port map( C1 => n18176, C2 => n17037, A => n17036, B => 
                           n17035, ZN => n17100);
   U1158 : INV_X1 port map( A => n17037, ZN => n17072);
   U1159 : OAI22_X1 port map( A1 => n14417, A2 => n17072, B1 => n14389, B2 => 
                           n17067, ZN => n17039);
   U1160 : INV_X1 port map( A => n17050, ZN => n17043);
   U1161 : OAI22_X1 port map( A1 => n14134, A2 => n17080, B1 => n17043, B2 => 
                           n14360, ZN => n17038);
   U1162 : AOI211_X1 port map( C1 => n14347, C2 => n17047, A => n17039, B => 
                           n17038, ZN => n17086);
   U1163 : OAI22_X1 port map( A1 => n14401, A2 => n17100, B1 => n17086, B2 => 
                           n14135, ZN => n17049);
   U1164 : OAI22_X1 port map( A1 => n14134, A2 => n17043, B1 => n14332, B2 => 
                           n17059, ZN => n17042);
   U1165 : OAI22_X1 port map( A1 => n14225, A2 => n17054, B1 => n14361, B2 => 
                           n17040, ZN => n17041);
   U1166 : AOI211_X1 port map( C1 => n13893, C2 => n17056, A => n17042, B => 
                           n17041, ZN => n17123);
   U1167 : OAI22_X1 port map( A1 => n14225, A2 => n17043, B1 => n17080, B2 => 
                           n14389, ZN => n17046);
   U1168 : INV_X1 port map( A => n17056, ZN => n17044);
   U1169 : OAI22_X1 port map( A1 => n17044, A2 => n14360, B1 => n14134, B2 => 
                           n17072, ZN => n17045);
   U1170 : AOI211_X1 port map( C1 => n13893, C2 => n17047, A => n17046, B => 
                           n17045, ZN => n17060);
   U1171 : OAI22_X1 port map( A1 => n17123, A2 => n14458, B1 => n17060, B2 => 
                           n14403, ZN => n17048);
   U1172 : AOI211_X1 port map( C1 => n14342, C2 => n17110, A => n17049, B => 
                           n17048, ZN => n17107);
   U1173 : AOI22_X1 port map( A1 => n17050, A2 => n18184, B1 => n17385, B2 => 
                           n14220, ZN => n17053);
   U1174 : AOI22_X1 port map( A1 => n18176, A2 => n17051, B1 => n17056, B2 => 
                           n18181, ZN => n17052);
   U1175 : OAI211_X1 port map( C1 => n18182, C2 => n17054, A => n17053, B => 
                           n17052, ZN => n17111);
   U1176 : INV_X1 port map( A => n17111, ZN => n17294);
   U1177 : AOI22_X1 port map( A1 => n14220, A2 => n17403, B1 => n18176, B2 => 
                           n17385, ZN => n17058);
   U1178 : AOI22_X1 port map( A1 => n14130, A2 => n17056, B1 => n14348, B2 => 
                           n17055, ZN => n17057);
   U1179 : OAI211_X1 port map( C1 => n17059, C2 => n18182, A => n17058, B => 
                           n17057, ZN => n17122);
   U1180 : INV_X1 port map( A => n17123, ZN => n17063);
   U1181 : AOI22_X1 port map( A1 => n14375, A2 => n17122, B1 => n13894, B2 => 
                           n17063, ZN => n17062);
   U1182 : INV_X1 port map( A => n17060, ZN => n17085);
   U1183 : AOI22_X1 port map( A1 => n14129, A2 => n17085, B1 => n14387, B2 => 
                           n17110, ZN => n17061);
   U1184 : OAI211_X1 port map( C1 => n17294, C2 => n14137, A => n17062, B => 
                           n17061, ZN => n17119);
   U1185 : AOI22_X1 port map( A1 => n14343, A2 => n17085, B1 => n14375, B2 => 
                           n17111, ZN => n17065);
   U1186 : AOI22_X1 port map( A1 => n14398, A2 => n17063, B1 => n13895, B2 => 
                           n17110, ZN => n17064);
   U1187 : OAI211_X1 port map( C1 => n14401, C2 => n17086, A => n17065, B => 
                           n17064, ZN => n17115);
   U1188 : AOI22_X1 port map( A1 => n14229, A2 => n17119, B1 => n14139, B2 => 
                           n17115, ZN => n17066);
   U1189 : OAI21_X1 port map( B1 => n17107, B2 => n18224, A => n17066, ZN => 
                           n17198);
   U1190 : INV_X1 port map( A => n17067, ZN => n17096);
   U1191 : AOI22_X1 port map( A1 => n14187, A2 => n13958, B1 => n14333, B2 => 
                           n14429, ZN => n17068);
   U1192 : OAI211_X1 port map( C1 => n14454, C2 => n13959, A => n13949, B => 
                           n17068, ZN => n17087);
   U1193 : AOI22_X1 port map( A1 => n14420, A2 => n17079, B1 => n14331, B2 => 
                           n17087, ZN => n17069);
   U1194 : INV_X1 port map( A => n17069, ZN => n17070);
   U1195 : AOI21_X1 port map( B1 => n17071, B2 => n14457, A => n17070, ZN => 
                           n17091);
   U1196 : OAI22_X1 port map( A1 => n14134, A2 => n17092, B1 => n14389, B2 => 
                           n17091, ZN => n17074);
   U1197 : OAI22_X1 port map( A1 => n18218, A2 => n17072, B1 => n14225, B2 => 
                           n17080, ZN => n17073);
   U1198 : AOI211_X1 port map( C1 => n18197, C2 => n17096, A => n17074, B => 
                           n17073, ZN => n17098);
   U1199 : OAI22_X1 port map( A1 => n18227, A2 => n17100, B1 => n18183, B2 => 
                           n17098, ZN => n17075);
   U1200 : INV_X1 port map( A => n17075, ZN => n17077);
   U1201 : AOI22_X1 port map( A1 => n14398, A2 => n17085, B1 => n14359, B2 => 
                           n17110, ZN => n17076);
   U1202 : OAI211_X1 port map( C1 => n17086, C2 => n14402, A => n17077, B => 
                           n17076, ZN => n17116);
   U1203 : OAI22_X1 port map( A1 => n14135, A2 => n17098, B1 => n17100, B2 => 
                           n18221, ZN => n17084);
   U1204 : AOI22_X1 port map( A1 => n14334, A2 => n14429, B1 => n14333, B2 => 
                           n14425, ZN => n17078);
   U1205 : OAI211_X1 port map( C1 => n14454, C2 => n14426, A => n13948, B => 
                           n17078, ZN => n17089);
   U1206 : AOI222_X1 port map( A1 => n17079, A2 => n14457, B1 => n17087, B2 => 
                           n14420, C1 => n17089, C2 => n14331, ZN => n17093);
   U1207 : OAI22_X1 port map( A1 => n14389, A2 => n17093, B1 => n17092, B2 => 
                           n18182, ZN => n17082);
   U1208 : OAI22_X1 port map( A1 => n14134, A2 => n17091, B1 => n14332, B2 => 
                           n17080, ZN => n17081);
   U1209 : AOI211_X1 port map( C1 => n18176, C2 => n17096, A => n17082, B => 
                           n17081, ZN => n17099);
   U1210 : OAI22_X1 port map( A1 => n14401, A2 => n17099, B1 => n17086, B2 => 
                           n14137, ZN => n17083);
   U1211 : AOI211_X1 port map( C1 => n17085, C2 => n18192, A => n17084, B => 
                           n17083, ZN => n17106);
   U1212 : INV_X1 port map( A => n17086, ZN => n17103);
   U1213 : OAI211_X1 port map( C1 => n14231, C2 => n13942, A => n13941, B => 
                           n13940, ZN => n17088);
   U1214 : AOI222_X1 port map( A1 => n17089, A2 => n14420, B1 => n17088, B2 => 
                           n14188, C1 => n17087, C2 => n14456, ZN => n17090);
   U1215 : OAI22_X1 port map( A1 => n14417, A2 => n17091, B1 => n14389, B2 => 
                           n17090, ZN => n17095);
   U1216 : OAI22_X1 port map( A1 => n14134, A2 => n17093, B1 => n17092, B2 => 
                           n18226, ZN => n17094);
   U1217 : AOI211_X1 port map( C1 => n14220, C2 => n17096, A => n17095, B => 
                           n17094, ZN => n17097);
   U1218 : OAI22_X1 port map( A1 => n14402, A2 => n17098, B1 => n17097, B2 => 
                           n18183, ZN => n17102);
   U1219 : OAI22_X1 port map( A1 => n14137, A2 => n17100, B1 => n14136, B2 => 
                           n17099, ZN => n17101);
   U1220 : AOI211_X1 port map( C1 => n17103, C2 => n18192, A => n17102, B => 
                           n17101, ZN => n17104);
   U1221 : OAI22_X1 port map( A1 => n17106, A2 => n18191, B1 => n17104, B2 => 
                           n18216, ZN => n17105);
   U1222 : AOI21_X1 port map( B1 => n14230, B2 => n17116, A => n17105, ZN => 
                           n17109);
   U1223 : INV_X1 port map( A => n17106, ZN => n17108);
   U1224 : INV_X1 port map( A => n17107, ZN => n17114);
   U1225 : AOI222_X1 port map( A1 => n17108, A2 => n14381, B1 => n17116, B2 => 
                           n14139, C1 => n17114, C2 => n14229, ZN => n17127);
   U1226 : OAI22_X1 port map( A1 => n14400, A2 => n17109, B1 => n17127, B2 => 
                           n18214, ZN => n17118);
   U1227 : AOI22_X1 port map( A1 => n14398, A2 => n17122, B1 => n14375, B2 => 
                           n17121, ZN => n17113);
   U1228 : AOI22_X1 port map( A1 => n13895, A2 => n17111, B1 => n14129, B2 => 
                           n17110, ZN => n17112);
   U1229 : OAI211_X1 port map( C1 => n17123, C2 => n14136, A => n17113, B => 
                           n17112, ZN => n17120);
   U1230 : AOI222_X1 port map( A1 => n17115, A2 => n14381, B1 => n17119, B2 => 
                           n14139, C1 => n17120, C2 => n14229, ZN => n17129);
   U1231 : AOI222_X1 port map( A1 => n17116, A2 => n14381, B1 => n17115, B2 => 
                           n14229, C1 => n17114, C2 => n14139, ZN => n17186);
   U1232 : OAI22_X1 port map( A1 => n17129, A2 => n14377, B1 => n17186, B2 => 
                           n14232, ZN => n17117);
   U1233 : AOI211_X1 port map( C1 => n17198, C2 => n18207, A => n17118, B => 
                           n17117, ZN => n17133);
   U1234 : INV_X1 port map( A => n17119, ZN => n17126);
   U1235 : INV_X1 port map( A => n17120, ZN => n17251);
   U1236 : INV_X1 port map( A => n17121, ZN => n17309);
   U1237 : INV_X1 port map( A => n17122, ZN => n17310);
   U1238 : OAI22_X1 port map( A1 => n17309, A2 => n18203, B1 => n17310, B2 => 
                           n14403, ZN => n17125);
   U1239 : OAI22_X1 port map( A1 => n17123, A2 => n14401, B1 => n17294, B2 => 
                           n14136, ZN => n17124);
   U1240 : AOI211_X1 port map( C1 => n18192, C2 => n17332, A => n17125, B => 
                           n17124, ZN => n17271);
   U1241 : OAI222_X1 port map( A1 => n17126, A2 => n14133, B1 => n17251, B2 => 
                           n14382, C1 => n14330, C2 => n17271, ZN => n17240);
   U1242 : INV_X1 port map( A => n17127, ZN => n17128);
   U1243 : AOI22_X1 port map( A1 => n14222, A2 => n17240, B1 => n18190, B2 => 
                           n17128, ZN => n17131);
   U1244 : INV_X1 port map( A => n17129, ZN => n17222);
   U1245 : AOI22_X1 port map( A1 => n14385, A2 => n17198, B1 => n14394, B2 => 
                           n17222, ZN => n17130);
   U1246 : OAI211_X1 port map( C1 => n17186, C2 => n18214, A => n17131, B => 
                           n17130, ZN => n17139);
   U1247 : NAND3_X1 port map( A1 => n14270, A2 => n14335, A3 => n17139, ZN => 
                           n17132);
   U1248 : OAI211_X1 port map( C1 => n14276, C2 => n17133, A => n14165, B => 
                           n17132, ZN => OUTALU(31));
   U1249 : AOI22_X1 port map( A1 => DATA2(30), A2 => n17493, B1 => n17713, B2 
                           => n1869, ZN => n17136);
   U1250 : INV_X1 port map( A => DATA2(30), ZN => n17771);
   U1251 : AOI22_X1 port map( A1 => DATA1(30), A2 => n17771, B1 => DATA2(30), 
                           B2 => n17702, ZN => n17618);
   U1252 : INV_X1 port map( A => n17618, ZN => n17696);
   U1253 : AOI22_X1 port map( A1 => n14011, A2 => n6095, B1 => n18171, B2 => 
                           n17696, ZN => n17135);
   U1254 : NAND3_X1 port map( A1 => DATA1(31), A2 => n1869, A3 => n17339, ZN =>
                           n17134);
   U1255 : OAI211_X1 port map( C1 => n17136, C2 => n17702, A => n17135, B => 
                           n17134, ZN => n8601);
   U1256 : NOR3_X1 port map( A1 => n17138, A2 => n18230, A3 => n17137, ZN => 
                           n12158);
   U1257 : AOI211_X1 port map( C1 => n14418, C2 => n17139, A => n13938, B => 
                           n14269, ZN => n17141);
   U1258 : OR2_X1 port map( A1 => n14338, A2 => n14424, ZN => n17140);
   U1259 : OAI211_X1 port map( C1 => n14450, C2 => n13937, A => n17141, B => 
                           n17140, ZN => OUTALU(30));
   U1260 : NAND2_X1 port map( A1 => n17339, A2 => n18194, ZN => n17709);
   U1261 : INV_X1 port map( A => n17709, ZN => n17142);
   U1262 : AOI211_X1 port map( C1 => n17144, C2 => n14461, A => n17143, B => 
                           n17142, ZN => n8600);
   U1263 : AOI211_X1 port map( C1 => n17146, C2 => n17150, A => n17145, B => 
                           n1866, ZN => n17156);
   U1264 : AOI22_X1 port map( A1 => DATA2(2), A2 => n14327, B1 => n14451, B2 =>
                           n18079, ZN => n17623);
   U1265 : INV_X1 port map( A => n17623, ZN => n17154);
   U1266 : OAI211_X1 port map( C1 => n14336, C2 => n17517, A => DATA2(2), B => 
                           n17493, ZN => n17153);
   U1267 : NOR2_X1 port map( A1 => n17147, A2 => n17336, ZN => n17149);
   U1268 : AOI211_X1 port map( C1 => n17150, C2 => n17149, A => n17335, B => 
                           n17148, ZN => n17151);
   U1269 : INV_X1 port map( A => n17151, ZN => n17152);
   U1270 : OAI211_X1 port map( C1 => n17154, C2 => n17521, A => n17153, B => 
                           n17152, ZN => n17155);
   U1271 : AOI211_X1 port map( C1 => n14170, C2 => n17538, A => n17156, B => 
                           n17155, ZN => n8599);
   U1272 : INV_X1 port map( A => n1862, ZN => n17732);
   U1273 : OAI22_X1 port map( A1 => n17732, A2 => n1896, B1 => n17731, B2 => 
                           n17728, ZN => n12189);
   U1274 : OAI22_X1 port map( A1 => n14227, A2 => n17158, B1 => n14232, B2 => 
                           n17157, ZN => n17172);
   U1275 : AOI22_X1 port map( A1 => n13893, A2 => n17739, B1 => n14356, B2 => 
                           n17738, ZN => n17164);
   U1276 : INV_X1 port map( A => n17159, ZN => n17161);
   U1277 : OAI22_X1 port map( A1 => n14231, A2 => n13934, B1 => n14391, B2 => 
                           n14405, ZN => n17160);
   U1278 : AOI211_X1 port map( C1 => n14364, C2 => n14406, A => n13933, B => 
                           n17160, ZN => n17740);
   U1279 : OAI222_X1 port map( A1 => n14228, A2 => n17361, B1 => n14373, B2 => 
                           n17161, C1 => n14390, C2 => n17740, ZN => n17737);
   U1280 : AOI22_X1 port map( A1 => n14220, A2 => n17162, B1 => n14130, B2 => 
                           n17737, ZN => n17163);
   U1281 : OAI211_X1 port map( C1 => n14225, C2 => n17165, A => n17164, B => 
                           n17163, ZN => n17749);
   U1282 : AOI22_X1 port map( A1 => n14129, A2 => n17749, B1 => n14387, B2 => 
                           n17736, ZN => n17168);
   U1283 : AOI22_X1 port map( A1 => n14398, A2 => n17166, B1 => n13894, B2 => 
                           n17748, ZN => n17167);
   U1284 : OAI211_X1 port map( C1 => n14458, C2 => n17169, A => n17168, B => 
                           n17167, ZN => n17754);
   U1285 : AOI222_X1 port map( A1 => n17754, A2 => n14381, B1 => n17371, B2 => 
                           n14139, C1 => n17170, C2 => n14229, ZN => n17760);
   U1286 : OAI22_X1 port map( A1 => n14400, A2 => n17760, B1 => n14397, B2 => 
                           n17373, ZN => n17171);
   U1287 : OAI21_X1 port map( B1 => n17172, B2 => n17171, A => n14386, ZN => 
                           n17173);
   U1288 : OAI211_X1 port map( C1 => n14276, C2 => n13936, A => n13935, B => 
                           n17173, ZN => OUTALU(2));
   U1289 : NOR2_X1 port map( A1 => DATA2(29), A2 => n17247, ZN => n17697);
   U1290 : NAND2_X1 port map( A1 => DATA2(29), A2 => n17247, ZN => n17698);
   U1291 : INV_X1 port map( A => n17698, ZN => n17556);
   U1292 : OR2_X1 port map( A1 => n17697, A2 => n17556, ZN => n17174);
   U1293 : AOI22_X1 port map( A1 => n17538, A2 => n14013, B1 => n18171, B2 => 
                           n17174, ZN => n8596);
   U1294 : OAI21_X1 port map( B1 => n17530, B2 => n17247, A => n17424, ZN => 
                           n17178);
   U1295 : NAND2_X1 port map( A1 => DATA1(29), A2 => n17713, ZN => n17176);
   U1296 : NAND2_X1 port map( A1 => DATA1(30), A2 => n17339, ZN => n17175);
   U1297 : OAI211_X1 port map( C1 => n17276, C2 => n17206, A => n17176, B => 
                           n17175, ZN => n17177);
   U1298 : AOI22_X1 port map( A1 => DATA2(29), A2 => n17178, B1 => n1869, B2 =>
                           n17177, ZN => n8595);
   U1299 : OAI22_X1 port map( A1 => n17182, A2 => n17181, B1 => n17180, B2 => 
                           n17179, ZN => n12213);
   U1300 : INV_X1 port map( A => n17183, ZN => n17184);
   U1301 : AOI21_X1 port map( B1 => n8847, B2 => n17185, A => n17184, ZN => 
                           n12212);
   U1302 : INV_X1 port map( A => n17186, ZN => n17187);
   U1303 : AOI22_X1 port map( A1 => n14131, A2 => n17187, B1 => n14138, B2 => 
                           n17198, ZN => n17189);
   U1304 : AOI22_X1 port map( A1 => n14394, A2 => n17240, B1 => n14385, B2 => 
                           n17222, ZN => n17188);
   U1305 : AOI21_X1 port map( B1 => n17189, B2 => n17188, A => n14276, ZN => 
                           n17190);
   U1306 : AOI211_X1 port map( C1 => n13930, C2 => n14167, A => n14164, B => 
                           n17190, ZN => n17191);
   U1307 : NAND3_X1 port map( A1 => n13932, A2 => n13931, A3 => n17191, ZN => 
                           OUTALU(29));
   U1308 : INV_X1 port map( A => DATA2(28), ZN => n17773);
   U1309 : NOR3_X1 port map( A1 => n18162, A2 => n17773, A3 => n17695, ZN => 
                           n17197);
   U1310 : AOI22_X1 port map( A1 => DATA1(28), A2 => n17773, B1 => DATA2(28), 
                           B2 => n17695, ZN => n17615);
   U1311 : OAI22_X1 port map( A1 => n17206, A2 => n17192, B1 => n17702, B2 => 
                           n17276, ZN => n17193);
   U1312 : AOI211_X1 port map( C1 => n17713, C2 => DATA1(28), A => n17194, B =>
                           n17193, ZN => n17195);
   U1313 : OAI22_X1 port map( A1 => n17615, A2 => n17521, B1 => n17195, B2 => 
                           n17292, ZN => n17196);
   U1314 : AOI211_X1 port map( C1 => n17538, C2 => n14015, A => n17197, B => 
                           n17196, ZN => n12230);
   U1315 : AOI222_X1 port map( A1 => n17198, A2 => n14131, B1 => n17240, B2 => 
                           n14385, C1 => n17222, C2 => n14138, ZN => n17199);
   U1316 : OAI211_X1 port map( C1 => n14276, C2 => n17199, A => n14163, B => 
                           n13929, ZN => OUTALU(28));
   U1317 : NAND2_X1 port map( A1 => n17260, A2 => n17200, ZN => n17217);
   U1318 : INV_X1 port map( A => n17217, ZN => n17221);
   U1319 : AOI21_X1 port map( B1 => n17518, B2 => DATA2(27), A => n17517, ZN =>
                           n17210);
   U1320 : NOR2_X1 port map( A1 => DATA2(27), A2 => n17209, ZN => n17691);
   U1321 : INV_X1 port map( A => n17691, ZN => n17201);
   U1322 : NAND2_X1 port map( A1 => DATA2(27), A2 => n17209, ZN => n17692);
   U1323 : NAND2_X1 port map( A1 => n17201, A2 => n17692, ZN => n17552);
   U1324 : AOI22_X1 port map( A1 => n17538, A2 => n14017, B1 => n18171, B2 => 
                           n17552, ZN => n17208);
   U1325 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(30), A => n17203, B =>
                           n17202, ZN => n17205);
   U1326 : OAI211_X1 port map( C1 => n17264, C2 => n17206, A => n17205, B => 
                           n17204, ZN => n17224);
   U1327 : NAND3_X1 port map( A1 => n17352, A2 => n1869, A3 => n17224, ZN => 
                           n17207);
   U1328 : OAI211_X1 port map( C1 => n17210, C2 => n17209, A => n17208, B => 
                           n17207, ZN => n17219);
   U1329 : AND2_X1 port map( A1 => n17258, A2 => n17211, ZN => n17212);
   U1330 : OAI21_X1 port map( B1 => n17214, B2 => n17213, A => n17212, ZN => 
                           n17215);
   U1331 : OAI21_X1 port map( B1 => n17217, B2 => n17216, A => n17215, ZN => 
                           n17218);
   U1332 : AOI211_X1 port map( C1 => n17221, C2 => n17220, A => n17219, B => 
                           n17218, ZN => n12246);
   U1333 : AOI22_X1 port map( A1 => n14138, A2 => n17240, B1 => n14131, B2 => 
                           n17222, ZN => n17223);
   U1334 : OAI21_X1 port map( B1 => n14276, B2 => n17223, A => n13928, ZN => 
                           OUTALU(27));
   U1335 : INV_X1 port map( A => n17224, ZN => n17250);
   U1336 : OAI211_X1 port map( C1 => n17264, C2 => n17702, A => n17226, B => 
                           n17225, ZN => n17227);
   U1337 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(29), A => n17228, B =>
                           n17227, ZN => n17267);
   U1338 : OAI22_X1 port map( A1 => n17250, A2 => n17349, B1 => n17267, B2 => 
                           n17318, ZN => n17229);
   U1339 : NAND2_X1 port map( A1 => n1869, A2 => n17229, ZN => n12255);
   U1340 : INV_X1 port map( A => DATA2(26), ZN => n17775);
   U1341 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2(26), B1 => n17775, 
                           B2 => n17689, ZN => n17684);
   U1342 : NOR3_X1 port map( A1 => n18162, A2 => n17775, A3 => n17689, ZN => 
                           n17239);
   U1343 : NAND2_X1 port map( A1 => n14019, A2 => n17538, ZN => n17237);
   U1344 : OAI211_X1 port map( C1 => n17234, C2 => n17231, A => n17258, B => 
                           n17230, ZN => n17236);
   U1345 : OAI211_X1 port map( C1 => n17234, C2 => n17233, A => n17260, B => 
                           n17232, ZN => n17235);
   U1346 : NAND3_X1 port map( A1 => n17237, A2 => n17236, A3 => n17235, ZN => 
                           n17238);
   U1347 : AOI211_X1 port map( C1 => n18171, C2 => n17684, A => n17239, B => 
                           n17238, ZN => n12254);
   U1348 : NAND3_X1 port map( A1 => n14418, A2 => n14131, A3 => n17240, ZN => 
                           n17241);
   U1349 : NAND3_X1 port map( A1 => n14268, A2 => n13927, A3 => n17241, ZN => 
                           OUTALU(26));
   U1350 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n17493, 
                           ZN => n8838);
   U1351 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n17257);
   U1352 : INV_X1 port map( A => n17257, ZN => n17244);
   U1353 : OAI211_X1 port map( C1 => n17244, C2 => n17243, A => n17258, B => 
                           n17242, ZN => n8946);
   U1354 : OAI211_X1 port map( C1 => n17264, C2 => n17247, A => n17246, B => 
                           n17245, ZN => n17248);
   U1355 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(28), A => n17249, B =>
                           n17248, ZN => n17280);
   U1356 : OAI222_X1 port map( A1 => n17318, A2 => n17280, B1 => n17718, B2 => 
                           n17267, C1 => n17315, C2 => n17250, ZN => n17319);
   U1357 : NAND3_X1 port map( A1 => n1869, A2 => n18159, A3 => n17319, ZN => 
                           n12263);
   U1358 : OAI22_X1 port map( A1 => n17251, A2 => n14133, B1 => n17271, B2 => 
                           n14382, ZN => n17252);
   U1359 : INV_X1 port map( A => n17252, ZN => n17255);
   U1360 : NAND2_X1 port map( A1 => n14162, A2 => n14267, ZN => n17253);
   U1361 : NOR3_X1 port map( A1 => n13926, A2 => n14413, A3 => n17253, ZN => 
                           n17254);
   U1362 : OAI211_X1 port map( C1 => n17255, C2 => n18212, A => n14161, B => 
                           n17254, ZN => OUTALU(25));
   U1363 : NAND3_X1 port map( A1 => n17258, A2 => n17257, A3 => n17256, ZN => 
                           n8837);
   U1364 : NAND2_X1 port map( A1 => n17260, A2 => n17259, ZN => n8945);
   U1365 : AOI22_X1 port map( A1 => DATA2(24), A2 => n17518, B1 => 
                           DATA2_I_24_port, B2 => n17260, ZN => n17261);
   U1366 : AOI21_X1 port map( B1 => n17261, B2 => n17424, A => n17683, ZN => 
                           n17270);
   U1367 : INV_X1 port map( A => DATA2(24), ZN => n17777);
   U1368 : AOI22_X1 port map( A1 => DATA1(24), A2 => n17777, B1 => DATA2(24), 
                           B2 => n17683, ZN => n17610);
   U1369 : OAI211_X1 port map( C1 => n17264, C2 => n17695, A => n17263, B => 
                           n17262, ZN => n17265);
   U1370 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(27), A => n17266, B =>
                           n17265, ZN => n17302);
   U1371 : OAI222_X1 port map( A1 => n17318, A2 => n17302, B1 => n17718, B2 => 
                           n17280, C1 => n17315, C2 => n17267, ZN => n18124);
   U1372 : AOI22_X1 port map( A1 => n18118, A2 => n17319, B1 => n18159, B2 => 
                           n18124, ZN => n17268);
   U1373 : OAI22_X1 port map( A1 => n17610, A2 => n17521, B1 => n17268, B2 => 
                           n17292, ZN => n17269);
   U1374 : AOI211_X1 port map( C1 => n14026, C2 => n17538, A => n17270, B => 
                           n17269, ZN => n12273);
   U1375 : OR3_X1 port map( A1 => n14133, A2 => n17271, A3 => n14276, ZN => 
                           n17272);
   U1376 : NAND4_X1 port map( A1 => n13925, A2 => n14160, A3 => n14266, A4 => 
                           n17272, ZN => OUTALU(24));
   U1377 : AOI21_X1 port map( B1 => DATA2(23), B2 => n17518, A => n17517, ZN =>
                           n8834);
   U1378 : NAND2_X1 port map( A1 => n17538, A2 => n14029, ZN => n8944);
   U1379 : OAI211_X1 port map( C1 => n17276, C2 => n17275, A => n17274, B => 
                           n17273, ZN => n17277);
   U1380 : AOI211_X1 port map( C1 => n17279, C2 => DATA1(26), A => n17278, B =>
                           n17277, ZN => n17314);
   U1381 : OAI222_X1 port map( A1 => n17318, A2 => n17314, B1 => n17718, B2 => 
                           n17302, C1 => n17315, C2 => n17280, ZN => n18129);
   U1382 : AOI222_X1 port map( A1 => n18129, A2 => n18159, B1 => n18124, B2 => 
                           n18118, C1 => n17319, C2 => n18116, ZN => n17293);
   U1383 : NOR2_X1 port map( A1 => DATA2(23), A2 => n1882, ZN => n17679);
   U1384 : INV_X1 port map( A => n17679, ZN => n17281);
   U1385 : NAND2_X1 port map( A1 => DATA2(23), A2 => n1882, ZN => n17680);
   U1386 : NAND2_X1 port map( A1 => n17281, A2 => n17680, ZN => n17551);
   U1387 : NOR2_X1 port map( A1 => n17288, A2 => n17300, ZN => n17282);
   U1388 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, B1 => 
                           n1809, B2 => n18174, ZN => n17284);
   U1389 : OAI22_X1 port map( A1 => n17286, A2 => n17413, B1 => n17284, B2 => 
                           n17409, ZN => n17298);
   U1390 : AOI22_X1 port map( A1 => n18171, A2 => n17551, B1 => n17282, B2 => 
                           n17298, ZN => n17291);
   U1391 : INV_X1 port map( A => n17283, ZN => n17289);
   U1392 : INV_X1 port map( A => n17409, ZN => n18175);
   U1393 : AND2_X1 port map( A1 => n18175, A2 => n17284, ZN => n17285);
   U1394 : AOI211_X1 port map( C1 => n17286, C2 => n18173, A => n17285, B => 
                           n17300, ZN => n17299);
   U1395 : OAI21_X1 port map( B1 => n17289, B2 => n17299, A => n17288, ZN => 
                           n17287);
   U1396 : OAI211_X1 port map( C1 => n17289, C2 => n17288, A => n17769, B => 
                           n17287, ZN => n17290);
   U1397 : OAI211_X1 port map( C1 => n17293, C2 => n17292, A => n17291, B => 
                           n17290, ZN => n12292);
   U1398 : OAI22_X1 port map( A1 => n14401, A2 => n17294, B1 => n17310, B2 => 
                           n14136, ZN => n17296);
   U1399 : INV_X1 port map( A => n17332, ZN => n17308);
   U1400 : OAI22_X1 port map( A1 => n14137, A2 => n17308, B1 => n17309, B2 => 
                           n14403, ZN => n17295);
   U1401 : AOI221_X1 port map( B1 => n17296, B2 => n14418, C1 => n17295, C2 => 
                           n14418, A => n14264, ZN => n17297);
   U1402 : OAI211_X1 port map( C1 => n14159, C2 => n14439, A => n14265, B => 
                           n17297, ZN => OUTALU(23));
   U1403 : AOI22_X1 port map( A1 => DATA1(22), A2 => DATA2(22), B1 => n17779, 
                           B2 => n17675, ZN => n17608);
   U1404 : AOI22_X1 port map( A1 => n14032, A2 => n17538, B1 => n18171, B2 => 
                           n17608, ZN => n8588);
   U1405 : INV_X1 port map( A => n17298, ZN => n17301);
   U1406 : AOI21_X1 port map( B1 => n17301, B2 => n17300, A => n17299, ZN => 
                           n8587);
   U1407 : INV_X1 port map( A => n17316, ZN => n17304);
   U1408 : OAI22_X1 port map( A1 => n17302, A2 => n17716, B1 => n17314, B2 => 
                           n17349, ZN => n17303);
   U1409 : AOI21_X1 port map( B1 => n17305, B2 => n17304, A => n17303, ZN => 
                           n18122);
   U1410 : AOI22_X1 port map( A1 => n18144, A2 => n17319, B1 => n18116, B2 => 
                           n18124, ZN => n17306);
   U1411 : OAI21_X1 port map( B1 => n18137, B2 => n18122, A => n17306, ZN => 
                           n17307);
   U1412 : AOI21_X1 port map( B1 => n18118, B2 => n18129, A => n17307, ZN => 
                           n12306);
   U1413 : OAI222_X1 port map( A1 => n14401, A2 => n17310, B1 => n14136, B2 => 
                           n17309, C1 => n14403, C2 => n17308, ZN => n17311);
   U1414 : AOI211_X1 port map( C1 => n14418, C2 => n17311, A => n14158, B => 
                           n14184, ZN => n17312);
   U1415 : OAI211_X1 port map( C1 => n14275, C2 => n14157, A => n13924, B => 
                           n17312, ZN => OUTALU(22));
   U1416 : INV_X1 port map( A => n17313, ZN => n17317);
   U1417 : OAI222_X1 port map( A1 => n17318, A2 => n17317, B1 => n17718, B2 => 
                           n17316, C1 => n17315, C2 => n17314, ZN => n18115);
   U1418 : AOI22_X1 port map( A1 => n18116, A2 => n18129, B1 => n18159, B2 => 
                           n18115, ZN => n17321);
   U1419 : AOI22_X1 port map( A1 => n18144, A2 => n18124, B1 => n17319, B2 => 
                           n18123, ZN => n17320);
   U1420 : OAI211_X1 port map( C1 => n18122, C2 => n18148, A => n17321, B => 
                           n17320, ZN => n12392);
   U1421 : NAND3_X1 port map( A1 => n1897, A2 => n1869, A3 => n12392, ZN => 
                           n12313);
   U1422 : OAI211_X1 port map( C1 => n17326, C2 => n17323, A => n18173, B => 
                           n17322, ZN => n17330);
   U1423 : OAI211_X1 port map( C1 => n17326, C2 => n17325, A => n18175, B => 
                           n17324, ZN => n17329);
   U1424 : NAND3_X1 port map( A1 => DATA2(20), A2 => DATA1(20), A3 => n17493, 
                           ZN => n17328);
   U1425 : INV_X1 port map( A => DATA2(20), ZN => n17781);
   U1426 : NAND2_X1 port map( A1 => DATA1(20), A2 => n17781, ZN => n17604);
   U1427 : INV_X1 port map( A => n17604, ZN => n17548);
   U1428 : NOR2_X1 port map( A1 => n17781, A2 => DATA1(20), ZN => n17669);
   U1429 : OAI21_X1 port map( B1 => n17548, B2 => n17669, A => n18171, ZN => 
                           n17327);
   U1430 : NAND4_X1 port map( A1 => n17330, A2 => n17329, A3 => n17328, A4 => 
                           n17327, ZN => n17331);
   U1431 : AOI21_X1 port map( B1 => n17538, B2 => n14038, A => n17331, ZN => 
                           n12325);
   U1432 : AOI22_X1 port map( A1 => n14341, A2 => n13985, B1 => n13986, B2 => 
                           n14362, ZN => n17334);
   U1433 : NAND3_X1 port map( A1 => n18189, A2 => n17332, A3 => n18210, ZN => 
                           n17333);
   U1434 : OAI211_X1 port map( C1 => n14275, C2 => n17334, A => n14263, B => 
                           n17333, ZN => OUTALU(20));
   U1435 : AOI211_X1 port map( C1 => n17531, C2 => n17340, A => n17336, B => 
                           n17335, ZN => n17338);
   U1436 : NOR2_X1 port map( A1 => n14463, A2 => n18059, ZN => n17574);
   U1437 : INV_X1 port map( A => n17574, ZN => n17626);
   U1438 : NAND2_X1 port map( A1 => n18059, A2 => n18194, ZN => n17622);
   U1439 : AOI21_X1 port map( B1 => n17626, B2 => n17622, A => n17521, ZN => 
                           n17337);
   U1440 : AOI211_X1 port map( C1 => n13848, C2 => n17538, A => n17338, B => 
                           n17337, ZN => n8581);
   U1441 : AOI21_X1 port map( B1 => n17713, B2 => n1868, A => n17517, ZN => 
                           n17529);
   U1442 : OAI21_X1 port map( B1 => n18059, B2 => n17530, A => n17529, ZN => 
                           n8832);
   U1443 : NAND3_X1 port map( A1 => n14461, A2 => n17339, A3 => n1868, ZN => 
                           n8831);
   U1444 : OAI221_X1 port map( B1 => n17532, B2 => n17342, C1 => n17341, C2 => 
                           n17340, A => n17537, ZN => n8553);
   U1445 : AOI211_X1 port map( C1 => n17345, C2 => n18194, A => n17344, B => 
                           n17343, ZN => n17347);
   U1446 : OAI211_X1 port map( C1 => n14451, C2 => n17348, A => n17347, B => 
                           n17346, ZN => n17714);
   U1447 : OAI22_X1 port map( A1 => n17350, A2 => n17716, B1 => n17715, B2 => 
                           n17349, ZN => n17351);
   U1448 : AOI21_X1 port map( B1 => n17352, B2 => n17714, A => n17351, ZN => 
                           n17727);
   U1449 : INV_X1 port map( A => n17724, ZN => n17353);
   U1450 : OAI22_X1 port map( A1 => n18137, A2 => n17727, B1 => n17353, B2 => 
                           n18150, ZN => n17357);
   U1451 : OAI22_X1 port map( A1 => n18155, A2 => n17355, B1 => n17354, B2 => 
                           n18152, ZN => n17356);
   U1452 : AOI211_X1 port map( C1 => n18118, C2 => n17722, A => n17357, B => 
                           n17356, ZN => n17729);
   U1453 : OAI22_X1 port map( A1 => n17731, A2 => n1896, B1 => n17729, B2 => 
                           n17499, ZN => n17360);
   U1454 : OAI22_X1 port map( A1 => n17358, A2 => n1895, B1 => n17732, B2 => 
                           n9020, ZN => n17359);
   U1455 : AOI211_X1 port map( C1 => n1898, C2 => n1861, A => n17360, B => 
                           n17359, ZN => n12722);
   U1456 : OAI222_X1 port map( A1 => n14228, A2 => n17740, B1 => n14373, B2 => 
                           n17361, C1 => n14390, C2 => n13921, ZN => n17741);
   U1457 : INV_X1 port map( A => n17741, ZN => n17365);
   U1458 : AOI22_X1 port map( A1 => n18176, A2 => n17739, B1 => n17738, B2 => 
                           n13893, ZN => n17364);
   U1459 : AOI22_X1 port map( A1 => n17362, A2 => n14221, B1 => n17737, B2 => 
                           n14384, ZN => n17363);
   U1460 : OAI211_X1 port map( C1 => n18196, C2 => n17365, A => n17364, B => 
                           n17363, ZN => n17746);
   U1461 : AOI22_X1 port map( A1 => n17736, A2 => n13894, B1 => n17746, B2 => 
                           n14129, ZN => n17366);
   U1462 : INV_X1 port map( A => n17366, ZN => n17370);
   U1463 : OAI22_X1 port map( A1 => n14458, A2 => n17368, B1 => n17367, B2 => 
                           n18215, ZN => n17369);
   U1464 : AOI211_X1 port map( C1 => n14343, C2 => n17749, A => n17370, B => 
                           n17369, ZN => n17756);
   U1465 : AOI22_X1 port map( A1 => n14139, A2 => n17754, B1 => n14230, B2 => 
                           n17371, ZN => n17372);
   U1466 : OAI21_X1 port map( B1 => n17756, B2 => n18216, A => n17372, ZN => 
                           n17763);
   U1467 : INV_X1 port map( A => n17373, ZN => n17757);
   U1468 : AOI22_X1 port map( A1 => n18190, A2 => n17763, B1 => n18220, B2 => 
                           n17757, ZN => n17376);
   U1469 : AOI22_X1 port map( A1 => n14222, A2 => n17374, B1 => n18207, B2 => 
                           n17758, ZN => n17375);
   U1470 : OAI211_X1 port map( C1 => n17760, C2 => n14397, A => n17376, B => 
                           n17375, ZN => n17764);
   U1471 : AOI22_X1 port map( A1 => n14462, A2 => n14155, B1 => n14386, B2 => 
                           n17764, ZN => n17377);
   U1472 : NAND4_X1 port map( A1 => n13922, A2 => n14154, A3 => n13867, A4 => 
                           n17377, ZN => OUTALU(1));
   U1473 : INV_X1 port map( A => DATA2(19), ZN => n17782);
   U1474 : OAI21_X1 port map( B1 => n17530, B2 => n17782, A => n17424, ZN => 
                           n17378);
   U1475 : AOI22_X1 port map( A1 => DATA1(19), A2 => n17378, B1 => n17538, B2 
                           => n14041, ZN => n8579);
   U1476 : NOR2_X1 port map( A1 => DATA2(19), A2 => n17379, ZN => n17601);
   U1477 : NAND2_X1 port map( A1 => DATA2(19), A2 => n17379, ZN => n17667);
   U1478 : INV_X1 port map( A => n17667, ZN => n17546);
   U1479 : OAI21_X1 port map( B1 => n17601, B2 => n17546, A => n18171, ZN => 
                           n8830);
   U1480 : XNOR2_X1 port map( A => n17380, B => n17381, ZN => n17384);
   U1481 : XNOR2_X1 port map( A => n17382, B => n17381, ZN => n17383);
   U1482 : OAI22_X1 port map( A1 => n17413, A2 => n17384, B1 => n17409, B2 => 
                           n17383, ZN => n8578);
   U1483 : AOI222_X1 port map( A1 => n14341, A2 => n13986, B1 => n14363, B2 => 
                           n13985, C1 => n14440, C2 => n14362, ZN => n17391);
   U1484 : AOI22_X1 port map( A1 => n14384, A2 => n17403, B1 => n14130, B2 => 
                           n17385, ZN => n17387);
   U1485 : AOI22_X1 port map( A1 => n13893, A2 => n17417, B1 => n18176, B2 => 
                           n17429, ZN => n17386);
   U1486 : AOI21_X1 port map( B1 => n17387, B2 => n17386, A => n14276, ZN => 
                           n17389);
   U1487 : NAND2_X1 port map( A1 => n14153, A2 => n13920, ZN => n17388);
   U1488 : NOR3_X1 port map( A1 => n13919, A2 => n17389, A3 => n17388, ZN => 
                           n17390);
   U1489 : OAI21_X1 port map( B1 => n14275, B2 => n17391, A => n17390, ZN => 
                           OUTALU(19));
   U1490 : NAND2_X1 port map( A1 => n17393, A2 => n17392, ZN => n17398);
   U1491 : INV_X1 port map( A => n17398, ZN => n17395);
   U1492 : AOI211_X1 port map( C1 => n17395, C2 => n17412, A => n17394, B => 
                           n17413, ZN => n17402);
   U1493 : INV_X1 port map( A => DATA2(18), ZN => n17783);
   U1494 : AOI22_X1 port map( A1 => DATA1(18), A2 => n17783, B1 => DATA2(18), 
                           B2 => n17600, ZN => n17664);
   U1495 : OAI211_X1 port map( C1 => n17517, C2 => n17518, A => DATA2(18), B =>
                           DATA1(18), ZN => n17400);
   U1496 : INV_X1 port map( A => n17396, ZN => n17410);
   U1497 : OAI211_X1 port map( C1 => n17410, C2 => n17398, A => n18175, B => 
                           n17397, ZN => n17399);
   U1498 : OAI211_X1 port map( C1 => n17664, C2 => n17521, A => n17400, B => 
                           n17399, ZN => n17401);
   U1499 : AOI211_X1 port map( C1 => n17538, C2 => n14044, A => n17402, B => 
                           n17401, ZN => n12400);
   U1500 : AOI222_X1 port map( A1 => n17429, A2 => n13893, B1 => n17403, B2 => 
                           n14130, C1 => n17417, C2 => n14384, ZN => n17407);
   U1501 : AOI22_X1 port map( A1 => n14435, A2 => n13985, B1 => n13986, B2 => 
                           n14396, ZN => n17404);
   U1502 : OAI21_X1 port map( B1 => n14231, B2 => n14444, A => n17404, ZN => 
                           n17405);
   U1503 : OAI221_X1 port map( B1 => n17405, B2 => n18185, C1 => n17405, C2 => 
                           n18223, A => n14351, ZN => n17406);
   U1504 : OAI211_X1 port map( C1 => n14276, C2 => n17407, A => n14262, B => 
                           n17406, ZN => OUTALU(18));
   U1505 : INV_X1 port map( A => DATA2(17), ZN => n17784);
   U1506 : NAND2_X1 port map( A1 => DATA1(17), A2 => n17784, ZN => n17663);
   U1507 : NOR2_X1 port map( A1 => DATA1(17), A2 => n17784, ZN => n17599);
   U1508 : INV_X1 port map( A => n17599, ZN => n17662);
   U1509 : NAND2_X1 port map( A1 => n17663, A2 => n17662, ZN => n17558);
   U1510 : AOI22_X1 port map( A1 => n17538, A2 => n14047, B1 => n18171, B2 => 
                           n17558, ZN => n8574);
   U1511 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n17411);
   U1512 : INV_X1 port map( A => n17408, ZN => n17416);
   U1513 : AOI211_X1 port map( C1 => n17411, C2 => n17416, A => n17410, B => 
                           n17409, ZN => n8573);
   U1514 : INV_X1 port map( A => n17412, ZN => n17414);
   U1515 : AOI211_X1 port map( C1 => n17416, C2 => n17415, A => n17414, B => 
                           n17413, ZN => n8572);
   U1516 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n17493, 
                           ZN => n8828);
   U1517 : AOI22_X1 port map( A1 => n17417, A2 => n14130, B1 => n17429, B2 => 
                           n14384, ZN => n17418);
   U1518 : INV_X1 port map( A => n17418, ZN => n17419);
   U1519 : AOI211_X1 port map( C1 => n14418, C2 => n17419, A => n13917, B => 
                           n13916, ZN => n17422);
   U1520 : NAND3_X1 port map( A1 => n14331, A2 => n14386, A3 => n17420, ZN => 
                           n17421);
   U1521 : NAND4_X1 port map( A1 => n13918, A2 => n14152, A3 => n17422, A4 => 
                           n17421, ZN => OUTALU(17));
   U1522 : INV_X1 port map( A => DATA2(16), ZN => n17785);
   U1523 : NAND2_X1 port map( A1 => DATA1(16), A2 => n17785, ZN => n17656);
   U1524 : NAND2_X1 port map( A1 => DATA2(16), A2 => n17423, ZN => n17661);
   U1525 : NAND2_X1 port map( A1 => n17656, A2 => n17661, ZN => n17559);
   U1526 : AOI22_X1 port map( A1 => n17538, A2 => n14050, B1 => n18171, B2 => 
                           n17559, ZN => n8571);
   U1527 : OAI21_X1 port map( B1 => n17530, B2 => n17785, A => n17424, ZN => 
                           n17426);
   U1528 : AOI22_X1 port map( A1 => DATA1(16), A2 => n17426, B1 => n17425, B2 
                           => n18173, ZN => n12423);
   U1529 : OAI22_X1 port map( A1 => n17428, A2 => n18198, B1 => n17427, B2 => 
                           n18177, ZN => n17431);
   U1530 : AND3_X1 port map( A1 => n17429, A2 => n14130, A3 => n14418, ZN => 
                           n17430);
   U1531 : AOI211_X1 port map( C1 => n18179, C2 => n17431, A => n14278, B => 
                           n17430, ZN => n17432);
   U1532 : NAND3_X1 port map( A1 => n14151, A2 => n13915, A3 => n17432, ZN => 
                           OUTALU(16));
   U1533 : INV_X1 port map( A => n17501, ZN => n17498);
   U1534 : INV_X1 port map( A => n17512, ZN => n17434);
   U1535 : INV_X1 port map( A => n17513, ZN => n17433);
   U1536 : OAI21_X1 port map( B1 => n17434, B2 => n17514, A => n17433, ZN => 
                           n17510);
   U1537 : NAND2_X1 port map( A1 => n17435, A2 => n17510, ZN => n17500);
   U1538 : NAND2_X1 port map( A1 => n17498, A2 => n17500, ZN => n17503);
   U1539 : NAND2_X1 port map( A1 => n17436, A2 => n17503, ZN => n18166);
   U1540 : AOI21_X1 port map( B1 => n17438, B2 => n18166, A => n17437, ZN => 
                           n17457);
   U1541 : NAND2_X1 port map( A1 => n17457, A2 => n17456, ZN => n17463);
   U1542 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n17467, B2 => n17463, ZN => n17440);
   U1543 : INV_X1 port map( A => n18163, ZN => n17515);
   U1544 : OAI21_X1 port map( B1 => n17440, B2 => n17444, A => n17515, ZN => 
                           n17439);
   U1545 : AOI21_X1 port map( B1 => n17440, B2 => n17444, A => n17439, ZN => 
                           n17449);
   U1546 : NOR2_X1 port map( A1 => n17441, A2 => DATA2(15), ZN => n17657);
   U1547 : INV_X1 port map( A => n17657, ZN => n17595);
   U1548 : NAND2_X1 port map( A1 => DATA2(15), A2 => n17441, ZN => n17659);
   U1549 : AND2_X1 port map( A1 => n17595, A2 => n17659, ZN => n17563);
   U1550 : NAND3_X1 port map( A1 => DATA2(15), A2 => DATA1(15), A3 => n17493, 
                           ZN => n17447);
   U1551 : INV_X1 port map( A => n17445, ZN => n17443);
   U1552 : INV_X1 port map( A => n17444, ZN => n17442);
   U1553 : OAI221_X1 port map( B1 => n17445, B2 => n17444, C1 => n17443, C2 => 
                           n17442, A => n17481, ZN => n17446);
   U1554 : OAI211_X1 port map( C1 => n17563, C2 => n17521, A => n17447, B => 
                           n17446, ZN => n17448);
   U1555 : AOI211_X1 port map( C1 => n14053, C2 => n17538, A => n17449, B => 
                           n17448, ZN => n12446);
   U1556 : INV_X1 port map( A => n17450, ZN => n17451);
   U1557 : AOI22_X1 port map( A1 => n14358, A2 => n17452, B1 => n14357, B2 => 
                           n17451, ZN => n17455);
   U1558 : NAND3_X1 port map( A1 => n18211, A2 => n17453, A3 => n18179, ZN => 
                           n17454);
   U1559 : OAI211_X1 port map( C1 => n14276, C2 => n17455, A => n13914, B => 
                           n17454, ZN => OUTALU(15));
   U1560 : INV_X1 port map( A => n17456, ZN => n17460);
   U1561 : AOI22_X1 port map( A1 => n17458, A2 => n17481, B1 => n17515, B2 => 
                           n17457, ZN => n17474);
   U1562 : NOR3_X1 port map( A1 => n17460, A2 => n17474, A3 => n17459, ZN => 
                           n8826);
   U1563 : NAND2_X1 port map( A1 => n14292, A2 => n16394, ZN => n17461);
   U1564 : OAI21_X1 port map( B1 => n14292, B2 => n16394, A => n17461, ZN => 
                           n18008);
   U1565 : NOR3_X1 port map( A1 => n14352, A2 => n16397, A3 => n18008, ZN => 
                           n3020);
   U1566 : AOI221_X1 port map( B1 => n14352, B2 => n16397, C1 => n18008, C2 => 
                           n16397, A => n3020, ZN => n8824);
   U1567 : AOI22_X1 port map( A1 => n17515, A2 => n17463, B1 => n17481, B2 => 
                           n17462, ZN => n17466);
   U1568 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2(14), B1 => n17787, 
                           B2 => n17655, ZN => n17650);
   U1569 : AOI22_X1 port map( A1 => n13864, A2 => n6095, B1 => n18171, B2 => 
                           n17650, ZN => n17465);
   U1570 : NAND3_X1 port map( A1 => DATA2(14), A2 => DATA1(14), A3 => n17493, 
                           ZN => n17464);
   U1571 : OAI211_X1 port map( C1 => n17467, C2 => n17466, A => n17465, B => 
                           n17464, ZN => n8942);
   U1572 : NAND2_X1 port map( A1 => n14357, A2 => n18210, ZN => n17471);
   U1573 : OAI22_X1 port map( A1 => n14134, A2 => n17488, B1 => n14339, B2 => 
                           n17487, ZN => n17468);
   U1574 : AOI211_X1 port map( C1 => n14351, C2 => n17468, A => n14150, B => 
                           n13913, ZN => n17469);
   U1575 : OAI21_X1 port map( B1 => n17471, B2 => n17470, A => n17469, ZN => 
                           OUTALU(14));
   U1576 : INV_X1 port map( A => n18166, ZN => n18164);
   U1577 : NOR3_X1 port map( A1 => n18164, A2 => n18165, A3 => n18230, ZN => 
                           n17472);
   U1578 : OAI211_X1 port map( C1 => n17473, C2 => n17483, A => n17472, B => 
                           n17476, ZN => n8823);
   U1579 : AOI21_X1 port map( B1 => n17476, B2 => n17475, A => n17474, ZN => 
                           n8821);
   U1580 : OAI22_X1 port map( A1 => n12526, A2 => n9020, B1 => n17484, B2 => 
                           n17728, ZN => n12473);
   U1581 : OAI211_X1 port map( C1 => DATA2(13), C2 => n17517, A => DATA1(13), B
                           => n17493, ZN => n12474);
   U1582 : OAI222_X1 port map( A1 => n14134, A2 => n17487, B1 => n14339, B2 => 
                           n17486, C1 => n14345, C2 => n17488, ZN => n17477);
   U1583 : AOI211_X1 port map( C1 => n14351, C2 => n17477, A => n14149, B => 
                           n14415, ZN => n17480);
   U1584 : OAI22_X1 port map( A1 => n14454, A2 => n13960, B1 => n14231, B2 => 
                           n14412, ZN => n17478);
   U1585 : OAI21_X1 port map( B1 => n13911, B2 => n17478, A => n14346, ZN => 
                           n17479);
   U1586 : NAND4_X1 port map( A1 => n13912, A2 => n14261, A3 => n17480, A4 => 
                           n17479, ZN => OUTALU(13));
   U1587 : INV_X1 port map( A => n18165, ZN => n18167);
   U1588 : INV_X1 port map( A => n17483, ZN => n17482);
   U1589 : OAI221_X1 port map( B1 => n18167, B2 => n17483, C1 => n18165, C2 => 
                           n17482, A => n17481, ZN => n8551);
   U1590 : OAI222_X1 port map( A1 => n17499, A2 => n17484, B1 => n1896, B2 => 
                           n12526, C1 => n17728, C2 => n8604, ZN => n12487);
   U1591 : AOI22_X1 port map( A1 => n14418, A2 => n13858, B1 => n14008, B2 => 
                           n13868, ZN => n17492);
   U1592 : OAI22_X1 port map( A1 => n14134, A2 => n17486, B1 => n14339, B2 => 
                           n17485, ZN => n17490);
   U1593 : OAI22_X1 port map( A1 => n14225, A2 => n17488, B1 => n14345, B2 => 
                           n17487, ZN => n17489);
   U1594 : OAI21_X1 port map( B1 => n17490, B2 => n17489, A => n14351, ZN => 
                           n17491);
   U1595 : NAND4_X1 port map( A1 => n13863, A2 => n14416, A3 => n17492, A4 => 
                           n17491, ZN => OUTALU(12));
   U1596 : AND3_X1 port map( A1 => n17493, A2 => DATA2(11), A3 => DATA1(11), ZN
                           => n17495);
   U1597 : INV_X1 port map( A => DATA2(11), ZN => n17789);
   U1598 : NOR2_X1 port map( A1 => DATA1(11), A2 => n17789, ZN => n17589);
   U1599 : INV_X1 port map( A => n17589, ZN => n17646);
   U1600 : NAND2_X1 port map( A1 => DATA1(11), A2 => n17789, ZN => n17590);
   U1601 : AOI21_X1 port map( B1 => n17646, B2 => n17590, A => n17521, ZN => 
                           n17494);
   U1602 : AOI211_X1 port map( C1 => n14080, C2 => n17538, A => n17495, B => 
                           n17494, ZN => n8567);
   U1603 : INV_X1 port map( A => n17496, ZN => n17497);
   U1604 : AOI221_X1 port map( B1 => n17498, B2 => n17497, C1 => n17501, C2 => 
                           n17496, A => n17508, ZN => n8550);
   U1605 : OAI22_X1 port map( A1 => n12526, A2 => n17728, B1 => n8604, B2 => 
                           n17499, ZN => n17505);
   U1606 : INV_X1 port map( A => n17500, ZN => n17502);
   U1607 : AOI21_X1 port map( B1 => n17502, B2 => n17501, A => n18163, ZN => 
                           n17504);
   U1608 : AOI22_X1 port map( A1 => n1868, A2 => n17505, B1 => n17504, B2 => 
                           n17503, ZN => n12509);
   U1609 : NOR2_X1 port map( A1 => n14401, A2 => n14275, ZN => n17506);
   U1610 : AOI21_X1 port map( B1 => n17506, B2 => n17524, A => n13862, ZN => 
                           n17507);
   U1611 : NAND3_X1 port map( A1 => n13910, A2 => n13909, A3 => n17507, ZN => 
                           OUTALU(11));
   U1612 : NOR2_X1 port map( A1 => n17509, A2 => n17508, ZN => n17516);
   U1613 : AOI21_X1 port map( B1 => n17515, B2 => n17510, A => n17516, ZN => 
                           n17511);
   U1614 : AOI21_X1 port map( B1 => n17513, B2 => n17512, A => n17511, ZN => 
                           n8566);
   U1615 : NAND3_X1 port map( A1 => n17515, A2 => n17514, A3 => n17513, ZN => 
                           n8820);
   U1616 : INV_X1 port map( A => n17516, ZN => n17522);
   U1617 : AOI22_X1 port map( A1 => DATA1(10), A2 => n17790, B1 => DATA2(10), 
                           B2 => n17520, ZN => n17642);
   U1618 : AOI21_X1 port map( B1 => n17518, B2 => DATA2(10), A => n17517, ZN =>
                           n17519);
   U1619 : OAI222_X1 port map( A1 => n17523, A2 => n17522, B1 => n17521, B2 => 
                           n17642, C1 => n17520, C2 => n17519, ZN => n8819);
   U1620 : NAND2_X1 port map( A1 => n17538, A2 => n13873, ZN => n8940);
   U1621 : AOI22_X1 port map( A1 => n18189, A2 => n17525, B1 => n18222, B2 => 
                           n17524, ZN => n17528);
   U1622 : NAND2_X1 port map( A1 => n14147, A2 => n14260, ZN => n17526);
   U1623 : NOR3_X1 port map( A1 => n14148, A2 => n13857, A3 => n17526, ZN => 
                           n17527);
   U1624 : OAI211_X1 port map( C1 => n17528, C2 => n18208, A => n14146, B => 
                           n17527, ZN => OUTALU(10));
   U1625 : OAI21_X1 port map( B1 => n18062, B2 => n17530, A => n17529, ZN => 
                           n17535);
   U1626 : NAND2_X1 port map( A1 => n14461, A2 => n18062, ZN => n17575);
   U1627 : NAND2_X1 port map( A1 => DATA2(0), A2 => n14329, ZN => n17625);
   U1628 : NAND2_X1 port map( A1 => n17575, A2 => n17625, ZN => n17550);
   U1629 : NOR2_X1 port map( A1 => n17532, A2 => n17531, ZN => n17536);
   U1630 : INV_X1 port map( A => n17536, ZN => n17534);
   U1631 : AOI222_X1 port map( A1 => n17535, A2 => n14461, B1 => n17550, B2 => 
                           n18171, C1 => n17534, C2 => n17533, ZN => n8818);
   U1632 : AOI22_X1 port map( A1 => n17538, A2 => n14253, B1 => n17537, B2 => 
                           n17536, ZN => n8565);
   U1633 : NOR2_X1 port map( A1 => n17540, A2 => n17539, ZN => n8626);
   U1634 : NAND2_X1 port map( A1 => FUNC(3), A2 => n8626, ZN => n12754);
   U1635 : INV_X1 port map( A => n17608, ZN => n17677);
   U1636 : INV_X1 port map( A => n17590, ZN => n17541);
   U1637 : INV_X1 port map( A => DATA2(12), ZN => n18160);
   U1638 : AOI22_X1 port map( A1 => DATA2(12), A2 => DATA1(12), B1 => n18161, 
                           B2 => n18160, ZN => n18170);
   U1639 : NOR2_X1 port map( A1 => n17541, A2 => n18170, ZN => n17648);
   U1640 : NOR4_X1 port map( A1 => n17684, A2 => n17544, A3 => n17543, A4 => 
                           n17542, ZN => n17545);
   U1641 : NAND4_X1 port map( A1 => n17677, A2 => n17664, A3 => n17648, A4 => 
                           n17545, ZN => n17571);
   U1642 : OR2_X1 port map( A1 => n17669, A2 => n17546, ZN => n17605);
   U1643 : INV_X1 port map( A => n17610, ZN => n17678);
   U1644 : INV_X1 port map( A => n17615, ZN => n17690);
   U1645 : NOR4_X1 port map( A1 => n17605, A2 => n17678, A3 => n17690, A4 => 
                           n17696, ZN => n17569);
   U1646 : INV_X1 port map( A => n17642, ZN => n17547);
   U1647 : INV_X1 port map( A => n17635, ZN => n17582);
   U1648 : NOR4_X1 port map( A1 => n17547, A2 => n17582, A3 => n17623, A4 => 
                           n17650, ZN => n17568);
   U1649 : NOR2_X1 port map( A1 => n17548, A2 => n17601, ZN => n17671);
   U1650 : NOR4_X1 port map( A1 => n17552, A2 => n17551, A3 => n17550, A4 => 
                           n17549, ZN => n17553);
   U1651 : NAND4_X1 port map( A1 => n17671, A2 => n17553, A3 => n17641, A4 => 
                           n17640, ZN => n17554);
   U1652 : NOR4_X1 port map( A1 => n17697, A2 => n17556, A3 => n17555, A4 => 
                           n17554, ZN => n17567);
   U1653 : AOI21_X1 port map( B1 => n16393, B2 => DATA2(7), A => n17557, ZN => 
                           n17585);
   U1654 : INV_X1 port map( A => n17585, ZN => n17565);
   U1655 : NOR4_X1 port map( A1 => n17561, A2 => n17560, A3 => n17559, A4 => 
                           n17558, ZN => n17562);
   U1656 : NAND4_X1 port map( A1 => n17563, A2 => n17562, A3 => n17626, A4 => 
                           n17622, ZN => n17564);
   U1657 : NOR4_X1 port map( A1 => n17589, A2 => n17636, A3 => n17565, A4 => 
                           n17564, ZN => n17566);
   U1658 : NAND4_X1 port map( A1 => n17569, A2 => n17568, A3 => n17567, A4 => 
                           n17566, ZN => n17570);
   U1659 : OAI21_X1 port map( B1 => n17571, B2 => n17570, A => n1870, ZN => 
                           n17573);
   U1660 : AOI211_X1 port map( C1 => FUNC(2), C2 => n17573, A => FUNC(1), B => 
                           n17572, ZN => n12751);
   U1661 : AOI211_X1 port map( C1 => n17622, C2 => n17575, A => n17574, B => 
                           n17623, ZN => n17576);
   U1662 : AOI21_X1 port map( B1 => n14336, B2 => n18079, A => n17576, ZN => 
                           n17577);
   U1663 : AOI22_X1 port map( A1 => DATA2(4), A2 => n14438, B1 => n17577, B2 =>
                           n17628, ZN => n17579);
   U1664 : INV_X1 port map( A => n17629, ZN => n17578);
   U1665 : AOI21_X1 port map( B1 => n17579, B2 => n17627, A => n17578, ZN => 
                           n17580);
   U1666 : OAI21_X1 port map( B1 => DATA2(5), B2 => n14453, A => n17580, ZN => 
                           n17581);
   U1667 : OAI21_X1 port map( B1 => n14465, B2 => n17797, A => n17581, ZN => 
                           n17583);
   U1668 : OAI22_X1 port map( A1 => DATA2(6), A2 => n14437, B1 => n17583, B2 =>
                           n17582, ZN => n17584);
   U1669 : AOI221_X1 port map( B1 => n17636, B2 => n17585, C1 => n17584, C2 => 
                           n17585, A => n17637, ZN => n17586);
   U1670 : OAI21_X1 port map( B1 => n17587, B2 => n17586, A => n17641, ZN => 
                           n17588);
   U1671 : AOI22_X1 port map( A1 => DATA1(10), A2 => n17790, B1 => n17642, B2 
                           => n17588, ZN => n17591);
   U1672 : AOI21_X1 port map( B1 => n17591, B2 => n17590, A => n17589, ZN => 
                           n17592);
   U1673 : AOI222_X1 port map( A1 => DATA1(12), A2 => n17592, B1 => DATA1(12), 
                           B2 => n18160, C1 => n17592, C2 => n18160, ZN => 
                           n17594);
   U1674 : AOI211_X1 port map( C1 => n17594, C2 => n17649, A => n17593, B => 
                           n17650, ZN => n17597);
   U1675 : OAI21_X1 port map( B1 => DATA2(14), B2 => n17655, A => n17595, ZN =>
                           n17596);
   U1676 : OAI211_X1 port map( C1 => n17597, C2 => n17596, A => n17661, B => 
                           n17659, ZN => n17598);
   U1677 : OAI221_X1 port map( B1 => n17599, B2 => n17656, C1 => n17599, C2 => 
                           n17598, A => n17663, ZN => n17603);
   U1678 : NOR2_X1 port map( A1 => DATA2(18), A2 => n17600, ZN => n17602);
   U1679 : AOI211_X1 port map( C1 => n17664, C2 => n17603, A => n17602, B => 
                           n17601, ZN => n17606);
   U1680 : OAI21_X1 port map( B1 => n17606, B2 => n17605, A => n17604, ZN => 
                           n17607);
   U1681 : AOI21_X1 port map( B1 => n17672, B2 => n17607, A => n17674, ZN => 
                           n17609);
   U1682 : OAI22_X1 port map( A1 => DATA2(22), A2 => n17675, B1 => n17609, B2 
                           => n17608, ZN => n17611);
   U1683 : OAI211_X1 port map( C1 => n17679, C2 => n17611, A => n17610, B => 
                           n17680, ZN => n17612);
   U1684 : OAI21_X1 port map( B1 => DATA2(24), B2 => n17683, A => n17612, ZN =>
                           n17613);
   U1685 : AOI21_X1 port map( B1 => n17686, B2 => n17613, A => n17685, ZN => 
                           n17614);
   U1686 : OAI22_X1 port map( A1 => DATA2(26), A2 => n17689, B1 => n17614, B2 
                           => n17684, ZN => n17616);
   U1687 : OAI211_X1 port map( C1 => n17691, C2 => n17616, A => n17615, B => 
                           n17692, ZN => n17617);
   U1688 : OAI21_X1 port map( B1 => DATA2(28), B2 => n17695, A => n17617, ZN =>
                           n17619);
   U1689 : OAI211_X1 port map( C1 => n17697, C2 => n17619, A => n17618, B => 
                           n17698, ZN => n17620);
   U1690 : OAI211_X1 port map( C1 => DATA2(30), C2 => n17702, A => n17620, B =>
                           n17621, ZN => n17706);
   U1691 : INV_X1 port map( A => n17621, ZN => n17704);
   U1692 : INV_X1 port map( A => n17707, ZN => n17701);
   U1693 : AOI22_X1 port map( A1 => DATA2(6), A2 => n14437, B1 => n16393, B2 =>
                           DATA2(7), ZN => n17639);
   U1694 : INV_X1 port map( A => n17622, ZN => n17624);
   U1695 : AOI211_X1 port map( C1 => n17626, C2 => n17625, A => n17624, B => 
                           n17623, ZN => n17631);
   U1696 : OAI21_X1 port map( B1 => n14327, B2 => n18079, A => n17627, ZN => 
                           n17630);
   U1697 : OAI211_X1 port map( C1 => n17631, C2 => n17630, A => n17629, B => 
                           n17628, ZN => n17632);
   U1698 : OAI211_X1 port map( C1 => n14465, C2 => n17797, A => n17633, B => 
                           n17632, ZN => n17634);
   U1699 : OAI211_X1 port map( C1 => DATA2(5), C2 => n14453, A => n17635, B => 
                           n17634, ZN => n17638);
   U1700 : AOI211_X1 port map( C1 => n17639, C2 => n17638, A => n17637, B => 
                           n17636, ZN => n17644);
   U1701 : OAI21_X1 port map( B1 => n14469, B2 => n17792, A => n17640, ZN => 
                           n17643);
   U1702 : OAI211_X1 port map( C1 => n17644, C2 => n17643, A => n17642, B => 
                           n17641, ZN => n17645);
   U1703 : OAI211_X1 port map( C1 => DATA1(10), C2 => n17790, A => n17646, B =>
                           n17645, ZN => n17647);
   U1704 : AOI22_X1 port map( A1 => DATA2(12), A2 => n18161, B1 => n17648, B2 
                           => n17647, ZN => n17653);
   U1705 : INV_X1 port map( A => n17649, ZN => n17651);
   U1706 : AOI211_X1 port map( C1 => n17653, C2 => n17652, A => n17651, B => 
                           n17650, ZN => n17654);
   U1707 : AOI21_X1 port map( B1 => DATA2(14), B2 => n17655, A => n17654, ZN =>
                           n17660);
   U1708 : INV_X1 port map( A => n17656, ZN => n17658);
   U1709 : AOI211_X1 port map( C1 => n17660, C2 => n17659, A => n17658, B => 
                           n17657, ZN => n17666);
   U1710 : NAND2_X1 port map( A1 => n17662, A2 => n17661, ZN => n17665);
   U1711 : OAI211_X1 port map( C1 => n17666, C2 => n17665, A => n17664, B => 
                           n17663, ZN => n17668);
   U1712 : OAI211_X1 port map( C1 => DATA1(18), C2 => n17783, A => n17668, B =>
                           n17667, ZN => n17670);
   U1713 : AOI21_X1 port map( B1 => n17671, B2 => n17670, A => n17669, ZN => 
                           n17673);
   U1714 : OAI21_X1 port map( B1 => n17674, B2 => n17673, A => n17672, ZN => 
                           n17676);
   U1715 : AOI22_X1 port map( A1 => n17677, A2 => n17676, B1 => DATA2(22), B2 
                           => n17675, ZN => n17681);
   U1716 : AOI211_X1 port map( C1 => n17681, C2 => n17680, A => n17679, B => 
                           n17678, ZN => n17682);
   U1717 : AOI21_X1 port map( B1 => DATA2(24), B2 => n17683, A => n17682, ZN =>
                           n17687);
   U1718 : AOI211_X1 port map( C1 => n17687, C2 => n17686, A => n17685, B => 
                           n17684, ZN => n17688);
   U1719 : AOI21_X1 port map( B1 => DATA2(26), B2 => n17689, A => n17688, ZN =>
                           n17693);
   U1720 : AOI211_X1 port map( C1 => n17693, C2 => n17692, A => n17691, B => 
                           n17690, ZN => n17694);
   U1721 : AOI21_X1 port map( B1 => DATA2(28), B2 => n17695, A => n17694, ZN =>
                           n17699);
   U1722 : AOI211_X1 port map( C1 => n17699, C2 => n17698, A => n17697, B => 
                           n17696, ZN => n17700);
   U1723 : AOI211_X1 port map( C1 => DATA2(30), C2 => n17702, A => n17701, B =>
                           n17700, ZN => n17703);
   U1724 : AOI221_X1 port map( B1 => n17704, B2 => n1870, C1 => n17703, C2 => 
                           n1870, A => FUNC(2), ZN => n17705);
   U1725 : OAI221_X1 port map( B1 => n1870, B2 => n17707, C1 => n1870, C2 => 
                           n17706, A => n17705, ZN => n12750);
   U1726 : OAI211_X1 port map( C1 => n14438, C2 => n17710, A => n17709, B => 
                           n17708, ZN => n17711);
   U1727 : AOI211_X1 port map( C1 => n17713, C2 => n14461, A => n17712, B => 
                           n17711, ZN => n17719);
   U1728 : INV_X1 port map( A => n17714, ZN => n17717);
   U1729 : OAI222_X1 port map( A1 => n17720, A2 => n17719, B1 => n17718, B2 => 
                           n17717, C1 => n17716, C2 => n17715, ZN => n17721);
   U1730 : AOI22_X1 port map( A1 => n18116, A2 => n17722, B1 => n18159, B2 => 
                           n17721, ZN => n17726);
   U1731 : AOI22_X1 port map( A1 => n18144, A2 => n17724, B1 => n18123, B2 => 
                           n17723, ZN => n17725);
   U1732 : OAI211_X1 port map( C1 => n17727, C2 => n18148, A => n17726, B => 
                           n17725, ZN => n17735);
   U1733 : INV_X1 port map( A => n1861, ZN => n17730);
   U1734 : OAI22_X1 port map( A1 => n17730, A2 => n1896, B1 => n17729, B2 => 
                           n17728, ZN => n17734);
   U1735 : OAI22_X1 port map( A1 => n17732, A2 => n1895, B1 => n17731, B2 => 
                           n9020, ZN => n17733);
   U1736 : AOI211_X1 port map( C1 => n1897, C2 => n17735, A => n17734, B => 
                           n17733, ZN => n12721);
   U1737 : INV_X1 port map( A => n17736, ZN => n17752);
   U1738 : INV_X1 port map( A => n17737, ZN => n17745);
   U1739 : AOI22_X1 port map( A1 => n14221, A2 => n17739, B1 => n18176, B2 => 
                           n17738, ZN => n17744);
   U1740 : OAI222_X1 port map( A1 => n14228, A2 => n13921, B1 => n14373, B2 => 
                           n17740, C1 => n14390, C2 => n13905, ZN => n17742);
   U1741 : AOI22_X1 port map( A1 => n14130, A2 => n17742, B1 => n14384, B2 => 
                           n17741, ZN => n17743);
   U1742 : OAI211_X1 port map( C1 => n17745, C2 => n18182, A => n17744, B => 
                           n17743, ZN => n17747);
   U1743 : AOI22_X1 port map( A1 => n14129, A2 => n17747, B1 => n14388, B2 => 
                           n17746, ZN => n17751);
   U1744 : AOI22_X1 port map( A1 => n13894, A2 => n17749, B1 => n18192, B2 => 
                           n17748, ZN => n17750);
   U1745 : OAI211_X1 port map( C1 => n17752, C2 => n18215, A => n17751, B => 
                           n17750, ZN => n17753);
   U1746 : AOI22_X1 port map( A1 => n14230, A2 => n17754, B1 => n14380, B2 => 
                           n17753, ZN => n17755);
   U1747 : AOI221_X1 port map( B1 => n17756, B2 => n17755, C1 => n18191, C2 => 
                           n17755, A => n14400, ZN => n17762);
   U1748 : AOI22_X1 port map( A1 => n14222, A2 => n17758, B1 => n18207, B2 => 
                           n17757, ZN => n17759);
   U1749 : OAI21_X1 port map( B1 => n14232, B2 => n17760, A => n17759, ZN => 
                           n17761);
   U1750 : AOI211_X1 port map( C1 => n18225, C2 => n17763, A => n17762, B => 
                           n17761, ZN => n17768);
   U1751 : INV_X1 port map( A => n17764, ZN => n17765);
   U1752 : OAI211_X1 port map( C1 => n17765, C2 => n14259, A => n13856, B => 
                           n13908, ZN => n17766);
   U1753 : AOI21_X1 port map( B1 => n13906, B2 => n13907, A => n17766, ZN => 
                           n17767);
   U1754 : OAI21_X1 port map( B1 => n14275, B2 => n17768, A => n17767, ZN => 
                           OUTALU(0));
   U1755 : NAND2_X1 port map( A1 => n17769, A2 => n1870, ZN => n17799);
   U1756 : CLKBUF_X1 port map( A => n17799, Z => n17794);
   U1757 : NAND2_X1 port map( A1 => FUNC(3), A2 => n17769, ZN => n17798);
   U1758 : CLKBUF_X1 port map( A => n17798, Z => n17793);
   U1759 : AOI22_X1 port map( A1 => DATA2(31), A2 => n17794, B1 => n17793, B2 
                           => n17770, ZN => N2548);
   U1760 : AOI22_X1 port map( A1 => DATA2(30), A2 => n17799, B1 => n17798, B2 
                           => n17771, ZN => N2547);
   U1761 : INV_X1 port map( A => DATA2(29), ZN => n17772);
   U1762 : AOI22_X1 port map( A1 => DATA2(29), A2 => n17794, B1 => n17793, B2 
                           => n17772, ZN => N2546);
   U1763 : AOI22_X1 port map( A1 => DATA2(28), A2 => n17799, B1 => n17798, B2 
                           => n17773, ZN => N2545);
   U1764 : INV_X1 port map( A => DATA2(27), ZN => n17774);
   U1765 : AOI22_X1 port map( A1 => DATA2(27), A2 => n17794, B1 => n17793, B2 
                           => n17774, ZN => N2544);
   U1766 : AOI22_X1 port map( A1 => DATA2(26), A2 => n17799, B1 => n17798, B2 
                           => n17775, ZN => N2543);
   U1767 : INV_X1 port map( A => DATA2(25), ZN => n17776);
   U1768 : AOI22_X1 port map( A1 => DATA2(25), A2 => n17794, B1 => n17793, B2 
                           => n17776, ZN => N2542);
   U1769 : AOI22_X1 port map( A1 => DATA2(24), A2 => n17799, B1 => n17798, B2 
                           => n17777, ZN => N2541);
   U1770 : INV_X1 port map( A => DATA2(23), ZN => n17778);
   U1771 : AOI22_X1 port map( A1 => DATA2(23), A2 => n17794, B1 => n17793, B2 
                           => n17778, ZN => N2540);
   U1772 : AOI22_X1 port map( A1 => DATA2(22), A2 => n17799, B1 => n17798, B2 
                           => n17779, ZN => N2539);
   U1773 : AOI22_X1 port map( A1 => DATA2(21), A2 => n17799, B1 => n17798, B2 
                           => n17780, ZN => N2538);
   U1774 : AOI22_X1 port map( A1 => DATA2(20), A2 => n17799, B1 => n17798, B2 
                           => n17781, ZN => N2537);
   U1775 : AOI22_X1 port map( A1 => DATA2(19), A2 => n17794, B1 => n17793, B2 
                           => n17782, ZN => N2536);
   U1776 : AOI22_X1 port map( A1 => DATA2(18), A2 => n17794, B1 => n17793, B2 
                           => n17783, ZN => N2535);
   U1777 : AOI22_X1 port map( A1 => DATA2(17), A2 => n17794, B1 => n17793, B2 
                           => n17784, ZN => N2534);
   U1778 : AOI22_X1 port map( A1 => DATA2(16), A2 => n17794, B1 => n17793, B2 
                           => n17785, ZN => N2533);
   U1779 : INV_X1 port map( A => DATA2(15), ZN => n17786);
   U1780 : AOI22_X1 port map( A1 => DATA2(15), A2 => n17794, B1 => n17793, B2 
                           => n17786, ZN => N2532);
   U1781 : AOI22_X1 port map( A1 => DATA2(14), A2 => n17794, B1 => n17793, B2 
                           => n17787, ZN => N2531);
   U1782 : AOI22_X1 port map( A1 => DATA2(13), A2 => n17794, B1 => n17793, B2 
                           => n17788, ZN => N2530);
   U1783 : AOI22_X1 port map( A1 => DATA2(12), A2 => n17794, B1 => n17793, B2 
                           => n18160, ZN => N2529);
   U1784 : AOI22_X1 port map( A1 => DATA2(11), A2 => n17794, B1 => n17793, B2 
                           => n17789, ZN => N2528);
   U1785 : AOI22_X1 port map( A1 => DATA2(10), A2 => n17794, B1 => n17793, B2 
                           => n17790, ZN => N2527);
   U1786 : AOI22_X1 port map( A1 => DATA2(9), A2 => n17794, B1 => n17793, B2 =>
                           n17791, ZN => N2526);
   U1787 : AOI22_X1 port map( A1 => DATA2(8), A2 => n17794, B1 => n17793, B2 =>
                           n17792, ZN => N2525);
   U1788 : INV_X1 port map( A => DATA2(7), ZN => n17795);
   U1789 : AOI22_X1 port map( A1 => DATA2(7), A2 => n17799, B1 => n17798, B2 =>
                           n17795, ZN => N2524);
   U1790 : AOI22_X1 port map( A1 => DATA2(6), A2 => n17799, B1 => n17798, B2 =>
                           n17796, ZN => N2523);
   U1791 : AOI22_X1 port map( A1 => DATA2(5), A2 => n17799, B1 => n17798, B2 =>
                           n17797, ZN => N2522);
   U1792 : AOI22_X1 port map( A1 => DATA2(4), A2 => n17799, B1 => n17798, B2 =>
                           n18058, ZN => N2521);
   U1793 : AOI22_X1 port map( A1 => DATA2(3), A2 => n17799, B1 => n17798, B2 =>
                           n18082, ZN => N2520);
   U1794 : AOI22_X1 port map( A1 => DATA2(2), A2 => n17799, B1 => n17798, B2 =>
                           n18079, ZN => N2519);
   U1795 : AOI22_X1 port map( A1 => DATA2(1), A2 => n17799, B1 => n17798, B2 =>
                           n18059, ZN => N2518);
   U1796 : AOI22_X1 port map( A1 => DATA2(0), A2 => n17799, B1 => n17798, B2 =>
                           n18062, ZN => N2517);
   U1797 : NOR2_X1 port map( A1 => n17800, A2 => n1844, ZN => n8933);
   U1798 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , ZN => n17801);
   U1799 : NAND2_X1 port map( A1 => n17803, A2 => n17801, ZN => n17835);
   U1800 : NAND2_X1 port map( A1 => n17836, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n17831);
   U1801 : INV_X1 port map( A => n17831, ZN => n17838);
   U1802 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, 
                           ZN => n17802);
   U1803 : NOR2_X1 port map( A1 => n17838, A2 => n17833, ZN => n17804);
   U1804 : NAND2_X1 port map( A1 => n17803, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n17840);
   U1805 : OAI222_X1 port map( A1 => n1843, A2 => n17835, B1 => n1844, B2 => 
                           n17804, C1 => n1842, C2 => n17840, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1806 : OAI22_X1 port map( A1 => n1840, A2 => n17840, B1 => n1842, B2 => 
                           n17831, ZN => n17805);
   U1807 : AOI21_X1 port map( B1 => n17833, B2 => n9084, A => n17805, ZN => 
                           n17806);
   U1808 : OAI21_X1 port map( B1 => n1841, B2 => n17835, A => n17806, ZN => 
                           boothmul_pipelined_i_mux_out_1_4_port);
   U1809 : OAI22_X1 port map( A1 => n1840, A2 => n17831, B1 => n17840, B2 => 
                           n1838, ZN => n17807);
   U1810 : AOI21_X1 port map( B1 => n9081, B2 => n17833, A => n17807, ZN => 
                           n17808);
   U1811 : OAI21_X1 port map( B1 => n17835, B2 => n1839, A => n17808, ZN => 
                           boothmul_pipelined_i_mux_out_1_5_port);
   U1812 : OAI22_X1 port map( A1 => n17840, A2 => n1836, B1 => n17831, B2 => 
                           n1838, ZN => n17809);
   U1813 : AOI21_X1 port map( B1 => n17833, B2 => n9078, A => n17809, ZN => 
                           n17810);
   U1814 : OAI21_X1 port map( B1 => n17835, B2 => n1837, A => n17810, ZN => 
                           boothmul_pipelined_i_mux_out_1_6_port);
   U1815 : OAI22_X1 port map( A1 => n17840, A2 => n1833, B1 => n17831, B2 => 
                           n1836, ZN => n17811);
   U1816 : AOI21_X1 port map( B1 => n17833, B2 => n9075, A => n17811, ZN => 
                           n17812);
   U1817 : OAI21_X1 port map( B1 => n17835, B2 => n1834, A => n17812, ZN => 
                           boothmul_pipelined_i_mux_out_1_7_port);
   U1818 : OAI22_X1 port map( A1 => n17840, A2 => n1831, B1 => n17831, B2 => 
                           n1833, ZN => n17813);
   U1819 : AOI21_X1 port map( B1 => n17833, B2 => n9072, A => n17813, ZN => 
                           n17814);
   U1820 : OAI21_X1 port map( B1 => n17835, B2 => n1832, A => n17814, ZN => 
                           boothmul_pipelined_i_mux_out_1_8_port);
   U1821 : OAI22_X1 port map( A1 => n17840, A2 => n1829, B1 => n17831, B2 => 
                           n1831, ZN => n17815);
   U1822 : AOI21_X1 port map( B1 => n17833, B2 => n9069, A => n17815, ZN => 
                           n17816);
   U1823 : OAI21_X1 port map( B1 => n17835, B2 => n1830, A => n17816, ZN => 
                           boothmul_pipelined_i_mux_out_1_9_port);
   U1824 : OAI22_X1 port map( A1 => n17840, A2 => n1827, B1 => n17831, B2 => 
                           n1829, ZN => n17817);
   U1825 : AOI21_X1 port map( B1 => n17833, B2 => n9066, A => n17817, ZN => 
                           n17818);
   U1826 : OAI21_X1 port map( B1 => n17835, B2 => n1828, A => n17818, ZN => 
                           boothmul_pipelined_i_mux_out_1_10_port);
   U1827 : OAI22_X1 port map( A1 => n17840, A2 => n1825, B1 => n17831, B2 => 
                           n1827, ZN => n17819);
   U1828 : AOI21_X1 port map( B1 => n17833, B2 => n9063, A => n17819, ZN => 
                           n17820);
   U1829 : OAI21_X1 port map( B1 => n17835, B2 => n1826, A => n17820, ZN => 
                           boothmul_pipelined_i_mux_out_1_11_port);
   U1830 : OAI22_X1 port map( A1 => n17840, A2 => n1823, B1 => n17831, B2 => 
                           n1825, ZN => n17821);
   U1831 : AOI21_X1 port map( B1 => n17833, B2 => n9060, A => n17821, ZN => 
                           n17822);
   U1832 : OAI21_X1 port map( B1 => n17835, B2 => n1824, A => n17822, ZN => 
                           boothmul_pipelined_i_mux_out_1_12_port);
   U1833 : OAI22_X1 port map( A1 => n17840, A2 => n1821, B1 => n17831, B2 => 
                           n1823, ZN => n17823);
   U1834 : AOI21_X1 port map( B1 => n17833, B2 => n9057, A => n17823, ZN => 
                           n17824);
   U1835 : OAI21_X1 port map( B1 => n17835, B2 => n1822, A => n17824, ZN => 
                           boothmul_pipelined_i_mux_out_1_13_port);
   U1836 : OAI22_X1 port map( A1 => n17840, A2 => n1819, B1 => n17831, B2 => 
                           n1821, ZN => n17825);
   U1837 : AOI21_X1 port map( B1 => n17833, B2 => n9054, A => n17825, ZN => 
                           n17826);
   U1838 : OAI21_X1 port map( B1 => n17835, B2 => n1820, A => n17826, ZN => 
                           boothmul_pipelined_i_mux_out_1_14_port);
   U1839 : OAI22_X1 port map( A1 => n17840, A2 => n1817, B1 => n17831, B2 => 
                           n1819, ZN => n17827);
   U1840 : AOI21_X1 port map( B1 => n17833, B2 => n9051, A => n17827, ZN => 
                           n17828);
   U1841 : OAI21_X1 port map( B1 => n17835, B2 => n1818, A => n17828, ZN => 
                           boothmul_pipelined_i_mux_out_1_15_port);
   U1842 : OAI22_X1 port map( A1 => n17840, A2 => n1815, B1 => n17831, B2 => 
                           n1817, ZN => n17829);
   U1843 : AOI21_X1 port map( B1 => n17833, B2 => n9048, A => n17829, ZN => 
                           n17830);
   U1844 : OAI21_X1 port map( B1 => n17835, B2 => n1816, A => n17830, ZN => 
                           boothmul_pipelined_i_mux_out_1_16_port);
   U1845 : OAI22_X1 port map( A1 => n17840, A2 => n1813, B1 => n17831, B2 => 
                           n1815, ZN => n17832);
   U1846 : AOI21_X1 port map( B1 => n17833, B2 => n9045, A => n17832, ZN => 
                           n17834);
   U1847 : OAI21_X1 port map( B1 => n17835, B2 => n1814, A => n17834, ZN => 
                           boothmul_pipelined_i_mux_out_1_17_port);
   U1848 : NOR3_X1 port map( A1 => n17836, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A3 
                           => n1814, ZN => n17837);
   U1849 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           B2 => n17838, A => n17837, ZN => n17839);
   U1850 : OAI21_X1 port map( B1 => n1812, B2 => n17840, A => n17839, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1851 : OR2_X1 port map( A1 => n17841, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n8932);
   U1852 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n14223, B1 => n9084, B2 => n14182, ZN => 
                           n17842);
   U1853 : OAI221_X1 port map( B1 => n1844, B2 => n14224, C1 => n1844, C2 => 
                           n14252, A => n17842, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1854 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n14223, B1 => n9081, B2 => n14182, ZN => 
                           n17844);
   U1855 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n14399, ZN => n17843);
   U1856 : OAI211_X1 port map( C1 => n14252, C2 => n1843, A => n17844, B => 
                           n17843, ZN => boothmul_pipelined_i_mux_out_2_6_port)
                           ;
   U1857 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n14223, ZN => n17846);
   U1858 : NAND2_X1 port map( A1 => n9078, A2 => n14182, ZN => n17845);
   U1859 : OAI211_X1 port map( C1 => n14252, C2 => n1841, A => n17846, B => 
                           n17845, ZN => boothmul_pipelined_i_mux_out_2_7_port)
                           ;
   U1860 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n14223, ZN => n17848);
   U1861 : NAND2_X1 port map( A1 => n9075, A2 => n14182, ZN => n17847);
   U1862 : OAI211_X1 port map( C1 => n14252, C2 => n1839, A => n17848, B => 
                           n17847, ZN => boothmul_pipelined_i_mux_out_2_8_port)
                           ;
   U1863 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n14223, ZN => n17850);
   U1864 : NAND2_X1 port map( A1 => n9072, A2 => n14182, ZN => n17849);
   U1865 : OAI211_X1 port map( C1 => n14252, C2 => n1837, A => n17850, B => 
                           n17849, ZN => boothmul_pipelined_i_mux_out_2_9_port)
                           ;
   U1866 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n14223, ZN => n17852);
   U1867 : NAND2_X1 port map( A1 => n9069, A2 => n14182, ZN => n17851);
   U1868 : OAI211_X1 port map( C1 => n14252, C2 => n1834, A => n17852, B => 
                           n17851, ZN => boothmul_pipelined_i_mux_out_2_10_port
                           );
   U1869 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n14223, ZN => n17854);
   U1870 : NAND2_X1 port map( A1 => n9066, A2 => n14182, ZN => n17853);
   U1871 : OAI211_X1 port map( C1 => n14252, C2 => n1832, A => n17854, B => 
                           n17853, ZN => boothmul_pipelined_i_mux_out_2_11_port
                           );
   U1872 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n14223, ZN => n17856);
   U1873 : NAND2_X1 port map( A1 => n9063, A2 => n14182, ZN => n17855);
   U1874 : OAI211_X1 port map( C1 => n14252, C2 => n1830, A => n17856, B => 
                           n17855, ZN => boothmul_pipelined_i_mux_out_2_12_port
                           );
   U1875 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n14223, ZN => n17858);
   U1876 : NAND2_X1 port map( A1 => n9060, A2 => n14182, ZN => n17857);
   U1877 : OAI211_X1 port map( C1 => n14252, C2 => n1828, A => n17858, B => 
                           n17857, ZN => boothmul_pipelined_i_mux_out_2_13_port
                           );
   U1878 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n14223, ZN => n17860);
   U1879 : NAND2_X1 port map( A1 => n9057, A2 => n14182, ZN => n17859);
   U1880 : OAI211_X1 port map( C1 => n14252, C2 => n1826, A => n17860, B => 
                           n17859, ZN => boothmul_pipelined_i_mux_out_2_14_port
                           );
   U1881 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n14223, ZN => n17862);
   U1882 : NAND2_X1 port map( A1 => n9054, A2 => n14182, ZN => n17861);
   U1883 : OAI211_X1 port map( C1 => n14252, C2 => n1824, A => n17862, B => 
                           n17861, ZN => boothmul_pipelined_i_mux_out_2_15_port
                           );
   U1884 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n14223, ZN => n17864);
   U1885 : NAND2_X1 port map( A1 => n9051, A2 => n14182, ZN => n17863);
   U1886 : OAI211_X1 port map( C1 => n14252, C2 => n1822, A => n17864, B => 
                           n17863, ZN => boothmul_pipelined_i_mux_out_2_16_port
                           );
   U1887 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n14223, ZN => n17866);
   U1888 : NAND2_X1 port map( A1 => n9048, A2 => n14182, ZN => n17865);
   U1889 : OAI211_X1 port map( C1 => n14252, C2 => n1820, A => n17866, B => 
                           n17865, ZN => boothmul_pipelined_i_mux_out_2_17_port
                           );
   U1890 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n14223, ZN => n17868);
   U1891 : NAND2_X1 port map( A1 => n9045, A2 => n14182, ZN => n17867);
   U1892 : OAI211_X1 port map( C1 => n14252, C2 => n1818, A => n17868, B => 
                           n17867, ZN => boothmul_pipelined_i_mux_out_2_18_port
                           );
   U1893 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n14399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n14223, ZN => n17870);
   U1894 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n14182, ZN => 
                           n17869);
   U1895 : OAI211_X1 port map( C1 => n14252, C2 => n1816, A => n17870, B => 
                           n17869, ZN => boothmul_pipelined_i_mux_out_2_19_port
                           );
   U1896 : OAI222_X1 port map( A1 => n1813, A2 => n14224, B1 => n1814, B2 => 
                           n14183, C1 => n14372, C2 => n1812, ZN => n8535);
   U1897 : NAND2_X1 port map( A1 => n7769, A2 => n17871, ZN => n8931);
   U1898 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n14419, B1 => n9084, B2 => n14379, ZN => 
                           n17872);
   U1899 : OAI221_X1 port map( B1 => n1844, B2 => n14251, C1 => n1844, C2 => 
                           n14282, A => n17872, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1900 : OAI22_X1 port map( A1 => n14282, A2 => n1843, B1 => n14283, B2 => 
                           n1841, ZN => n17873);
   U1901 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           B2 => n14419, A => n17873, ZN => n17874);
   U1902 : OAI21_X1 port map( B1 => n14251, B2 => n1842, A => n17874, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1903 : OAI22_X1 port map( A1 => n14251, A2 => n1840, B1 => n14283, B2 => 
                           n1839, ZN => n17875);
   U1904 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           B2 => n14419, A => n17875, ZN => n17876);
   U1905 : OAI21_X1 port map( B1 => n14282, B2 => n1841, A => n17876, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1906 : OAI22_X1 port map( A1 => n14251, A2 => n1838, B1 => n14283, B2 => 
                           n1837, ZN => n17877);
   U1907 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           B2 => n14419, A => n17877, ZN => n17878);
   U1908 : OAI21_X1 port map( B1 => n14282, B2 => n1839, A => n17878, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1909 : OAI22_X1 port map( A1 => n14251, A2 => n1836, B1 => n14283, B2 => 
                           n1834, ZN => n17879);
   U1910 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           B2 => n14419, A => n17879, ZN => n17880);
   U1911 : OAI21_X1 port map( B1 => n14282, B2 => n1837, A => n17880, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1912 : OAI22_X1 port map( A1 => n14251, A2 => n1833, B1 => n14283, B2 => 
                           n1832, ZN => n17881);
   U1913 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           B2 => n14419, A => n17881, ZN => n17882);
   U1914 : OAI21_X1 port map( B1 => n14282, B2 => n1834, A => n17882, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1915 : OAI22_X1 port map( A1 => n14251, A2 => n1831, B1 => n14283, B2 => 
                           n1830, ZN => n17883);
   U1916 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           B2 => n14419, A => n17883, ZN => n17884);
   U1917 : OAI21_X1 port map( B1 => n14282, B2 => n1832, A => n17884, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1918 : OAI22_X1 port map( A1 => n14251, A2 => n1829, B1 => n14283, B2 => 
                           n1828, ZN => n17885);
   U1919 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           B2 => n14419, A => n17885, ZN => n17886);
   U1920 : OAI21_X1 port map( B1 => n14282, B2 => n1830, A => n17886, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U1921 : OAI22_X1 port map( A1 => n14251, A2 => n1827, B1 => n14283, B2 => 
                           n1826, ZN => n17887);
   U1922 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           B2 => n14419, A => n17887, ZN => n17888);
   U1923 : OAI21_X1 port map( B1 => n14282, B2 => n1828, A => n17888, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U1924 : OAI22_X1 port map( A1 => n14251, A2 => n1825, B1 => n14283, B2 => 
                           n1824, ZN => n17889);
   U1925 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           B2 => n14419, A => n17889, ZN => n17890);
   U1926 : OAI21_X1 port map( B1 => n14282, B2 => n1826, A => n17890, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U1927 : OAI22_X1 port map( A1 => n14251, A2 => n1823, B1 => n14283, B2 => 
                           n1822, ZN => n17891);
   U1928 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           B2 => n14419, A => n17891, ZN => n17892);
   U1929 : OAI21_X1 port map( B1 => n14282, B2 => n1824, A => n17892, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U1930 : OAI22_X1 port map( A1 => n14251, A2 => n1821, B1 => n14283, B2 => 
                           n1820, ZN => n17893);
   U1931 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           B2 => n14419, A => n17893, ZN => n17894);
   U1932 : OAI21_X1 port map( B1 => n14282, B2 => n1822, A => n17894, ZN => 
                           n8813);
   U1933 : OAI22_X1 port map( A1 => n14251, A2 => n1819, B1 => n14283, B2 => 
                           n1818, ZN => n17895);
   U1934 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           B2 => n14419, A => n17895, ZN => n17896);
   U1935 : OAI21_X1 port map( B1 => n14282, B2 => n1820, A => n17896, ZN => 
                           n8812);
   U1936 : OAI22_X1 port map( A1 => n14251, A2 => n1817, B1 => n14283, B2 => 
                           n1816, ZN => n17897);
   U1937 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           B2 => n14419, A => n17897, ZN => n17898);
   U1938 : OAI21_X1 port map( B1 => n14282, B2 => n1818, A => n17898, ZN => 
                           n8811);
   U1939 : OAI22_X1 port map( A1 => n14251, A2 => n1815, B1 => n14283, B2 => 
                           n1814, ZN => n17899);
   U1940 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           B2 => n14419, A => n17899, ZN => n17900);
   U1941 : OAI21_X1 port map( B1 => n14282, B2 => n1816, A => n17900, ZN => 
                           n8810);
   U1942 : OAI222_X1 port map( A1 => n1813, A2 => n14251, B1 => n1814, B2 => 
                           n14281, C1 => n14233, C2 => n1812, ZN => n8534);
   U1943 : NAND3_X1 port map( A1 => n7769, A2 => n8978, A3 => n1845, ZN => 
                           n12927);
   U1944 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n14285, B1 => n9084, B2 => n14421, ZN => 
                           n17901);
   U1945 : OAI221_X1 port map( B1 => n1844, B2 => n14141, C1 => n1844, C2 => 
                           n14422, A => n17901, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U1946 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n14285, B1 => n9081, B2 => n14421, ZN => 
                           n17903);
   U1947 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n14284, ZN => n17902);
   U1948 : OAI211_X1 port map( C1 => n14141, C2 => n1843, A => n17903, B => 
                           n17902, ZN => boothmul_pipelined_i_mux_out_4_10_port
                           );
   U1949 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n14285, ZN => n17905);
   U1950 : NAND2_X1 port map( A1 => n9078, A2 => n14421, ZN => n17904);
   U1951 : OAI211_X1 port map( C1 => n14141, C2 => n1841, A => n17905, B => 
                           n17904, ZN => boothmul_pipelined_i_mux_out_4_11_port
                           );
   U1952 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n14285, ZN => n17907);
   U1953 : NAND2_X1 port map( A1 => n9075, A2 => n14421, ZN => n17906);
   U1954 : OAI211_X1 port map( C1 => n14141, C2 => n1839, A => n17907, B => 
                           n17906, ZN => boothmul_pipelined_i_mux_out_4_12_port
                           );
   U1955 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n14285, ZN => n17909);
   U1956 : NAND2_X1 port map( A1 => n9072, A2 => n14421, ZN => n17908);
   U1957 : OAI211_X1 port map( C1 => n14141, C2 => n1837, A => n17909, B => 
                           n17908, ZN => boothmul_pipelined_i_mux_out_4_13_port
                           );
   U1958 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n14285, ZN => n17911);
   U1959 : NAND2_X1 port map( A1 => n9069, A2 => n14421, ZN => n17910);
   U1960 : OAI211_X1 port map( C1 => n14141, C2 => n1834, A => n17911, B => 
                           n17910, ZN => boothmul_pipelined_i_mux_out_4_14_port
                           );
   U1961 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n14285, ZN => n17913);
   U1962 : NAND2_X1 port map( A1 => n9066, A2 => n14421, ZN => n17912);
   U1963 : OAI211_X1 port map( C1 => n14141, C2 => n1832, A => n17913, B => 
                           n17912, ZN => boothmul_pipelined_i_mux_out_4_15_port
                           );
   U1964 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n14285, ZN => n17915);
   U1965 : NAND2_X1 port map( A1 => n9063, A2 => n14421, ZN => n17914);
   U1966 : OAI211_X1 port map( C1 => n14141, C2 => n1830, A => n17915, B => 
                           n17914, ZN => n8928);
   U1967 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n14285, ZN => n17917);
   U1968 : NAND2_X1 port map( A1 => n9060, A2 => n14421, ZN => n17916);
   U1969 : OAI211_X1 port map( C1 => n14141, C2 => n1828, A => n17917, B => 
                           n17916, ZN => n8927);
   U1970 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n14285, ZN => n17919);
   U1971 : NAND2_X1 port map( A1 => n9057, A2 => n14421, ZN => n17918);
   U1972 : OAI211_X1 port map( C1 => n14141, C2 => n1826, A => n17919, B => 
                           n17918, ZN => n8926);
   U1973 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n14285, ZN => n17921);
   U1974 : NAND2_X1 port map( A1 => n9054, A2 => n14421, ZN => n17920);
   U1975 : OAI211_X1 port map( C1 => n14141, C2 => n1824, A => n17921, B => 
                           n17920, ZN => n8925);
   U1976 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n14285, ZN => n17923);
   U1977 : NAND2_X1 port map( A1 => n9051, A2 => n14421, ZN => n17922);
   U1978 : OAI211_X1 port map( C1 => n14141, C2 => n1822, A => n17923, B => 
                           n17922, ZN => n8924);
   U1979 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n14285, ZN => n17925);
   U1980 : NAND2_X1 port map( A1 => n9048, A2 => n14421, ZN => n17924);
   U1981 : OAI211_X1 port map( C1 => n14141, C2 => n1820, A => n17925, B => 
                           n17924, ZN => n8923);
   U1982 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n14285, ZN => n17927);
   U1983 : NAND2_X1 port map( A1 => n9045, A2 => n14421, ZN => n17926);
   U1984 : OAI211_X1 port map( C1 => n14141, C2 => n1818, A => n17927, B => 
                           n17926, ZN => n8922);
   U1985 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n14284, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n14285, ZN => n17929);
   U1986 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n14421, ZN => 
                           n17928);
   U1987 : OAI211_X1 port map( C1 => n14141, C2 => n1816, A => n17929, B => 
                           n17928, ZN => n8921);
   U1988 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n14284, B1 => n14285, B2 => n18051, ZN => 
                           n17930);
   U1989 : OAI221_X1 port map( B1 => n1814, B2 => n14141, C1 => n1814, C2 => 
                           n14250, A => n17930, ZN => n8549);
   U1990 : NAND3_X1 port map( A1 => n14286, A2 => n16410, A3 => n16391, ZN => 
                           n17963);
   U1991 : NOR2_X1 port map( A1 => n16410, A2 => n14286, ZN => n17931);
   U1992 : NAND2_X1 port map( A1 => n17931, A2 => n14287, ZN => n17968);
   U1993 : NOR2_X1 port map( A1 => n17932, A2 => n16391, ZN => n17934);
   U1994 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n17934, B1 => n9084, B2 => n17965, ZN => 
                           n17933);
   U1995 : OAI221_X1 port map( B1 => n1844, B2 => n17963, C1 => n1844, C2 => 
                           n17968, A => n17933, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U1996 : INV_X1 port map( A => n17934, ZN => n17967);
   U1997 : OAI22_X1 port map( A1 => n1842, A2 => n17968, B1 => n1843, B2 => 
                           n17963, ZN => n17935);
   U1998 : AOI21_X1 port map( B1 => n9081, B2 => n17965, A => n17935, ZN => 
                           n17936);
   U1999 : OAI21_X1 port map( B1 => n1840, B2 => n17967, A => n17936, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2000 : OAI22_X1 port map( A1 => n1840, A2 => n17968, B1 => n1841, B2 => 
                           n17963, ZN => n17937);
   U2001 : AOI21_X1 port map( B1 => n9078, B2 => n17965, A => n17937, ZN => 
                           n17938);
   U2002 : OAI21_X1 port map( B1 => n1838, B2 => n17967, A => n17938, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2003 : OAI22_X1 port map( A1 => n1839, A2 => n17963, B1 => n1838, B2 => 
                           n17968, ZN => n17939);
   U2004 : AOI21_X1 port map( B1 => n9075, B2 => n17965, A => n17939, ZN => 
                           n17940);
   U2005 : OAI21_X1 port map( B1 => n1836, B2 => n17967, A => n17940, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2006 : OAI22_X1 port map( A1 => n1837, A2 => n17963, B1 => n1836, B2 => 
                           n17968, ZN => n17941);
   U2007 : AOI21_X1 port map( B1 => n9072, B2 => n17965, A => n17941, ZN => 
                           n17942);
   U2008 : OAI21_X1 port map( B1 => n1833, B2 => n17967, A => n17942, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2009 : OAI22_X1 port map( A1 => n1834, A2 => n17963, B1 => n1833, B2 => 
                           n17968, ZN => n17943);
   U2010 : AOI21_X1 port map( B1 => n9069, B2 => n17965, A => n17943, ZN => 
                           n17944);
   U2011 : OAI21_X1 port map( B1 => n1831, B2 => n17967, A => n17944, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2012 : OAI22_X1 port map( A1 => n1832, A2 => n17963, B1 => n1831, B2 => 
                           n17968, ZN => n17945);
   U2013 : AOI21_X1 port map( B1 => n9066, B2 => n17965, A => n17945, ZN => 
                           n17946);
   U2014 : OAI21_X1 port map( B1 => n1829, B2 => n17967, A => n17946, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2015 : OAI22_X1 port map( A1 => n1830, A2 => n17963, B1 => n1829, B2 => 
                           n17968, ZN => n17947);
   U2016 : AOI21_X1 port map( B1 => n9063, B2 => n17965, A => n17947, ZN => 
                           n17948);
   U2017 : OAI21_X1 port map( B1 => n1827, B2 => n17967, A => n17948, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2018 : OAI22_X1 port map( A1 => n1828, A2 => n17963, B1 => n1827, B2 => 
                           n17968, ZN => n17949);
   U2019 : AOI21_X1 port map( B1 => n9060, B2 => n17965, A => n17949, ZN => 
                           n17950);
   U2020 : OAI21_X1 port map( B1 => n1825, B2 => n17967, A => n17950, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2021 : OAI22_X1 port map( A1 => n1826, A2 => n17963, B1 => n1825, B2 => 
                           n17968, ZN => n17951);
   U2022 : AOI21_X1 port map( B1 => n9057, B2 => n17965, A => n17951, ZN => 
                           n17952);
   U2023 : OAI21_X1 port map( B1 => n1823, B2 => n17967, A => n17952, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2024 : OAI22_X1 port map( A1 => n1824, A2 => n17963, B1 => n1823, B2 => 
                           n17968, ZN => n17953);
   U2025 : AOI21_X1 port map( B1 => n9054, B2 => n17965, A => n17953, ZN => 
                           n17954);
   U2026 : OAI21_X1 port map( B1 => n1821, B2 => n17967, A => n17954, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2027 : OAI22_X1 port map( A1 => n1822, A2 => n17963, B1 => n1821, B2 => 
                           n17968, ZN => n17955);
   U2028 : AOI21_X1 port map( B1 => n9051, B2 => n17965, A => n17955, ZN => 
                           n17956);
   U2029 : OAI21_X1 port map( B1 => n1819, B2 => n17967, A => n17956, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2030 : OAI22_X1 port map( A1 => n1820, A2 => n17963, B1 => n1819, B2 => 
                           n17968, ZN => n17957);
   U2031 : AOI21_X1 port map( B1 => n9048, B2 => n17965, A => n17957, ZN => 
                           n17958);
   U2032 : OAI21_X1 port map( B1 => n1817, B2 => n17967, A => n17958, ZN => 
                           n8920);
   U2033 : OAI22_X1 port map( A1 => n1818, A2 => n17963, B1 => n1817, B2 => 
                           n17968, ZN => n17959);
   U2034 : AOI21_X1 port map( B1 => n9045, B2 => n17965, A => n17959, ZN => 
                           n17960);
   U2035 : OAI21_X1 port map( B1 => n1815, B2 => n17967, A => n17960, ZN => 
                           n8919);
   U2036 : OAI22_X1 port map( A1 => n1816, A2 => n17963, B1 => n1815, B2 => 
                           n17968, ZN => n17961);
   U2037 : AOI21_X1 port map( B1 => data1_mul_15_port, B2 => n17965, A => 
                           n17961, ZN => n17962);
   U2038 : OAI21_X1 port map( B1 => n1813, B2 => n17967, A => n17962, ZN => 
                           n8918);
   U2039 : INV_X1 port map( A => n17963, ZN => n17964);
   U2040 : NOR2_X1 port map( A1 => n17965, A2 => n17964, ZN => n17966);
   U2041 : OAI222_X1 port map( A1 => n17968, A2 => n1813, B1 => n17967, B2 => 
                           n1812, C1 => n1814, C2 => n17966, ZN => n8548);
   U2042 : NAND3_X1 port map( A1 => n14288, A2 => n16396, A3 => n16390, ZN => 
                           n18006);
   U2043 : NOR2_X1 port map( A1 => n16396, A2 => n14288, ZN => n17969);
   U2044 : NAND2_X1 port map( A1 => n17969, A2 => n14290, ZN => n17972);
   U2045 : AOI22_X1 port map( A1 => n17999, A2 => n14299, B1 => n18003, B2 => 
                           n14219, ZN => n17971);
   U2046 : OAI221_X1 port map( B1 => n14353, B2 => n18006, C1 => n14353, C2 => 
                           n17972, A => n17971, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2047 : INV_X1 port map( A => n18006, ZN => n18000);
   U2048 : INV_X1 port map( A => n17972, ZN => n18004);
   U2049 : AOI22_X1 port map( A1 => n14299, A2 => n18000, B1 => n18004, B2 => 
                           n14219, ZN => n17974);
   U2050 : AOI22_X1 port map( A1 => n17999, A2 => n14301, B1 => n18003, B2 => 
                           n14217, ZN => n17973);
   U2051 : NAND2_X1 port map( A1 => n17974, A2 => n17973, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2052 : AOI22_X1 port map( A1 => n18000, A2 => n14301, B1 => n18004, B2 => 
                           n14217, ZN => n17976);
   U2053 : AOI22_X1 port map( A1 => n17999, A2 => n14303, B1 => n18003, B2 => 
                           n14215, ZN => n17975);
   U2054 : NAND2_X1 port map( A1 => n17976, A2 => n17975, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2055 : AOI22_X1 port map( A1 => n18000, A2 => n14303, B1 => n18004, B2 => 
                           n14215, ZN => n17978);
   U2056 : AOI22_X1 port map( A1 => n17999, A2 => n14305, B1 => n18003, B2 => 
                           n14213, ZN => n17977);
   U2057 : NAND2_X1 port map( A1 => n17978, A2 => n17977, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2058 : AOI22_X1 port map( A1 => n18000, A2 => n14305, B1 => n18004, B2 => 
                           n14213, ZN => n17980);
   U2059 : AOI22_X1 port map( A1 => n17999, A2 => n14307, B1 => n18003, B2 => 
                           n14211, ZN => n17979);
   U2060 : NAND2_X1 port map( A1 => n17980, A2 => n17979, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2061 : AOI22_X1 port map( A1 => n18000, A2 => n14307, B1 => n18004, B2 => 
                           n14211, ZN => n17982);
   U2062 : AOI22_X1 port map( A1 => n17999, A2 => n14309, B1 => n18003, B2 => 
                           n14209, ZN => n17981);
   U2063 : NAND2_X1 port map( A1 => n17982, A2 => n17981, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2064 : AOI22_X1 port map( A1 => n18000, A2 => n14309, B1 => n18004, B2 => 
                           n14209, ZN => n17984);
   U2065 : AOI22_X1 port map( A1 => n17999, A2 => n14311, B1 => n18003, B2 => 
                           n14207, ZN => n17983);
   U2066 : NAND2_X1 port map( A1 => n17984, A2 => n17983, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2067 : AOI22_X1 port map( A1 => n18000, A2 => n14311, B1 => n18004, B2 => 
                           n14207, ZN => n17986);
   U2068 : AOI22_X1 port map( A1 => n17999, A2 => n14313, B1 => n18003, B2 => 
                           n14205, ZN => n17985);
   U2069 : NAND2_X1 port map( A1 => n17986, A2 => n17985, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2070 : AOI22_X1 port map( A1 => n18000, A2 => n14313, B1 => n18004, B2 => 
                           n14205, ZN => n17988);
   U2071 : AOI22_X1 port map( A1 => n17999, A2 => n14315, B1 => n18003, B2 => 
                           n14203, ZN => n17987);
   U2072 : NAND2_X1 port map( A1 => n17988, A2 => n17987, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2073 : AOI22_X1 port map( A1 => n18000, A2 => n14315, B1 => n18004, B2 => 
                           n14203, ZN => n17990);
   U2074 : AOI22_X1 port map( A1 => n17999, A2 => n14317, B1 => n18003, B2 => 
                           n14201, ZN => n17989);
   U2075 : NAND2_X1 port map( A1 => n17990, A2 => n17989, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2076 : AOI22_X1 port map( A1 => n18000, A2 => n14317, B1 => n18004, B2 => 
                           n14201, ZN => n17992);
   U2077 : AOI22_X1 port map( A1 => n17999, A2 => n14319, B1 => n18003, B2 => 
                           n14199, ZN => n17991);
   U2078 : NAND2_X1 port map( A1 => n17992, A2 => n17991, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2079 : AOI22_X1 port map( A1 => n18000, A2 => n14319, B1 => n18004, B2 => 
                           n14199, ZN => n17994);
   U2080 : AOI22_X1 port map( A1 => n17999, A2 => n14321, B1 => n18003, B2 => 
                           n14197, ZN => n17993);
   U2081 : NAND2_X1 port map( A1 => n17994, A2 => n17993, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2082 : AOI22_X1 port map( A1 => n18000, A2 => n14321, B1 => n18004, B2 => 
                           n14197, ZN => n17996);
   U2083 : AOI22_X1 port map( A1 => n17999, A2 => n14323, B1 => n18003, B2 => 
                           n14195, ZN => n17995);
   U2084 : NAND2_X1 port map( A1 => n17996, A2 => n17995, ZN => n8917);
   U2085 : AOI22_X1 port map( A1 => n18000, A2 => n14323, B1 => n18004, B2 => 
                           n14195, ZN => n17998);
   U2086 : AOI22_X1 port map( A1 => n17999, A2 => n14325, B1 => n18003, B2 => 
                           n14193, ZN => n17997);
   U2087 : NAND2_X1 port map( A1 => n17998, A2 => n17997, ZN => n8916);
   U2088 : INV_X1 port map( A => n17999, ZN => n18007);
   U2089 : AOI22_X1 port map( A1 => n18000, A2 => n14325, B1 => n18004, B2 => 
                           n14193, ZN => n18002);
   U2090 : NAND2_X1 port map( A1 => n18003, A2 => n14191, ZN => n18001);
   U2091 : OAI211_X1 port map( C1 => n14355, C2 => n18007, A => n18002, B => 
                           n18001, ZN => n8915);
   U2092 : AOI22_X1 port map( A1 => n18004, A2 => n14191, B1 => n18003, B2 => 
                           n14280, ZN => n18005);
   U2093 : OAI221_X1 port map( B1 => n14355, B2 => n18007, C1 => n14355, C2 => 
                           n18006, A => n18005, ZN => n8547);
   U2094 : NAND3_X1 port map( A1 => n16389, A2 => n14292, A3 => n16394, ZN => 
                           n18011);
   U2095 : INV_X1 port map( A => n18043, ZN => n18010);
   U2096 : AOI22_X1 port map( A1 => n18041, A2 => n14298, B1 => n18042, B2 => 
                           n14218, ZN => n18009);
   U2097 : OAI221_X1 port map( B1 => n14352, B2 => n18011, C1 => n14352, C2 => 
                           n18010, A => n18009, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2098 : INV_X1 port map( A => n18011, ZN => n18040);
   U2099 : AOI22_X1 port map( A1 => n14298, A2 => n18040, B1 => n18043, B2 => 
                           n14218, ZN => n18013);
   U2100 : AOI22_X1 port map( A1 => n18041, A2 => n14300, B1 => n18042, B2 => 
                           n14216, ZN => n18012);
   U2101 : NAND2_X1 port map( A1 => n18013, A2 => n18012, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2102 : AOI22_X1 port map( A1 => n18040, A2 => n14300, B1 => n18043, B2 => 
                           n14216, ZN => n18015);
   U2103 : AOI22_X1 port map( A1 => n18041, A2 => n14302, B1 => n18042, B2 => 
                           n14214, ZN => n18014);
   U2104 : NAND2_X1 port map( A1 => n18015, A2 => n18014, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2105 : AOI22_X1 port map( A1 => n18040, A2 => n14302, B1 => n18043, B2 => 
                           n14214, ZN => n18017);
   U2106 : AOI22_X1 port map( A1 => n18041, A2 => n14304, B1 => n18042, B2 => 
                           n14212, ZN => n18016);
   U2107 : NAND2_X1 port map( A1 => n18017, A2 => n18016, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2108 : AOI22_X1 port map( A1 => n18040, A2 => n14304, B1 => n18043, B2 => 
                           n14212, ZN => n18019);
   U2109 : AOI22_X1 port map( A1 => n18041, A2 => n14306, B1 => n18042, B2 => 
                           n14210, ZN => n18018);
   U2110 : NAND2_X1 port map( A1 => n18019, A2 => n18018, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2111 : AOI22_X1 port map( A1 => n18040, A2 => n14306, B1 => n18043, B2 => 
                           n14210, ZN => n18021);
   U2112 : AOI22_X1 port map( A1 => n18041, A2 => n14308, B1 => n18042, B2 => 
                           n14208, ZN => n18020);
   U2113 : NAND2_X1 port map( A1 => n18021, A2 => n18020, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2114 : AOI22_X1 port map( A1 => n18040, A2 => n14308, B1 => n18043, B2 => 
                           n14208, ZN => n18023);
   U2115 : AOI22_X1 port map( A1 => n18041, A2 => n14310, B1 => n18042, B2 => 
                           n14206, ZN => n18022);
   U2116 : NAND2_X1 port map( A1 => n18023, A2 => n18022, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2117 : AOI22_X1 port map( A1 => n18040, A2 => n14310, B1 => n18043, B2 => 
                           n14206, ZN => n18025);
   U2118 : AOI22_X1 port map( A1 => n18041, A2 => n14312, B1 => n18042, B2 => 
                           n14204, ZN => n18024);
   U2119 : NAND2_X1 port map( A1 => n18025, A2 => n18024, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2120 : AOI22_X1 port map( A1 => n18040, A2 => n14312, B1 => n18043, B2 => 
                           n14204, ZN => n18027);
   U2121 : AOI22_X1 port map( A1 => n18041, A2 => n14314, B1 => n18042, B2 => 
                           n14202, ZN => n18026);
   U2122 : NAND2_X1 port map( A1 => n18027, A2 => n18026, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2123 : AOI22_X1 port map( A1 => n18040, A2 => n14314, B1 => n18043, B2 => 
                           n14202, ZN => n18029);
   U2124 : AOI22_X1 port map( A1 => n18041, A2 => n14316, B1 => n18042, B2 => 
                           n14200, ZN => n18028);
   U2125 : NAND2_X1 port map( A1 => n18029, A2 => n18028, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2126 : AOI22_X1 port map( A1 => n18040, A2 => n14316, B1 => n18043, B2 => 
                           n14200, ZN => n18031);
   U2127 : AOI22_X1 port map( A1 => n18041, A2 => n14318, B1 => n18042, B2 => 
                           n14198, ZN => n18030);
   U2128 : NAND2_X1 port map( A1 => n18031, A2 => n18030, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2129 : AOI22_X1 port map( A1 => n18040, A2 => n14318, B1 => n18043, B2 => 
                           n14198, ZN => n18033);
   U2130 : AOI22_X1 port map( A1 => n18041, A2 => n14320, B1 => n18042, B2 => 
                           n14196, ZN => n18032);
   U2131 : NAND2_X1 port map( A1 => n18033, A2 => n18032, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2132 : AOI22_X1 port map( A1 => n18040, A2 => n14320, B1 => n18043, B2 => 
                           n14196, ZN => n18035);
   U2133 : AOI22_X1 port map( A1 => n18041, A2 => n14322, B1 => n18042, B2 => 
                           n14194, ZN => n18034);
   U2134 : NAND2_X1 port map( A1 => n18035, A2 => n18034, ZN => n8914);
   U2135 : AOI22_X1 port map( A1 => n18040, A2 => n14322, B1 => n18043, B2 => 
                           n14194, ZN => n18037);
   U2136 : AOI22_X1 port map( A1 => n18041, A2 => n14324, B1 => n18042, B2 => 
                           n14192, ZN => n18036);
   U2137 : NAND2_X1 port map( A1 => n18037, A2 => n18036, ZN => n8913);
   U2138 : AOI22_X1 port map( A1 => n18040, A2 => n14324, B1 => n18043, B2 => 
                           n14192, ZN => n18039);
   U2139 : AOI22_X1 port map( A1 => n18041, A2 => n16414, B1 => n18042, B2 => 
                           n14190, ZN => n18038);
   U2140 : NAND2_X1 port map( A1 => n18039, A2 => n18038, ZN => n8912);
   U2141 : OAI21_X1 port map( B1 => n18041, B2 => n18040, A => n16414, ZN => 
                           n18045);
   U2142 : AOI22_X1 port map( A1 => n18043, A2 => n14190, B1 => n18042, B2 => 
                           n14279, ZN => n18044);
   U2143 : NAND2_X1 port map( A1 => n18045, A2 => n18044, ZN => n8911);
   U2144 : INV_X1 port map( A => n18046, ZN => n18054);
   U2145 : OAI222_X1 port map( A1 => n1844, A2 => n18047, B1 => n1842, B2 => 
                           n18048, C1 => n18054, C2 => n1843, ZN => n8528);
   U2146 : OAI222_X1 port map( A1 => n1840, A2 => n18047, B1 => n1838, B2 => 
                           n18048, C1 => n1839, C2 => n18054, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2147 : OAI222_X1 port map( A1 => n1837, A2 => n18054, B1 => n1836, B2 => 
                           n18048, C1 => n1838, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2148 : OAI222_X1 port map( A1 => n1834, A2 => n18054, B1 => n1833, B2 => 
                           n18048, C1 => n1836, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2149 : OAI222_X1 port map( A1 => n1832, A2 => n18054, B1 => n1831, B2 => 
                           n18048, C1 => n1833, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2150 : OAI222_X1 port map( A1 => n1830, A2 => n18054, B1 => n1829, B2 => 
                           n18048, C1 => n1831, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2151 : OAI222_X1 port map( A1 => n1828, A2 => n18054, B1 => n1827, B2 => 
                           n18048, C1 => n1829, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2152 : OAI222_X1 port map( A1 => n1826, A2 => n18054, B1 => n1825, B2 => 
                           n18048, C1 => n1827, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2153 : OAI222_X1 port map( A1 => n1824, A2 => n18054, B1 => n1823, B2 => 
                           n18048, C1 => n1825, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2154 : OAI222_X1 port map( A1 => n1822, A2 => n18054, B1 => n1821, B2 => 
                           n18048, C1 => n1823, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2155 : OAI222_X1 port map( A1 => n1820, A2 => n18054, B1 => n1819, B2 => 
                           n18048, C1 => n1821, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2156 : OAI222_X1 port map( A1 => n1818, A2 => n18054, B1 => n1817, B2 => 
                           n18048, C1 => n1819, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2157 : OAI222_X1 port map( A1 => n1816, A2 => n18054, B1 => n1815, B2 => 
                           n18048, C1 => n1817, C2 => n18047, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2158 : AOI22_X1 port map( A1 => n18052, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n18050, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n18049);
   U2159 : OAI21_X1 port map( B1 => n18054, B2 => n1814, A => n18049, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2160 : AOI22_X1 port map( A1 => n18052, A2 => n18051, B1 => n18050, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n18053);
   U2161 : OAI21_X1 port map( B1 => n18054, B2 => n1814, A => n18053, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U2162 : AOI21_X1 port map( B1 => n18057, B2 => n18056, A => n18055, ZN => 
                           n8800);
   U2163 : NOR2_X1 port map( A1 => n18058, A2 => n18079, ZN => n18064);
   U2164 : NOR2_X1 port map( A1 => n13096, A2 => n18064, ZN => n1900);
   U2165 : AOI22_X1 port map( A1 => DATA2(4), A2 => n18060, B1 => n18079, B2 =>
                           n18059, ZN => n18061);
   U2166 : INV_X1 port map( A => n13099, ZN => n18067);
   U2167 : NAND3_X1 port map( A1 => n1900, A2 => n18061, A3 => n18067, ZN => 
                           n16400);
   U2168 : NAND4_X1 port map( A1 => DATA2(1), A2 => n18064, A3 => n18082, A4 =>
                           n18062, ZN => n16401);
   U2169 : INV_X1 port map( A => n18077, ZN => n18076);
   U2170 : NAND2_X1 port map( A1 => n18076, A2 => n18063, ZN => n16403);
   U2171 : NOR4_X1 port map( A1 => DATA2(2), A2 => DATA2(3), A3 => n13099, A4 
                           => n18069, ZN => n16404);
   U2172 : NAND2_X1 port map( A1 => n18064, A2 => n18082, ZN => n18065);
   U2173 : NOR2_X1 port map( A1 => n18069, A2 => n18065, ZN => n16405);
   U2174 : NOR2_X1 port map( A1 => n18078, A2 => n18065, ZN => n16406);
   U2175 : INV_X1 port map( A => n18068, ZN => n18070);
   U2176 : NOR2_X1 port map( A1 => n18066, A2 => n18070, ZN => n16407);
   U2177 : NOR2_X1 port map( A1 => n18067, A2 => n9011, ZN => n16408);
   U2178 : NAND2_X1 port map( A1 => DATA2(1), A2 => n18068, ZN => n16409);
   U2179 : NOR2_X1 port map( A1 => n18070, A2 => n18069, ZN => n16413);
   U2180 : NOR2_X1 port map( A1 => n4302, A2 => n18071, ZN => n16415);
   U2181 : NAND2_X1 port map( A1 => n4302, A2 => n18072, ZN => n16416);
   U2182 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           A3 => n18073, ZN => n16418);
   U2183 : NOR2_X1 port map( A1 => n18075, A2 => n18074, ZN => n16419);
   U2184 : OAI21_X1 port map( B1 => DATA2(2), B2 => DATA2(1), A => n18076, ZN 
                           => n1903);
   U2185 : AOI21_X1 port map( B1 => n18079, B2 => n18078, A => n18077, ZN => 
                           n1902);
   U2186 : INV_X1 port map( A => n13096, ZN => n18080);
   U2187 : AOI21_X1 port map( B1 => n18081, B2 => n18080, A => n1900, ZN => 
                           n1901);
   U2188 : AOI21_X1 port map( B1 => n18083, B2 => n18082, A => n13099, ZN => 
                           n1893);
   U2189 : OAI22_X1 port map( A1 => n18137, A2 => n18140, B1 => n18084, B2 => 
                           n18138, ZN => n18088);
   U2190 : OAI22_X1 port map( A1 => n18086, A2 => n18150, B1 => n18085, B2 => 
                           n18152, ZN => n18087);
   U2191 : AOI211_X1 port map( C1 => n18123, C2 => n18089, A => n18088, B => 
                           n18087, ZN => n1886);
   U2192 : AOI22_X1 port map( A1 => n18144, A2 => n18091, B1 => n18123, B2 => 
                           n18090, ZN => n18094);
   U2193 : AOI22_X1 port map( A1 => n18116, A2 => n18092, B1 => n18159, B2 => 
                           n18106, ZN => n18093);
   U2194 : OAI211_X1 port map( C1 => n18100, C2 => n18148, A => n18094, B => 
                           n18093, ZN => n1885);
   U2195 : OAI22_X1 port map( A1 => n18155, A2 => n18095, B1 => n18099, B2 => 
                           n18138, ZN => n18098);
   U2196 : OAI22_X1 port map( A1 => n18137, A2 => n18096, B1 => n18100, B2 => 
                           n18152, ZN => n18097);
   U2197 : AOI211_X1 port map( C1 => n18114, C2 => n18106, A => n18098, B => 
                           n18097, ZN => n1884);
   U2198 : OAI22_X1 port map( A1 => n18155, A2 => n18100, B1 => n18099, B2 => 
                           n18150, ZN => n18105);
   U2199 : AOI22_X1 port map( A1 => n18159, A2 => n18102, B1 => n18101, B2 => 
                           n18118, ZN => n18103);
   U2200 : INV_X1 port map( A => n18103, ZN => n18104);
   U2201 : AOI211_X1 port map( C1 => n18144, C2 => n18106, A => n18105, B => 
                           n18104, ZN => n1881);
   U2202 : INV_X1 port map( A => n18115, ZN => n18121);
   U2203 : OAI22_X1 port map( A1 => n18155, A2 => n18121, B1 => n18110, B2 => 
                           n18150, ZN => n18109);
   U2204 : OAI22_X1 port map( A1 => n18137, A2 => n18107, B1 => n18111, B2 => 
                           n18138, ZN => n18108);
   U2205 : AOI211_X1 port map( C1 => n18144, C2 => n18125, A => n18109, B => 
                           n18108, ZN => n1876);
   U2206 : OAI22_X1 port map( A1 => n18110, A2 => n18148, B1 => n18121, B2 => 
                           n18152, ZN => n18113);
   U2207 : OAI22_X1 port map( A1 => n18137, A2 => n18111, B1 => n18155, B2 => 
                           n18122, ZN => n18112);
   U2208 : AOI211_X1 port map( C1 => n18114, C2 => n18125, A => n18113, B => 
                           n18112, ZN => n1874);
   U2209 : AOI22_X1 port map( A1 => n18116, A2 => n18115, B1 => n18129, B2 => 
                           n18123, ZN => n18120);
   U2210 : AOI22_X1 port map( A1 => n18118, A2 => n18125, B1 => n18159, B2 => 
                           n18117, ZN => n18119);
   U2211 : OAI211_X1 port map( C1 => n18122, C2 => n18152, A => n18120, B => 
                           n18119, ZN => n1872);
   U2212 : OAI22_X1 port map( A1 => n18122, A2 => n18150, B1 => n18121, B2 => 
                           n18138, ZN => n18128);
   U2213 : AOI22_X1 port map( A1 => n18159, A2 => n18125, B1 => n18124, B2 => 
                           n18123, ZN => n18126);
   U2214 : INV_X1 port map( A => n18126, ZN => n18127);
   U2215 : AOI211_X1 port map( C1 => n18144, C2 => n18129, A => n18128, B => 
                           n18127, ZN => n1871);
   U2216 : OAI22_X1 port map( A1 => n14133, A2 => n18131, B1 => n14382, B2 => 
                           n18130, ZN => n18132);
   U2217 : NAND2_X1 port map( A1 => n14368, A2 => n18132, ZN => n18134);
   U2218 : AOI211_X1 port map( C1 => n13878, C2 => n14008, A => n14007, B => 
                           n13975, ZN => n18133);
   U2219 : NAND3_X1 port map( A1 => n18134, A2 => n18133, A3 => n14272, ZN => 
                           OUTALU(6));
   U2220 : INV_X1 port map( A => n8647, ZN => n18145);
   U2221 : AOI22_X1 port map( A1 => n1894, A2 => n18145, B1 => n11927, B2 => 
                           n1865, ZN => n1864);
   U2222 : OAI22_X1 port map( A1 => n18137, A2 => n18136, B1 => n18135, B2 => 
                           n18150, ZN => n18142);
   U2223 : OAI22_X1 port map( A1 => n18155, A2 => n18140, B1 => n18139, B2 => 
                           n18138, ZN => n18141);
   U2224 : AOI211_X1 port map( C1 => n18144, C2 => n18143, A => n18142, B => 
                           n18141, ZN => n1863);
   U2225 : AOI22_X1 port map( A1 => n1898, A2 => n1859, B1 => n13151, B2 => 
                           n18145, ZN => n1860);
   U2226 : INV_X1 port map( A => n8604, ZN => n18146);
   U2227 : AOI22_X1 port map( A1 => n11927, A2 => n1857, B1 => n1894, B2 => 
                           n18146, ZN => n1858);
   U2228 : INV_X1 port map( A => n18147, ZN => n18149);
   U2229 : OAI22_X1 port map( A1 => n18151, A2 => n18150, B1 => n18149, B2 => 
                           n18148, ZN => n18157);
   U2230 : OAI22_X1 port map( A1 => n18155, A2 => n18154, B1 => n18153, B2 => 
                           n18152, ZN => n18156);
   U2231 : AOI211_X1 port map( C1 => n18159, C2 => n18158, A => n18157, B => 
                           n18156, ZN => n1856);
   U2232 : NOR3_X1 port map( A1 => n18162, A2 => n18161, A3 => n18160, ZN => 
                           n18169);
   U2233 : AOI221_X1 port map( B1 => n18167, B2 => n18166, C1 => n18165, C2 => 
                           n18164, A => n18163, ZN => n18168);
   U2234 : AOI211_X1 port map( C1 => n18171, C2 => n18170, A => n18169, B => 
                           n18168, ZN => n1811);
   U2235 : AOI22_X1 port map( A1 => n18175, A2 => n18174, B1 => n18173, B2 => 
                           n18172, ZN => n1810);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n18281, n18282, n18283, n18284, n18293, n18294, n18295, n18296, 
      n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, 
      n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, 
      n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, 
      n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, 
      n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, 
      n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, 
      n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, 
      n18360, n19395, n19396, n19397, n19398, n19399, n19400, n19402, n29018, 
      n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, 
      n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, 
      n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, 
      n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, 
      n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, 
      n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, 
      n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, 
      n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, 
      n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, 
      n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, 
      n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, 
      n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, 
      n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, 
      n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, 
      n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, 
      n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, 
      n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, 
      n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, 
      n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, 
      n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, 
      n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, 
      n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, 
      n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, 
      n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, 
      n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, 
      n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, 
      n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, 
      n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, 
      n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, 
      n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, 
      n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, 
      n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, 
      n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, 
      n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, 
      n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, 
      n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, 
      n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, 
      n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, 
      n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, 
      n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, 
      n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, 
      n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, 
      n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, 
      n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, 
      n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, 
      n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, 
      n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, 
      n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, 
      n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, 
      n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, 
      n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, 
      n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, 
      n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, 
      n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, 
      n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, 
      n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, 
      n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, 
      n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, 
      n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, 
      n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, 
      n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, 
      n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, 
      n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, 
      n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, 
      n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, 
      n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, 
      n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, 
      n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, 
      n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, 
      n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, 
      n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, 
      n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, 
      n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, 
      n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, 
      n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, 
      n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, 
      n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, 
      n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, 
      n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, 
      n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, 
      n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, 
      n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, 
      n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, 
      n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, 
      n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, 
      n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, 
      n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, 
      n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, 
      n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, 
      n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, 
      n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, 
      n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, 
      n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, 
      n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, 
      n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, 
      n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, 
      n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, 
      n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, 
      n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, 
      n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, 
      n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, 
      n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, 
      n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, 
      n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, 
      n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, 
      n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, 
      n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, 
      n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, 
      n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, 
      n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, 
      n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, 
      n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, 
      n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, 
      n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, 
      n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, 
      n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, 
      n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, 
      n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, 
      n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, 
      n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, 
      n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, 
      n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, 
      n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, 
      n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, 
      n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, 
      n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, 
      n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, 
      n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, 
      n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, 
      n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, 
      n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, 
      n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, 
      n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, 
      n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, 
      n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, 
      n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, 
      n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, 
      n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, 
      n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, 
      n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, 
      n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, 
      n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, 
      n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, 
      n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, 
      n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, 
      n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, 
      n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, 
      n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, 
      n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, 
      n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, 
      n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, 
      n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, 
      n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, 
      n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, 
      n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, 
      n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, 
      n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, 
      n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, 
      n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, 
      n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, 
      n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, 
      n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, 
      n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, 
      n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, 
      n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, 
      n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, 
      n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, 
      n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, 
      n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, 
      n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, 
      n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, 
      n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, 
      n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, 
      n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, 
      n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, 
      n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, 
      n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, 
      n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, 
      n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, 
      n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, 
      n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, 
      n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, 
      n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, 
      n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, 
      n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, 
      n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, 
      n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, 
      n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, 
      n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, 
      n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, 
      n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, 
      n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, 
      n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, 
      n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, 
      n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, 
      n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, 
      n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, 
      n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, 
      n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, 
      n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, 
      n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, 
      n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, 
      n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, 
      n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, 
      n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, 
      n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, 
      n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, 
      n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, 
      n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, 
      n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, 
      n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, 
      n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, 
      n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, 
      n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, 
      n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, 
      n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, 
      n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, 
      n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, 
      n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, 
      n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, 
      n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, 
      n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, 
      n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, 
      n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, 
      n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, 
      n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, 
      n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, 
      n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, 
      n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, 
      n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, 
      n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, 
      n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, 
      n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, 
      n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, 
      n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, 
      n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, 
      n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, 
      n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, 
      n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, 
      n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, 
      n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, 
      n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, 
      n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, 
      n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, 
      n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, 
      n31224, n31225, n31226, n31227, n31228, n31229, n31231, n31233, n31234, 
      n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, 
      n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, 
      n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, 
      n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, 
      n31271, n31273, n35759, n35760, n2534, n2535, n2536, n2537, n2538, n2539,
      n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
      n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, 
      n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
      n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
      n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
      n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
      n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
      n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
      n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
      n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
      n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
      n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
      n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
      n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
      n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, 
      n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
      n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
      n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
      n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
      n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
      n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
      n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
      n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
      n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
      n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
      n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
      n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, 
      n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, 
      n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
      n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
      n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
      n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
      n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
      n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
      n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
      n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
      n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
      n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
      n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
      n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
      n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
      n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
      n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
      n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
      n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
      n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
      n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
      n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
      n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
      n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
      n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
      n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
      n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
      n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
      n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, 
      n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
      n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
      n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
      n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
      n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
      n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
      n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
      n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, 
      n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
      n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
      n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
      n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, 
      n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, 
      n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
      n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
      n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
      n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, 
      n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
      n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, 
      n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, 
      n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, 
      n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, 
      n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, 
      n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, 
      n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, 
      n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, 
      n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n35761, n35762, 
      n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, 
      n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, 
      n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, 
      n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, 
      n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, 
      n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, 
      n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, 
      n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, 
      n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, 
      n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, 
      n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, 
      n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, 
      n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, 
      n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, 
      n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, 
      n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, 
      n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, 
      n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, 
      n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, 
      n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, 
      n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, 
      n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, 
      n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, 
      n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, 
      n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, 
      n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, 
      n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, 
      n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, 
      n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, 
      n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, 
      n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, 
      n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, 
      n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, 
      n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, 
      n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, 
      n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, 
      n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, 
      n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, 
      n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, 
      n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, 
      n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, 
      n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, 
      n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, 
      n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, 
      n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, 
      n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, 
      n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, 
      n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, 
      n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, 
      n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, 
      n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, 
      n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, 
      n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, 
      n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, 
      n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, 
      n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, 
      n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, 
      n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, 
      n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, 
      n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, 
      n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, 
      n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, 
      n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, 
      n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, 
      n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, 
      n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, 
      n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, 
      n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, 
      n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, 
      n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, 
      n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, 
      n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, 
      n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, 
      n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, 
      n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, 
      n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, 
      n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, 
      n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, 
      n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, 
      n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, 
      n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, 
      n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, 
      n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, 
      n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, 
      n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, 
      n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, 
      n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, 
      n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, 
      n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, 
      n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, 
      n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, 
      n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, 
      n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, 
      n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, 
      n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, 
      n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, 
      n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, 
      n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, 
      n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, 
      n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, 
      n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, 
      n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, 
      n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, 
      n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, 
      n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, 
      n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, 
      n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, 
      n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, 
      n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, 
      n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, 
      n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, 
      n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, 
      n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, 
      n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, 
      n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, 
      n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, 
      n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, 
      n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, 
      n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, 
      n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, 
      n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, 
      n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, 
      n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, 
      n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, 
      n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, 
      n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896, 
      n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905, 
      n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, 
      n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923, 
      n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932, 
      n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941, 
      n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950, 
      n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959, 
      n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968, 
      n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977, 
      n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986, 
      n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995, 
      n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004, 
      n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013, 
      n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022, 
      n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031, 
      n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040, 
      n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049, 
      n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058, 
      n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067, 
      n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076, 
      n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085, 
      n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094, 
      n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103, 
      n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112, 
      n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121, 
      n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, 
      n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, 
      n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, 
      n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, 
      n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, 
      n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, 
      n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, 
      n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, 
      n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, 
      n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, 
      n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, 
      n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, 
      n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, 
      n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, 
      n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, 
      n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, 
      n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, 
      n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, 
      n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, 
      n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, 
      n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, 
      n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, 
      n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, 
      n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, 
      n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, 
      n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, 
      n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, 
      n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, 
      n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, 
      n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, 
      n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, 
      n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, 
      n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, 
      n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, 
      n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, 
      n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, 
      n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, 
      n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, 
      n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, 
      n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, 
      n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, 
      n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, 
      n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, 
      n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, 
      n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, 
      n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, 
      n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, 
      n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, 
      n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, 
      n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, 
      n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, 
      n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, 
      n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, 
      n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, 
      n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, 
      n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, 
      n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, 
      n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, 
      n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, 
      n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, 
      n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, 
      n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, 
      n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, 
      n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, 
      n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, 
      n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, 
      n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, 
      n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, 
      n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, 
      n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, 
      n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, 
      n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, 
      n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, 
      n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, 
      n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, 
      n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, 
      n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, 
      n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, 
      n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, 
      n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, 
      n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, 
      n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, 
      n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, 
      n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, 
      n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, 
      n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, 
      n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, 
      n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, 
      n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922, 
      n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, 
      n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940, 
      n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949, 
      n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958, 
      n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967, 
      n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976, 
      n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985, 
      n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994, 
      n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003, 
      n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012, 
      n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, 
      n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, 
      n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, 
      n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, 
      n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, 
      n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066, 
      n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075, 
      n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084, 
      n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093, 
      n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102, 
      n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111, 
      n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120, 
      n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129, 
      n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138, 
      n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147, 
      n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156, 
      n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165, 
      n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174, 
      n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183, 
      n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192, 
      n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, 
      n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, 
      n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, 
      n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, 
      n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, 
      n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, 
      n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, 
      n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, 
      n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, 
      n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282, 
      n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291, 
      n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300, 
      n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309, 
      n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318, 
      n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327, 
      n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336, 
      n38337, n38338, n38339, n38340, n38341, n38342, n_1576, n_1577, n_1578, 
      n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, 
      n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, 
      n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, 
      n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, 
      n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, 
      n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, 
      n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, 
      n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, 
      n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, 
      n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, 
      n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, 
      n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, 
      n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, 
      n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, 
      n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, 
      n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, 
      n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, 
      n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, 
      n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, 
      n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, 
      n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, 
      n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, 
      n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, 
      n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, 
      n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, 
      n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, 
      n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, 
      n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, 
      n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, 
      n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, 
      n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, 
      n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, 
      n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, 
      n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, 
      n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, 
      n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, 
      n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, 
      n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, 
      n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, 
      n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, 
      n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, 
      n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, 
      n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, 
      n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, 
      n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, 
      n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, 
      n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, 
      n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, 
      n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, 
      n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, 
      n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, 
      n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, 
      n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, 
      n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, 
      n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, 
      n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, 
      n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, 
      n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, 
      n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, 
      n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, 
      n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, 
      n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, 
      n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, 
      n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, 
      n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, 
      n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, 
      n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, 
      n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, 
      n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, 
      n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, 
      n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, 
      n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, 
      n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, 
      n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, 
      n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, 
      n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, 
      n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, 
      n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, 
      n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, 
      n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, 
      n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, 
      n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, 
      n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, 
      n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, 
      n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, 
      n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, 
      n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, 
      n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, 
      n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, 
      n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, 
      n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, 
      n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, 
      n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, 
      n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, 
      n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, 
      n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, 
      n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, 
      n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, 
      n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, 
      n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, 
      n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, 
      n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, 
      n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, 
      n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, 
      n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, 
      n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, 
      n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, 
      n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, 
      n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, 
      n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, 
      n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, 
      n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, 
      n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, 
      n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, 
      n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, 
      n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, 
      n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, 
      n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, 
      n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, 
      n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, 
      n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, 
      n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, 
      n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, 
      n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, 
      n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, 
      n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, 
      n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, 
      n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, 
      n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, 
      n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, 
      n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, 
      n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, 
      n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, 
      n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, 
      n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, 
      n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, 
      n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, 
      n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, 
      n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, 
      n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, 
      n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, 
      n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, 
      n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, 
      n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, 
      n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, 
      n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, 
      n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, 
      n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, 
      n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, 
      n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, 
      n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, 
      n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, 
      n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, 
      n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, 
      n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, 
      n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, 
      n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, 
      n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, 
      n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, 
      n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, 
      n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, 
      n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, 
      n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, 
      n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, 
      n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, 
      n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, 
      n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, 
      n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, 
      n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, 
      n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, 
      n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, 
      n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, 
      n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, 
      n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, 
      n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, 
      n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, 
      n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, 
      n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, 
      n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, 
      n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, 
      n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, 
      n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, 
      n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, 
      n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, 
      n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, 
      n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, 
      n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, 
      n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, 
      n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, 
      n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, 
      n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, 
      n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, 
      n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, 
      n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, 
      n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, 
      n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, 
      n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, 
      n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, 
      n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, 
      n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, 
      n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, 
      n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, 
      n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, 
      n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, 
      n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, 
      n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, 
      n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, 
      n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, 
      n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, 
      n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, 
      n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, 
      n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, 
      n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, 
      n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, 
      n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, 
      n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, 
      n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, 
      n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, 
      n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, 
      n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, 
      n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, 
      n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, 
      n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, 
      n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, 
      n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, 
      n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, 
      n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, 
      n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, 
      n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, 
      n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, 
      n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, 
      n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, 
      n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, 
      n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, 
      n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, 
      n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, 
      n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, 
      n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, 
      n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, 
      n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, 
      n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, 
      n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, 
      n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, 
      n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, 
      n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, 
      n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, 
      n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, 
      n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, 
      n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, 
      n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, 
      n_3829, n_3830 : std_logic;

begin
   
   clk_r_REG9980_S1 : DFFR_X1 port map( D => ENABLE, CK => CLK, RN => RESET_BAR
                           , Q => n31273, QN => n_1576);
   clk_r_REG10013_S1 : DFFR_X1 port map( D => RD1, CK => CLK, RN => RESET_BAR, 
                           Q => n31271, QN => n_1577);
   clk_r_REG10116_S2 : DFFR_X1 port map( D => RD2, CK => CLK, RN => RESET_BAR, 
                           Q => n31270, QN => n_1578);
   clk_r_REG10287_S7 : DFFR_X1 port map( D => ADD_RD1(4), CK => CLK, RN => 
                           RESET_BAR, Q => n31269, QN => n_1579);
   clk_r_REG10289_S7 : DFFS_X1 port map( D => n3560, CK => CLK, SN => RESET_BAR
                           , Q => n_1580, QN => n31268);
   clk_r_REG10244_S7 : DFFR_X1 port map( D => ADD_RD2(4), CK => CLK, RN => 
                           RESET_BAR, Q => n31267, QN => n_1581);
   clk_r_REG10247_S7 : DFFS_X1 port map( D => n3569, CK => CLK, SN => RESET_BAR
                           , Q => n_1582, QN => n31266);
   clk_r_REG7003_S6 : DFFR_X1 port map( D => DATAIN(31), CK => CLK, RN => 
                           RESET_BAR, Q => n31265, QN => n_1583);
   clk_r_REG6994_S6 : DFFR_X1 port map( D => DATAIN(30), CK => CLK, RN => 
                           RESET_BAR, Q => n31264, QN => n_1584);
   clk_r_REG6985_S5 : DFFR_X1 port map( D => DATAIN(29), CK => CLK, RN => 
                           RESET_BAR, Q => n31263, QN => n_1585);
   clk_r_REG6978_S6 : DFFR_X1 port map( D => DATAIN(28), CK => CLK, RN => 
                           RESET_BAR, Q => n31262, QN => n_1586);
   clk_r_REG6971_S5 : DFFR_X1 port map( D => DATAIN(27), CK => CLK, RN => 
                           RESET_BAR, Q => n31261, QN => n_1587);
   clk_r_REG6964_S6 : DFFR_X1 port map( D => DATAIN(26), CK => CLK, RN => 
                           RESET_BAR, Q => n31260, QN => n_1588);
   clk_r_REG6956_S5 : DFFR_X1 port map( D => DATAIN(25), CK => CLK, RN => 
                           RESET_BAR, Q => n31259, QN => n_1589);
   clk_r_REG7104_S12 : DFFR_X1 port map( D => DATAIN(24), CK => CLK, RN => 
                           RESET_BAR, Q => n31258, QN => n_1590);
   clk_r_REG7025_S5 : DFFR_X1 port map( D => DATAIN(23), CK => CLK, RN => 
                           RESET_BAR, Q => n31257, QN => n_1591);
   clk_r_REG7017_S5 : DFFR_X1 port map( D => DATAIN(22), CK => CLK, RN => 
                           RESET_BAR, Q => n31256, QN => n_1592);
   clk_r_REG7144_S5 : DFFR_X1 port map( D => DATAIN(21), CK => CLK, RN => 
                           RESET_BAR, Q => n31255, QN => n_1593);
   clk_r_REG6949_S11 : DFFR_X1 port map( D => DATAIN(20), CK => CLK, RN => 
                           RESET_BAR, Q => n31254, QN => n_1594);
   clk_r_REG7137_S5 : DFFR_X1 port map( D => DATAIN(19), CK => CLK, RN => 
                           RESET_BAR, Q => n31253, QN => n_1595);
   clk_r_REG7130_S5 : DFFR_X1 port map( D => DATAIN(18), CK => CLK, RN => 
                           RESET_BAR, Q => n31252, QN => n_1596);
   clk_r_REG7123_S5 : DFFR_X1 port map( D => DATAIN(17), CK => CLK, RN => 
                           RESET_BAR, Q => n31251, QN => n_1597);
   clk_r_REG7116_S5 : DFFR_X1 port map( D => DATAIN(16), CK => CLK, RN => 
                           RESET_BAR, Q => n31250, QN => n_1598);
   clk_r_REG7235_S11 : DFFR_X1 port map( D => DATAIN(15), CK => CLK, RN => 
                           RESET_BAR, Q => n31249, QN => n_1599);
   clk_r_REG7254_S4 : DFFR_X1 port map( D => DATAIN(14), CK => CLK, RN => 
                           RESET_BAR, Q => n31248, QN => n_1600);
   clk_r_REG7184_S11 : DFFR_X1 port map( D => DATAIN(13), CK => CLK, RN => 
                           RESET_BAR, Q => n31247, QN => n_1601);
   clk_r_REG7166_S5 : DFFR_X1 port map( D => DATAIN(12), CK => CLK, RN => 
                           RESET_BAR, Q => n31246, QN => n_1602);
   clk_r_REG7063_S12 : DFFR_X1 port map( D => DATAIN(11), CK => CLK, RN => 
                           RESET_BAR, Q => n31245, QN => n_1603);
   clk_r_REG7044_S5 : DFFR_X1 port map( D => DATAIN(10), CK => CLK, RN => 
                           RESET_BAR, Q => n31244, QN => n_1604);
   clk_r_REG7327_S4 : DFFR_X1 port map( D => DATAIN(9), CK => CLK, RN => 
                           RESET_BAR, Q => n31243, QN => n_1605);
   clk_r_REG7397_S4 : DFFR_X1 port map( D => DATAIN(8), CK => CLK, RN => 
                           RESET_BAR, Q => n31242, QN => n_1606);
   clk_r_REG7546_S4 : DFFR_X1 port map( D => DATAIN(7), CK => CLK, RN => 
                           RESET_BAR, Q => n31241, QN => n_1607);
   clk_r_REG7641_S11 : DFFR_X1 port map( D => DATAIN(6), CK => CLK, RN => 
                           RESET_BAR, Q => n31240, QN => n_1608);
   clk_r_REG7532_S10 : DFFR_X1 port map( D => DATAIN(5), CK => CLK, RN => 
                           RESET_BAR, Q => n31239, QN => n_1609);
   clk_r_REG7742_S8 : DFFR_X1 port map( D => DATAIN(4), CK => CLK, RN => 
                           RESET_BAR, Q => n31238, QN => n_1610);
   clk_r_REG6934_S7 : DFFR_X1 port map( D => DATAIN(3), CK => CLK, RN => 
                           RESET_BAR, Q => n31237, QN => n_1611);
   clk_r_REG7384_S5 : DFFR_X1 port map( D => DATAIN(2), CK => CLK, RN => 
                           RESET_BAR, Q => n31236, QN => n_1612);
   clk_r_REG7308_S5 : DFFR_X1 port map( D => DATAIN(1), CK => CLK, RN => 
                           RESET_BAR, Q => n31235, QN => n_1613);
   clk_r_REG6921_S11 : DFFR_X1 port map( D => DATAIN(0), CK => CLK, RN => 
                           RESET_BAR, Q => n31234, QN => n_1614);
   clk_r_REG10240_S7 : DFFS_X1 port map( D => n3570, CK => CLK, SN => RESET_BAR
                           , Q => n31233, QN => n_1615);
   clk_r_REG10059_S3 : DFFS_X1 port map( D => n3559, CK => CLK, SN => RESET_BAR
                           , Q => n_1616, QN => n35760);
   clk_r_REG10060_S4 : DFFR_X1 port map( D => n35760, CK => CLK, RN => 
                           RESET_BAR, Q => n_1617, QN => n31231);
   clk_r_REG10055_S3 : DFFS_X1 port map( D => n3558, CK => CLK, SN => RESET_BAR
                           , Q => n_1618, QN => n35759);
   clk_r_REG10056_S4 : DFFR_X1 port map( D => n35759, CK => CLK, RN => 
                           RESET_BAR, Q => n_1619, QN => n31229);
   clk_r_REG10237_S7 : DFFR_X1 port map( D => n18314, CK => CLK, RN => 
                           RESET_BAR, Q => n31228, QN => n_1620);
   clk_r_REG10209_S7 : DFFR_X1 port map( D => n18317, CK => CLK, RN => 
                           RESET_BAR, Q => n31227, QN => n_1621);
   clk_r_REG10217_S7 : DFFR_X1 port map( D => n18320, CK => CLK, RN => 
                           RESET_BAR, Q => n31226, QN => n_1622);
   clk_r_REG10239_S7 : DFFR_X1 port map( D => n18316, CK => CLK, RN => 
                           RESET_BAR, Q => n31225, QN => n_1623);
   clk_r_REG10211_S7 : DFFR_X1 port map( D => n18321, CK => CLK, RN => 
                           RESET_BAR, Q => n31224, QN => n_1624);
   clk_r_REG10223_S7 : DFFR_X1 port map( D => n18310, CK => CLK, RN => 
                           RESET_BAR, Q => n31223, QN => n_1625);
   clk_r_REG10230_S7 : DFFR_X1 port map( D => n18315, CK => CLK, RN => 
                           RESET_BAR, Q => n31222, QN => n_1626);
   clk_r_REG10234_S7 : DFFR_X1 port map( D => n3573, CK => CLK, RN => RESET_BAR
                           , Q => n31221, QN => n_1627);
   clk_r_REG10228_S7 : DFFR_X1 port map( D => n3574, CK => CLK, RN => RESET_BAR
                           , Q => n31220, QN => n_1628);
   clk_r_REG10242_S7 : DFFS_X1 port map( D => n3570, CK => CLK, SN => RESET_BAR
                           , Q => n31219, QN => n_1629);
   clk_r_REG10199_S7 : DFFR_X1 port map( D => n3571, CK => CLK, RN => RESET_BAR
                           , Q => n31218, QN => n_1630);
   clk_r_REG10206_S7 : DFFR_X1 port map( D => n3576, CK => CLK, RN => RESET_BAR
                           , Q => n31217, QN => n_1631);
   clk_r_REG10214_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR
                           , Q => n31215, QN => n_1632);
   clk_r_REG10227_S7 : DFFR_X1 port map( D => n3574, CK => CLK, RN => RESET_BAR
                           , Q => n31214, QN => n_1633);
   clk_r_REG10190_S7 : DFFR_X1 port map( D => n18313, CK => CLK, RN => 
                           RESET_BAR, Q => n31213, QN => n_1634);
   clk_r_REG10188_S7 : DFFR_X1 port map( D => n18312, CK => CLK, RN => 
                           RESET_BAR, Q => n31212, QN => n_1635);
   clk_r_REG10232_S7 : DFFR_X1 port map( D => n18324, CK => CLK, RN => 
                           RESET_BAR, Q => n31211, QN => n_1636);
   clk_r_REG10200_S7 : DFFR_X1 port map( D => n3571, CK => CLK, RN => RESET_BAR
                           , Q => n31210, QN => n_1637);
   clk_r_REG10221_S7 : DFFR_X1 port map( D => n19402, CK => CLK, RN => 
                           RESET_BAR, Q => n31209, QN => n_1638);
   clk_r_REG10192_S7 : DFFR_X1 port map( D => n3577, CK => CLK, RN => RESET_BAR
                           , Q => n31208, QN => n_1639);
   clk_r_REG10219_S7 : DFFR_X1 port map( D => n18322, CK => CLK, RN => 
                           RESET_BAR, Q => n31207, QN => n_1640);
   clk_r_REG10195_S7 : DFFR_X1 port map( D => n18309, CK => CLK, RN => 
                           RESET_BAR, Q => n31206, QN => n_1641);
   clk_r_REG10225_S7 : DFFR_X1 port map( D => n18323, CK => CLK, RN => 
                           RESET_BAR, Q => n31205, QN => n_1642);
   clk_r_REG10235_S7 : DFFR_X1 port map( D => n3573, CK => CLK, RN => RESET_BAR
                           , Q => n31204, QN => n_1643);
   clk_r_REG10204_S7 : DFFR_X1 port map( D => n18319, CK => CLK, RN => 
                           RESET_BAR, Q => n31203, QN => n_1644);
   clk_r_REG10213_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR
                           , Q => n31202, QN => n_1645);
   clk_r_REG10193_S7 : DFFR_X1 port map( D => n3577, CK => CLK, RN => RESET_BAR
                           , Q => n31201, QN => n_1646);
   clk_r_REG10202_S7 : DFFR_X1 port map( D => n18311, CK => CLK, RN => 
                           RESET_BAR, Q => n31200, QN => n_1647);
   clk_r_REG10197_S7 : DFFR_X1 port map( D => n18318, CK => CLK, RN => 
                           RESET_BAR, Q => n31199, QN => n_1648);
   clk_r_REG10174_S7 : DFFR_X1 port map( D => n18299, CK => CLK, RN => 
                           RESET_BAR, Q => n31198, QN => n_1649);
   clk_r_REG10167_S7 : DFFR_X1 port map( D => n18294, CK => CLK, RN => 
                           RESET_BAR, Q => n31197, QN => n_1650);
   clk_r_REG10155_S7 : DFFR_X1 port map( D => n18302, CK => CLK, RN => 
                           RESET_BAR, Q => n31196, QN => n_1651);
   clk_r_REG10169_S7 : DFFR_X1 port map( D => n18304, CK => CLK, RN => 
                           RESET_BAR, Q => n31195, QN => n_1652);
   clk_r_REG10157_S7 : DFFR_X1 port map( D => n19397, CK => CLK, RN => 
                           RESET_BAR, Q => n31194, QN => n_1653);
   clk_r_REG10135_S7 : DFFR_X1 port map( D => n3568, CK => CLK, RN => RESET_BAR
                           , Q => n31193, QN => n_1654);
   clk_r_REG10143_S7 : DFFR_X1 port map( D => n19396, CK => CLK, RN => 
                           RESET_BAR, Q => n31192, QN => n_1655);
   clk_r_REG10184_S7 : DFFR_X1 port map( D => n3563, CK => CLK, RN => RESET_BAR
                           , Q => n31191, QN => n_1656);
   clk_r_REG10133_S7 : DFFR_X1 port map( D => n18307, CK => CLK, RN => 
                           RESET_BAR, Q => n31189, QN => n_1657);
   clk_r_REG10176_S7 : DFFR_X1 port map( D => n18303, CK => CLK, RN => 
                           RESET_BAR, Q => n31188, QN => n_1658);
   clk_r_REG10171_S7 : DFFR_X1 port map( D => n19395, CK => CLK, RN => 
                           RESET_BAR, Q => n31187, QN => n_1659);
   clk_r_REG10150_S7 : DFFS_X1 port map( D => n19400, CK => CLK, SN => 
                           RESET_BAR, Q => n31186, QN => n_1660);
   clk_r_REG10162_S7 : DFFR_X1 port map( D => n18305, CK => CLK, RN => 
                           RESET_BAR, Q => n31185, QN => n_1661);
   clk_r_REG10148_S7 : DFFR_X1 port map( D => n18308, CK => CLK, RN => 
                           RESET_BAR, Q => n31184, QN => n_1662);
   clk_r_REG10146_S7 : DFFR_X1 port map( D => n18306, CK => CLK, RN => 
                           RESET_BAR, Q => n31183, QN => n_1663);
   clk_r_REG10164_S7 : DFFR_X1 port map( D => n19399, CK => CLK, RN => 
                           RESET_BAR, Q => n31182, QN => n_1664);
   clk_r_REG10180_S7 : DFFR_X1 port map( D => n18297, CK => CLK, RN => 
                           RESET_BAR, Q => n31181, QN => n_1665);
   clk_r_REG10178_S7 : DFFR_X1 port map( D => n19398, CK => CLK, RN => 
                           RESET_BAR, Q => n31180, QN => n_1666);
   clk_r_REG10185_S7 : DFFR_X1 port map( D => n3563, CK => CLK, RN => RESET_BAR
                           , Q => n31179, QN => n_1667);
   clk_r_REG10160_S7 : DFFR_X1 port map( D => n18301, CK => CLK, RN => 
                           RESET_BAR, Q => n31178, QN => n_1668);
   clk_r_REG10182_S7 : DFFR_X1 port map( D => n18298, CK => CLK, RN => 
                           RESET_BAR, Q => n31177, QN => n_1669);
   clk_r_REG10131_S7 : DFFR_X1 port map( D => n18300, CK => CLK, RN => 
                           RESET_BAR, Q => n31176, QN => n_1670);
   clk_r_REG10139_S7 : DFFR_X1 port map( D => n18293, CK => CLK, RN => 
                           RESET_BAR, Q => n31175, QN => n_1671);
   clk_r_REG10153_S7 : DFFR_X1 port map( D => n18295, CK => CLK, RN => 
                           RESET_BAR, Q => n31174, QN => n_1672);
   clk_r_REG10141_S7 : DFFR_X1 port map( D => n18296, CK => CLK, RN => 
                           RESET_BAR, Q => n31173, QN => n_1673);
   clk_r_REG8974_S1 : DFF_X1 port map( D => n3024, CK => CLK, Q => n31172, QN 
                           => n_1674);
   clk_r_REG10156_S7 : DFFR_X1 port map( D => n19397, CK => CLK, RN => 
                           RESET_BAR, Q => n31171, QN => n_1675);
   clk_r_REG10163_S7 : DFFR_X1 port map( D => n19399, CK => CLK, RN => 
                           RESET_BAR, Q => n31170, QN => n_1676);
   clk_r_REG10177_S7 : DFFR_X1 port map( D => n19398, CK => CLK, RN => 
                           RESET_BAR, Q => n31169, QN => n_1677);
   clk_r_REG10220_S7 : DFFR_X1 port map( D => n19402, CK => CLK, RN => 
                           RESET_BAR, Q => n31168, QN => n_1678);
   clk_r_REG10142_S7 : DFFR_X1 port map( D => n19396, CK => CLK, RN => 
                           RESET_BAR, Q => n31167, QN => n_1679);
   clk_r_REG10149_S7 : DFFS_X1 port map( D => n19400, CK => CLK, SN => 
                           RESET_BAR, Q => n31166, QN => n_1680);
   clk_r_REG10241_S7 : DFFS_X1 port map( D => n3570, CK => CLK, SN => RESET_BAR
                           , Q => n31165, QN => n_1681);
   clk_r_REG10170_S7 : DFFR_X1 port map( D => n19395, CK => CLK, RN => 
                           RESET_BAR, Q => n31164, QN => n_1682);
   clk_r_REG9038_S1 : DFF_X1 port map( D => n2767, CK => CLK, Q => n31163, QN 
                           => n_1683);
   clk_r_REG10233_S7 : DFFR_X1 port map( D => n3573, CK => CLK, RN => RESET_BAR
                           , Q => n31162, QN => n_1684);
   clk_r_REG10226_S7 : DFFR_X1 port map( D => n3574, CK => CLK, RN => RESET_BAR
                           , Q => n31161, QN => n_1685);
   clk_r_REG10183_S7 : DFFR_X1 port map( D => n3563, CK => CLK, RN => RESET_BAR
                           , Q => n31160, QN => n_1686);
   clk_r_REG10134_S7 : DFFR_X1 port map( D => n3568, CK => CLK, RN => RESET_BAR
                           , Q => n31159, QN => n_1687);
   clk_r_REG10191_S7 : DFFR_X1 port map( D => n3577, CK => CLK, RN => RESET_BAR
                           , Q => n31158, QN => n_1688);
   clk_r_REG10198_S7 : DFFR_X1 port map( D => n3571, CK => CLK, RN => RESET_BAR
                           , Q => n31157, QN => n_1689);
   clk_r_REG10212_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR
                           , Q => n31156, QN => n_1690);
   clk_r_REG10205_S7 : DFFR_X1 port map( D => n3576, CK => CLK, RN => RESET_BAR
                           , Q => n31155, QN => n_1691);
   clk_r_REG7614_S1 : DFF_X1 port map( D => n3309, CK => CLK, Q => n31154, QN 
                           => n_1692);
   clk_r_REG7616_S1 : DFF_X1 port map( D => n3308, CK => CLK, Q => n31153, QN 
                           => n_1693);
   clk_r_REG7618_S1 : DFF_X1 port map( D => n3307, CK => CLK, Q => n31152, QN 
                           => n_1694);
   clk_r_REG7620_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n31151, QN 
                           => n_1695);
   clk_r_REG7704_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n31150, QN 
                           => n_1696);
   clk_r_REG7622_S1 : DFF_X1 port map( D => n3305, CK => CLK, Q => n31149, QN 
                           => n_1697);
   clk_r_REG7624_S1 : DFF_X1 port map( D => n3304, CK => CLK, Q => n31148, QN 
                           => n_1698);
   clk_r_REG7918_S1 : DFF_X1 port map( D => n3406, CK => CLK, Q => n31147, QN 
                           => n_1699);
   clk_r_REG7706_S1 : DFF_X1 port map( D => n3341, CK => CLK, Q => n31146, QN 
                           => n_1700);
   clk_r_REG9874_S1 : DFF_X1 port map( D => n3438, CK => CLK, Q => n31145, QN 
                           => n_1701);
   clk_r_REG7626_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n31144, QN 
                           => n_1702);
   clk_r_REG7708_S1 : DFF_X1 port map( D => n3340, CK => CLK, Q => n31143, QN 
                           => n_1703);
   clk_r_REG8259_S1 : DFF_X1 port map( D => n3470, CK => CLK, Q => n31142, QN 
                           => n_1704);
   clk_r_REG8261_S1 : DFF_X1 port map( D => n3469, CK => CLK, Q => n31141, QN 
                           => n_1705);
   clk_r_REG8399_S1 : DFF_X1 port map( D => n3502, CK => CLK, Q => n31140, QN 
                           => n_1706);
   clk_r_REG7628_S1 : DFF_X1 port map( D => n3302, CK => CLK, Q => n31139, QN 
                           => n_1707);
   clk_r_REG8263_S1 : DFF_X1 port map( D => n3468, CK => CLK, Q => n31138, QN 
                           => n_1708);
   clk_r_REG7548_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n31137, QN 
                           => n_1709);
   clk_r_REG8265_S1 : DFF_X1 port map( D => n3467, CK => CLK, Q => n31136, QN 
                           => n_1710);
   clk_r_REG8267_S1 : DFF_X1 port map( D => n3466, CK => CLK, Q => n31135, QN 
                           => n_1711);
   clk_r_REG7568_S1 : DFF_X1 port map( D => n3332, CK => CLK, Q => n31134, QN 
                           => n_1712);
   clk_r_REG7710_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n31133, QN 
                           => n_1713);
   clk_r_REG7712_S1 : DFF_X1 port map( D => n3338, CK => CLK, Q => n31132, QN 
                           => n_1714);
   clk_r_REG7714_S1 : DFF_X1 port map( D => n3337, CK => CLK, Q => n31131, QN 
                           => n_1715);
   clk_r_REG8269_S1 : DFF_X1 port map( D => n3465, CK => CLK, Q => n31130, QN 
                           => n_1716);
   clk_r_REG8271_S1 : DFF_X1 port map( D => n3464, CK => CLK, Q => n31129, QN 
                           => n_1717);
   clk_r_REG7716_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n31128, QN 
                           => n_1718);
   clk_r_REG8273_S1 : DFF_X1 port map( D => n3463, CK => CLK, Q => n31127, QN 
                           => n_1719);
   clk_r_REG8000_S1 : DFF_X1 port map( D => n3374, CK => CLK, Q => n31126, QN 
                           => n_1720);
   clk_r_REG7570_S1 : DFF_X1 port map( D => n3331, CK => CLK, Q => n31125, QN 
                           => n_1721);
   clk_r_REG7718_S1 : DFF_X1 port map( D => n3335, CK => CLK, Q => n31124, QN 
                           => n_1722);
   clk_r_REG7643_S1 : DFF_X1 port map( D => n3365, CK => CLK, Q => n31123, QN 
                           => n_1723);
   clk_r_REG7660_S1 : DFF_X1 port map( D => n3364, CK => CLK, Q => n31122, QN 
                           => n_1724);
   clk_r_REG7662_S1 : DFF_X1 port map( D => n3363, CK => CLK, Q => n31121, QN 
                           => n_1725);
   clk_r_REG8002_S1 : DFF_X1 port map( D => n3373, CK => CLK, Q => n31120, QN 
                           => n_1726);
   clk_r_REG7920_S1 : DFF_X1 port map( D => n3405, CK => CLK, Q => n31119, QN 
                           => n_1727);
   clk_r_REG7664_S1 : DFF_X1 port map( D => n3362, CK => CLK, Q => n31118, QN 
                           => n_1728);
   clk_r_REG9876_S1 : DFF_X1 port map( D => n3437, CK => CLK, Q => n31117, QN 
                           => n_1729);
   clk_r_REG7922_S1 : DFF_X1 port map( D => n3404, CK => CLK, Q => n31116, QN 
                           => n_1730);
   clk_r_REG8004_S1 : DFF_X1 port map( D => n3372, CK => CLK, Q => n31115, QN 
                           => n_1731);
   clk_r_REG8006_S1 : DFF_X1 port map( D => n3371, CK => CLK, Q => n31114, QN 
                           => n_1732);
   clk_r_REG9878_S1 : DFF_X1 port map( D => n3436, CK => CLK, Q => n31113, QN 
                           => n_1733);
   clk_r_REG8008_S1 : DFF_X1 port map( D => n3370, CK => CLK, Q => n31112, QN 
                           => n_1734);
   clk_r_REG8010_S1 : DFF_X1 port map( D => n3369, CK => CLK, Q => n31111, QN 
                           => n_1735);
   clk_r_REG8401_S1 : DFF_X1 port map( D => n3501, CK => CLK, Q => n31110, QN 
                           => n_1736);
   clk_r_REG8012_S1 : DFF_X1 port map( D => n3368, CK => CLK, Q => n31109, QN 
                           => n_1737);
   clk_r_REG8403_S1 : DFF_X1 port map( D => n3500, CK => CLK, Q => n31108, QN 
                           => n_1738);
   clk_r_REG8014_S1 : DFF_X1 port map( D => n3367, CK => CLK, Q => n31107, QN 
                           => n_1739);
   clk_r_REG7924_S1 : DFF_X1 port map( D => n3403, CK => CLK, Q => n31106, QN 
                           => n_1740);
   clk_r_REG9880_S1 : DFF_X1 port map( D => n3435, CK => CLK, Q => n31105, QN 
                           => n_1741);
   clk_r_REG7534_S1 : DFF_X1 port map( D => n3397, CK => CLK, Q => n31104, QN 
                           => n_1742);
   clk_r_REG7956_S1 : DFF_X1 port map( D => n3396, CK => CLK, Q => n31103, QN 
                           => n_1743);
   clk_r_REG7386_S1 : DFF_X1 port map( D => n3493, CK => CLK, Q => n31102, QN 
                           => n_1744);
   clk_r_REG7958_S1 : DFF_X1 port map( D => n3395, CK => CLK, Q => n31101, QN 
                           => n_1745);
   clk_r_REG8405_S1 : DFF_X1 port map( D => n3499, CK => CLK, Q => n31100, QN 
                           => n_1746);
   clk_r_REG7960_S1 : DFF_X1 port map( D => n3394, CK => CLK, Q => n31099, QN 
                           => n_1747);
   clk_r_REG8407_S1 : DFF_X1 port map( D => n3498, CK => CLK, Q => n31098, QN 
                           => n_1748);
   clk_r_REG8215_S1 : DFF_X1 port map( D => n3492, CK => CLK, Q => n31097, QN 
                           => n_1749);
   clk_r_REG9882_S1 : DFF_X1 port map( D => n3434, CK => CLK, Q => n31096, QN 
                           => n_1750);
   clk_r_REG7926_S1 : DFF_X1 port map( D => n3402, CK => CLK, Q => n31095, QN 
                           => n_1751);
   clk_r_REG7928_S1 : DFF_X1 port map( D => n3401, CK => CLK, Q => n31094, QN 
                           => n_1752);
   clk_r_REG7930_S1 : DFF_X1 port map( D => n3400, CK => CLK, Q => n31093, QN 
                           => n_1753);
   clk_r_REG7932_S1 : DFF_X1 port map( D => n3399, CK => CLK, Q => n31092, QN 
                           => n_1754);
   clk_r_REG9884_S1 : DFF_X1 port map( D => n3433, CK => CLK, Q => n31091, QN 
                           => n_1755);
   clk_r_REG9886_S1 : DFF_X1 port map( D => n3432, CK => CLK, Q => n31090, QN 
                           => n_1756);
   clk_r_REG8409_S1 : DFF_X1 port map( D => n3497, CK => CLK, Q => n31089, QN 
                           => n_1757);
   clk_r_REG8411_S1 : DFF_X1 port map( D => n3496, CK => CLK, Q => n31088, QN 
                           => n_1758);
   clk_r_REG7744_S1 : DFF_X1 port map( D => n3429, CK => CLK, Q => n31087, QN 
                           => n_1759);
   clk_r_REG7572_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n31086, QN 
                           => n_1760);
   clk_r_REG8413_S1 : DFF_X1 port map( D => n3495, CK => CLK, Q => n31085, QN 
                           => n_1761);
   clk_r_REG9888_S1 : DFF_X1 port map( D => n3431, CK => CLK, Q => n31084, QN 
                           => n_1762);
   clk_r_REG6936_S1 : DFF_X1 port map( D => n3461, CK => CLK, Q => n31083, QN 
                           => n_1763);
   clk_r_REG8217_S1 : DFF_X1 port map( D => n3491, CK => CLK, Q => n31082, QN 
                           => n_1764);
   clk_r_REG9830_S1 : DFF_X1 port map( D => n3460, CK => CLK, Q => n31081, QN 
                           => n_1765);
   clk_r_REG9832_S1 : DFF_X1 port map( D => n3459, CK => CLK, Q => n31080, QN 
                           => n_1766);
   clk_r_REG8219_S1 : DFF_X1 port map( D => n3490, CK => CLK, Q => n31079, QN 
                           => n_1767);
   clk_r_REG9834_S1 : DFF_X1 port map( D => n3458, CK => CLK, Q => n31078, QN 
                           => n_1768);
   clk_r_REG7310_S1 : DFF_X1 port map( D => n3525, CK => CLK, Q => n31077, QN 
                           => n_1769);
   clk_r_REG7874_S1 : DFF_X1 port map( D => n3428, CK => CLK, Q => n31076, QN 
                           => n_1770);
   clk_r_REG8355_S1 : DFF_X1 port map( D => n3524, CK => CLK, Q => n31075, QN 
                           => n_1771);
   clk_r_REG8357_S1 : DFF_X1 port map( D => n3523, CK => CLK, Q => n31074, QN 
                           => n_1772);
   clk_r_REG8359_S1 : DFF_X1 port map( D => n3522, CK => CLK, Q => n31073, QN 
                           => n_1773);
   clk_r_REG7876_S1 : DFF_X1 port map( D => n3427, CK => CLK, Q => n31072, QN 
                           => n_1774);
   clk_r_REG7878_S1 : DFF_X1 port map( D => n3426, CK => CLK, Q => n31071, QN 
                           => n_1775);
   clk_r_REG7880_S1 : DFF_X1 port map( D => n3425, CK => CLK, Q => n31070, QN 
                           => n_1776);
   clk_r_REG8361_S1 : DFF_X1 port map( D => n3521, CK => CLK, Q => n31069, QN 
                           => n_1777);
   clk_r_REG9836_S1 : DFF_X1 port map( D => n3457, CK => CLK, Q => n31068, QN 
                           => n_1778);
   clk_r_REG7666_S1 : DFF_X1 port map( D => n3361, CK => CLK, Q => n31067, QN 
                           => n_1779);
   clk_r_REG9838_S1 : DFF_X1 port map( D => n3456, CK => CLK, Q => n31066, QN 
                           => n_1780);
   clk_r_REG8221_S1 : DFF_X1 port map( D => n3489, CK => CLK, Q => n31065, QN 
                           => n_1781);
   clk_r_REG8363_S1 : DFF_X1 port map( D => n3520, CK => CLK, Q => n31064, QN 
                           => n_1782);
   clk_r_REG7962_S1 : DFF_X1 port map( D => n3393, CK => CLK, Q => n31063, QN 
                           => n_1783);
   clk_r_REG7964_S1 : DFF_X1 port map( D => n3392, CK => CLK, Q => n31062, QN 
                           => n_1784);
   clk_r_REG7574_S1 : DFF_X1 port map( D => n3329, CK => CLK, Q => n31061, QN 
                           => n_1785);
   clk_r_REG7882_S1 : DFF_X1 port map( D => n3424, CK => CLK, Q => n31060, QN 
                           => n_1786);
   clk_r_REG8223_S1 : DFF_X1 port map( D => n3488, CK => CLK, Q => n31059, QN 
                           => n_1787);
   clk_r_REG7576_S1 : DFF_X1 port map( D => n3328, CK => CLK, Q => n31058, QN 
                           => n_1788);
   clk_r_REG7668_S1 : DFF_X1 port map( D => n3360, CK => CLK, Q => n31057, QN 
                           => n_1789);
   clk_r_REG8365_S1 : DFF_X1 port map( D => n3519, CK => CLK, Q => n31056, QN 
                           => n_1790);
   clk_r_REG7884_S1 : DFF_X1 port map( D => n3423, CK => CLK, Q => n31055, QN 
                           => n_1791);
   clk_r_REG8914_S1 : DFF_X1 port map( D => n2990, CK => CLK, Q => n31054, QN 
                           => n_1792);
   clk_r_REG9809_S1 : DFF_X1 port map( D => n2893, CK => CLK, Q => n31053, QN 
                           => n_1793);
   clk_r_REG7670_S1 : DFF_X1 port map( D => n3359, CK => CLK, Q => n31052, QN 
                           => n_1794);
   clk_r_REG7966_S1 : DFF_X1 port map( D => n3391, CK => CLK, Q => n31051, QN 
                           => n_1795);
   clk_r_REG8531_S1 : DFF_X1 port map( D => n3054, CK => CLK, Q => n31050, QN 
                           => n_1796);
   clk_r_REG8225_S1 : DFF_X1 port map( D => n3487, CK => CLK, Q => n31049, QN 
                           => n_1797);
   clk_r_REG7578_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n31048, QN 
                           => n_1798);
   clk_r_REG9840_S1 : DFF_X1 port map( D => n3455, CK => CLK, Q => n31047, QN 
                           => n_1799);
   clk_r_REG9963_S1 : DFF_X1 port map( D => n3534, CK => CLK, Q => n31046, QN 
                           => n_1800);
   clk_r_REG9965_S1 : DFF_X1 port map( D => n3533, CK => CLK, Q => n31045, QN 
                           => n_1801);
   clk_r_REG9967_S1 : DFF_X1 port map( D => n3532, CK => CLK, Q => n31044, QN 
                           => n_1802);
   clk_r_REG9969_S1 : DFF_X1 port map( D => n3531, CK => CLK, Q => n31043, QN 
                           => n_1803);
   clk_r_REG9971_S1 : DFF_X1 port map( D => n3530, CK => CLK, Q => n31042, QN 
                           => n_1804);
   clk_r_REG9973_S1 : DFF_X1 port map( D => n3529, CK => CLK, Q => n31041, QN 
                           => n_1805);
   clk_r_REG9975_S1 : DFF_X1 port map( D => n3528, CK => CLK, Q => n31040, QN 
                           => n_1806);
   clk_r_REG9977_S1 : DFF_X1 port map( D => n3527, CK => CLK, Q => n31039, QN 
                           => n_1807);
   clk_r_REG6923_S1 : DFF_X1 port map( D => n3557, CK => CLK, Q => n31038, QN 
                           => n_1808);
   clk_r_REG9919_S1 : DFF_X1 port map( D => n3556, CK => CLK, Q => n31037, QN 
                           => n_1809);
   clk_r_REG9921_S1 : DFF_X1 port map( D => n3555, CK => CLK, Q => n31036, QN 
                           => n_1810);
   clk_r_REG7968_S1 : DFF_X1 port map( D => n3390, CK => CLK, Q => n31035, QN 
                           => n_1811);
   clk_r_REG7970_S1 : DFF_X1 port map( D => n3389, CK => CLK, Q => n31034, QN 
                           => n_1812);
   clk_r_REG8367_S1 : DFF_X1 port map( D => n3518, CK => CLK, Q => n31033, QN 
                           => n_1813);
   clk_r_REG7672_S1 : DFF_X1 port map( D => n3358, CK => CLK, Q => n31032, QN 
                           => n_1814);
   clk_r_REG7674_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n31031, QN 
                           => n_1815);
   clk_r_REG7886_S1 : DFF_X1 port map( D => n3422, CK => CLK, Q => n31030, QN 
                           => n_1816);
   clk_r_REG8369_S1 : DFF_X1 port map( D => n3517, CK => CLK, Q => n31029, QN 
                           => n_1817);
   clk_r_REG7888_S1 : DFF_X1 port map( D => n3421, CK => CLK, Q => n31028, QN 
                           => n_1818);
   clk_r_REG8916_S1 : DFF_X1 port map( D => n2989, CK => CLK, Q => n31027, QN 
                           => n_1819);
   clk_r_REG8533_S1 : DFF_X1 port map( D => n3053, CK => CLK, Q => n31026, QN 
                           => n_1820);
   clk_r_REG9842_S1 : DFF_X1 port map( D => n3454, CK => CLK, Q => n31025, QN 
                           => n_1821);
   clk_r_REG8535_S1 : DFF_X1 port map( D => n3052, CK => CLK, Q => n31024, QN 
                           => n_1822);
   clk_r_REG8371_S1 : DFF_X1 port map( D => n3516, CK => CLK, Q => n31023, QN 
                           => n_1823);
   clk_r_REG7580_S1 : DFF_X1 port map( D => n3326, CK => CLK, Q => n31022, QN 
                           => n_1824);
   clk_r_REG7972_S1 : DFF_X1 port map( D => n3388, CK => CLK, Q => n31021, QN 
                           => n_1825);
   clk_r_REG7582_S1 : DFF_X1 port map( D => n3325, CK => CLK, Q => n31020, QN 
                           => n_1826);
   clk_r_REG7890_S1 : DFF_X1 port map( D => n3420, CK => CLK, Q => n31019, QN 
                           => n_1827);
   clk_r_REG9844_S1 : DFF_X1 port map( D => n3453, CK => CLK, Q => n31018, QN 
                           => n_1828);
   clk_r_REG7584_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n31017, QN 
                           => n_1829);
   clk_r_REG7676_S1 : DFF_X1 port map( D => n3356, CK => CLK, Q => n31016, QN 
                           => n_1830);
   clk_r_REG9811_S1 : DFF_X1 port map( D => n2892, CK => CLK, Q => n31015, QN 
                           => n_1831);
   clk_r_REG9846_S1 : DFF_X1 port map( D => n3452, CK => CLK, Q => n31014, QN 
                           => n_1832);
   clk_r_REG8227_S1 : DFF_X1 port map( D => n3486, CK => CLK, Q => n31013, QN 
                           => n_1833);
   clk_r_REG8918_S1 : DFF_X1 port map( D => n2988, CK => CLK, Q => n31012, QN 
                           => n_1834);
   clk_r_REG9813_S1 : DFF_X1 port map( D => n2891, CK => CLK, Q => n31011, QN 
                           => n_1835);
   clk_r_REG8537_S1 : DFF_X1 port map( D => n3051, CK => CLK, Q => n31010, QN 
                           => n_1836);
   clk_r_REG8920_S1 : DFF_X1 port map( D => n2987, CK => CLK, Q => n31009, QN 
                           => n_1837);
   clk_r_REG9815_S1 : DFF_X1 port map( D => n2890, CK => CLK, Q => n31008, QN 
                           => n_1838);
   clk_r_REG8229_S1 : DFF_X1 port map( D => n3485, CK => CLK, Q => n31007, QN 
                           => n_1839);
   clk_r_REG8231_S1 : DFF_X1 port map( D => n3484, CK => CLK, Q => n31006, QN 
                           => n_1840);
   clk_r_REG9617_S1 : DFF_X1 port map( D => n2669, CK => CLK, Q => n31005, QN 
                           => n_1841);
   clk_r_REG9743_S1 : DFF_X1 port map( D => n2734, CK => CLK, Q => n31004, QN 
                           => n_1842);
   clk_r_REG9745_S1 : DFF_X1 port map( D => n2733, CK => CLK, Q => n31003, QN 
                           => n_1843);
   clk_r_REG9747_S1 : DFF_X1 port map( D => n2732, CK => CLK, Q => n31002, QN 
                           => n_1844);
   clk_r_REG9749_S1 : DFF_X1 port map( D => n2731, CK => CLK, Q => n31001, QN 
                           => n_1845);
   clk_r_REG9817_S1 : DFF_X1 port map( D => n2889, CK => CLK, Q => n31000, QN 
                           => n_1846);
   clk_r_REG9751_S1 : DFF_X1 port map( D => n2730, CK => CLK, Q => n30999, QN 
                           => n_1847);
   clk_r_REG9753_S1 : DFF_X1 port map( D => n2729, CK => CLK, Q => n30998, QN 
                           => n_1848);
   clk_r_REG9619_S1 : DFF_X1 port map( D => n2668, CK => CLK, Q => n30997, QN 
                           => n_1849);
   clk_r_REG9755_S1 : DFF_X1 port map( D => n2728, CK => CLK, Q => n30996, QN 
                           => n_1850);
   clk_r_REG9621_S1 : DFF_X1 port map( D => n2667, CK => CLK, Q => n30995, QN 
                           => n_1851);
   clk_r_REG9623_S1 : DFF_X1 port map( D => n2666, CK => CLK, Q => n30994, QN 
                           => n_1852);
   clk_r_REG9425_S1 : DFF_X1 port map( D => n2573, CK => CLK, Q => n30993, QN 
                           => n_1853);
   clk_r_REG9625_S1 : DFF_X1 port map( D => n2665, CK => CLK, Q => n30992, QN 
                           => n_1854);
   clk_r_REG9627_S1 : DFF_X1 port map( D => n2664, CK => CLK, Q => n30991, QN 
                           => n_1855);
   clk_r_REG9629_S1 : DFF_X1 port map( D => n2663, CK => CLK, Q => n30990, QN 
                           => n_1856);
   clk_r_REG9553_S1 : DFF_X1 port map( D => n2637, CK => CLK, Q => n30989, QN 
                           => n_1857);
   clk_r_REG9555_S1 : DFF_X1 port map( D => n2636, CK => CLK, Q => n30988, QN 
                           => n_1858);
   clk_r_REG9557_S1 : DFF_X1 port map( D => n2635, CK => CLK, Q => n30987, QN 
                           => n_1859);
   clk_r_REG9559_S1 : DFF_X1 port map( D => n2634, CK => CLK, Q => n30986, QN 
                           => n_1860);
   clk_r_REG9631_S1 : DFF_X1 port map( D => n2662, CK => CLK, Q => n30985, QN 
                           => n_1861);
   clk_r_REG6973_S1 : DFF_X1 port map( D => n2693, CK => CLK, Q => n30984, QN 
                           => n_1862);
   clk_r_REG9427_S1 : DFF_X1 port map( D => n2572, CK => CLK, Q => n30983, QN 
                           => n_1863);
   clk_r_REG9561_S1 : DFF_X1 port map( D => n2633, CK => CLK, Q => n30982, QN 
                           => n_1864);
   clk_r_REG9563_S1 : DFF_X1 port map( D => n2632, CK => CLK, Q => n30981, QN 
                           => n_1865);
   clk_r_REG9757_S1 : DFF_X1 port map( D => n2727, CK => CLK, Q => n30980, QN 
                           => n_1866);
   clk_r_REG9571_S1 : DFF_X1 port map( D => n2692, CK => CLK, Q => n30979, QN 
                           => n_1867);
   clk_r_REG9429_S1 : DFF_X1 port map( D => n2571, CK => CLK, Q => n30978, QN 
                           => n_1868);
   clk_r_REG9233_S1 : DFF_X1 port map( D => n2797, CK => CLK, Q => n30977, QN 
                           => n_1869);
   clk_r_REG9565_S1 : DFF_X1 port map( D => n2631, CK => CLK, Q => n30976, QN 
                           => n_1870);
   clk_r_REG9567_S1 : DFF_X1 port map( D => n2630, CK => CLK, Q => n30975, QN 
                           => n_1871);
   clk_r_REG6980_S1 : DFF_X1 port map( D => n2661, CK => CLK, Q => n30974, QN 
                           => n_1872);
   clk_r_REG9431_S1 : DFF_X1 port map( D => n2570, CK => CLK, Q => n30973, QN 
                           => n_1873);
   clk_r_REG9507_S1 : DFF_X1 port map( D => n2660, CK => CLK, Q => n30972, QN 
                           => n_1874);
   clk_r_REG9923_S1 : DFF_X1 port map( D => n3554, CK => CLK, Q => n30971, QN 
                           => n_1875);
   clk_r_REG9433_S1 : DFF_X1 port map( D => n2569, CK => CLK, Q => n30970, QN 
                           => n_1876);
   clk_r_REG9435_S1 : DFF_X1 port map( D => n2568, CK => CLK, Q => n30969, QN 
                           => n_1877);
   clk_r_REG9437_S1 : DFF_X1 port map( D => n2567, CK => CLK, Q => n30968, QN 
                           => n_1878);
   clk_r_REG9439_S1 : DFF_X1 port map( D => n2566, CK => CLK, Q => n30967, QN 
                           => n_1879);
   clk_r_REG6996_S1 : DFF_X1 port map( D => n2597, CK => CLK, Q => n30966, QN 
                           => n_1880);
   clk_r_REG9235_S1 : DFF_X1 port map( D => n2796, CK => CLK, Q => n30965, QN 
                           => n_1881);
   clk_r_REG9237_S1 : DFF_X1 port map( D => n2795, CK => CLK, Q => n30964, QN 
                           => n_1882);
   clk_r_REG9379_S1 : DFF_X1 port map( D => n2596, CK => CLK, Q => n30963, QN 
                           => n_1883);
   clk_r_REG9925_S1 : DFF_X1 port map( D => n3553, CK => CLK, Q => n30962, QN 
                           => n_1884);
   clk_r_REG9819_S1 : DFF_X1 port map( D => n2888, CK => CLK, Q => n30961, QN 
                           => n_1885);
   clk_r_REG9239_S1 : DFF_X1 port map( D => n2794, CK => CLK, Q => n30960, QN 
                           => n_1886);
   clk_r_REG6958_S1 : DFF_X1 port map( D => n2757, CK => CLK, Q => n30959, QN 
                           => n_1887);
   clk_r_REG9297_S1 : DFF_X1 port map( D => n2829, CK => CLK, Q => n30958, QN 
                           => n_1888);
   clk_r_REG9927_S1 : DFF_X1 port map( D => n3552, CK => CLK, Q => n30957, QN 
                           => n_1889);
   clk_r_REG9299_S1 : DFF_X1 port map( D => n2828, CK => CLK, Q => n30956, QN 
                           => n_1890);
   clk_r_REG9301_S1 : DFF_X1 port map( D => n2827, CK => CLK, Q => n30955, QN 
                           => n_1891);
   clk_r_REG9303_S1 : DFF_X1 port map( D => n2826, CK => CLK, Q => n30954, QN 
                           => n_1892);
   clk_r_REG9305_S1 : DFF_X1 port map( D => n2825, CK => CLK, Q => n30953, QN 
                           => n_1893);
   clk_r_REG9307_S1 : DFF_X1 port map( D => n2824, CK => CLK, Q => n30952, QN 
                           => n_1894);
   clk_r_REG9241_S1 : DFF_X1 port map( D => n2793, CK => CLK, Q => n30951, QN 
                           => n_1895);
   clk_r_REG9309_S1 : DFF_X1 port map( D => n2823, CK => CLK, Q => n30950, QN 
                           => n_1896);
   clk_r_REG9699_S1 : DFF_X1 port map( D => n2756, CK => CLK, Q => n30949, QN 
                           => n_1897);
   clk_r_REG9311_S1 : DFF_X1 port map( D => n2822, CK => CLK, Q => n30948, QN 
                           => n_1898);
   clk_r_REG9243_S1 : DFF_X1 port map( D => n2792, CK => CLK, Q => n30947, QN 
                           => n_1899);
   clk_r_REG9245_S1 : DFF_X1 port map( D => n2791, CK => CLK, Q => n30946, QN 
                           => n_1900);
   clk_r_REG7019_S1 : DFF_X1 port map( D => n2853, CK => CLK, Q => n30945, QN 
                           => n_1901);
   clk_r_REG9247_S1 : DFF_X1 port map( D => n2790, CK => CLK, Q => n30944, QN 
                           => n_1902);
   clk_r_REG9251_S1 : DFF_X1 port map( D => n2852, CK => CLK, Q => n30943, QN 
                           => n_1903);
   clk_r_REG7027_S1 : DFF_X1 port map( D => n2821, CK => CLK, Q => n30942, QN 
                           => n_1904);
   clk_r_REG9187_S1 : DFF_X1 port map( D => n2820, CK => CLK, Q => n30941, QN 
                           => n_1905);
   clk_r_REG9821_S1 : DFF_X1 port map( D => n2887, CK => CLK, Q => n30940, QN 
                           => n_1906);
   clk_r_REG7586_S1 : DFF_X1 port map( D => n3323, CK => CLK, Q => n30939, QN 
                           => n_1907);
   clk_r_REG9823_S1 : DFF_X1 port map( D => n2886, CK => CLK, Q => n30938, QN 
                           => n_1908);
   clk_r_REG6951_S1 : DFF_X1 port map( D => n2917, CK => CLK, Q => n30937, QN 
                           => n_1909);
   clk_r_REG7588_S1 : DFF_X1 port map( D => n3322, CK => CLK, Q => n30936, QN 
                           => n_1910);
   clk_r_REG7590_S1 : DFF_X1 port map( D => n3321, CK => CLK, Q => n30935, QN 
                           => n_1911);
   clk_r_REG9763_S1 : DFF_X1 port map( D => n2916, CK => CLK, Q => n30934, QN 
                           => n_1912);
   clk_r_REG7592_S1 : DFF_X1 port map( D => n3320, CK => CLK, Q => n30933, QN 
                           => n_1913);
   clk_r_REG9765_S1 : DFF_X1 port map( D => n2915, CK => CLK, Q => n30932, QN 
                           => n_1914);
   clk_r_REG9767_S1 : DFF_X1 port map( D => n2914, CK => CLK, Q => n30931, QN 
                           => n_1915);
   clk_r_REG9769_S1 : DFF_X1 port map( D => n2913, CK => CLK, Q => n30930, QN 
                           => n_1916);
   clk_r_REG9771_S1 : DFF_X1 port map( D => n2912, CK => CLK, Q => n30929, QN 
                           => n_1917);
   clk_r_REG7594_S1 : DFF_X1 port map( D => n3319, CK => CLK, Q => n30928, QN 
                           => n_1918);
   clk_r_REG7596_S1 : DFF_X1 port map( D => n3318, CK => CLK, Q => n30927, QN 
                           => n_1919);
   clk_r_REG7598_S1 : DFF_X1 port map( D => n3317, CK => CLK, Q => n30926, QN 
                           => n_1920);
   clk_r_REG7600_S1 : DFF_X1 port map( D => n3316, CK => CLK, Q => n30925, QN 
                           => n_1921);
   clk_r_REG9929_S1 : DFF_X1 port map( D => n3551, CK => CLK, Q => n30924, QN 
                           => n_1922);
   clk_r_REG9167_S1 : DFF_X1 port map( D => n3214, CK => CLK, Q => n30923, QN 
                           => n_1923);
   clk_r_REG9169_S1 : DFF_X1 port map( D => n3213, CK => CLK, Q => n30922, QN 
                           => n_1924);
   clk_r_REG9171_S1 : DFF_X1 port map( D => n3212, CK => CLK, Q => n30921, QN 
                           => n_1925);
   clk_r_REG9173_S1 : DFF_X1 port map( D => n3211, CK => CLK, Q => n30920, QN 
                           => n_1926);
   clk_r_REG9175_S1 : DFF_X1 port map( D => n3210, CK => CLK, Q => n30919, QN 
                           => n_1927);
   clk_r_REG9177_S1 : DFF_X1 port map( D => n3209, CK => CLK, Q => n30918, QN 
                           => n_1928);
   clk_r_REG9179_S1 : DFF_X1 port map( D => n3208, CK => CLK, Q => n30917, QN 
                           => n_1929);
   clk_r_REG9181_S1 : DFF_X1 port map( D => n3207, CK => CLK, Q => n30916, QN 
                           => n_1930);
   clk_r_REG7046_S1 : DFF_X1 port map( D => n3237, CK => CLK, Q => n30915, QN 
                           => n_1931);
   clk_r_REG9123_S1 : DFF_X1 port map( D => n3236, CK => CLK, Q => n30914, QN 
                           => n_1932);
   clk_r_REG9125_S1 : DFF_X1 port map( D => n3235, CK => CLK, Q => n30913, QN 
                           => n_1933);
   clk_r_REG9931_S1 : DFF_X1 port map( D => n3550, CK => CLK, Q => n30912, QN 
                           => n_1934);
   clk_r_REG9933_S1 : DFF_X1 port map( D => n3549, CK => CLK, Q => n30911, QN 
                           => n_1935);
   clk_r_REG9935_S1 : DFF_X1 port map( D => n3548, CK => CLK, Q => n30910, QN 
                           => n_1936);
   clk_r_REG8661_S1 : DFF_X1 port map( D => n3149, CK => CLK, Q => n30909, QN 
                           => n_1937);
   clk_r_REG8976_S1 : DFF_X1 port map( D => n3023, CK => CLK, Q => n30908, QN 
                           => n_1938);
   clk_r_REG8978_S1 : DFF_X1 port map( D => n3022, CK => CLK, Q => n30907, QN 
                           => n_1939);
   clk_r_REG8467_S1 : DFF_X1 port map( D => n3086, CK => CLK, Q => n30906, QN 
                           => n_1940);
   clk_r_REG8593_S1 : DFF_X1 port map( D => n3119, CK => CLK, Q => n30905, QN 
                           => n_1941);
   clk_r_REG8980_S1 : DFF_X1 port map( D => n3021, CK => CLK, Q => n30904, QN 
                           => n_1942);
   clk_r_REG8539_S1 : DFF_X1 port map( D => n3050, CK => CLK, Q => n30903, QN 
                           => n_1943);
   clk_r_REG8850_S1 : DFF_X1 port map( D => n2958, CK => CLK, Q => n30902, QN 
                           => n_1944);
   clk_r_REG8786_S1 : DFF_X1 port map( D => n2926, CK => CLK, Q => n30901, QN 
                           => n_1945);
   clk_r_REG9773_S1 : DFF_X1 port map( D => n2911, CK => CLK, Q => n30900, QN 
                           => n_1946);
   clk_r_REG8722_S1 : DFF_X1 port map( D => n2862, CK => CLK, Q => n30899, QN 
                           => n_1947);
   clk_r_REG9253_S1 : DFF_X1 port map( D => n2851, CK => CLK, Q => n30898, QN 
                           => n_1948);
   clk_r_REG9189_S1 : DFF_X1 port map( D => n2819, CK => CLK, Q => n30897, QN 
                           => n_1949);
   clk_r_REG9040_S1 : DFF_X1 port map( D => n2766, CK => CLK, Q => n30896, QN 
                           => n_1950);
   clk_r_REG8982_S1 : DFF_X1 port map( D => n3020, CK => CLK, Q => n30895, QN 
                           => n_1951);
   clk_r_REG9701_S1 : DFF_X1 port map( D => n2755, CK => CLK, Q => n30894, QN 
                           => n_1952);
   clk_r_REG8984_S1 : DFF_X1 port map( D => n3019, CK => CLK, Q => n30893, QN 
                           => n_1953);
   clk_r_REG8986_S1 : DFF_X1 port map( D => n3018, CK => CLK, Q => n30892, QN 
                           => n_1954);
   clk_r_REG9465_S1 : DFF_X1 port map( D => n2598, CK => CLK, Q => n30891, QN 
                           => n_1955);
   clk_r_REG8922_S1 : DFF_X1 port map( D => n2986, CK => CLK, Q => n30890, QN 
                           => n_1956);
   clk_r_REG9042_S1 : DFF_X1 port map( D => n2765, CK => CLK, Q => n30889, QN 
                           => n_1957);
   clk_r_REG9044_S1 : DFF_X1 port map( D => n2764, CK => CLK, Q => n30888, QN 
                           => n_1958);
   clk_r_REG8988_S1 : DFF_X1 port map( D => n3017, CK => CLK, Q => n30887, QN 
                           => n_1959);
   clk_r_REG9046_S1 : DFF_X1 port map( D => n2763, CK => CLK, Q => n30886, QN 
                           => n_1960);
   clk_r_REG9048_S1 : DFF_X1 port map( D => n2762, CK => CLK, Q => n30885, QN 
                           => n_1961);
   clk_r_REG9050_S1 : DFF_X1 port map( D => n2761, CK => CLK, Q => n30884, QN 
                           => n_1962);
   clk_r_REG8990_S1 : DFF_X1 port map( D => n3016, CK => CLK, Q => n30883, QN 
                           => n_1963);
   clk_r_REG7118_S1 : DFF_X1 port map( D => n3045, CK => CLK, Q => n30882, QN 
                           => n_1964);
   clk_r_REG8934_S1 : DFF_X1 port map( D => n3044, CK => CLK, Q => n30881, QN 
                           => n_1965);
   clk_r_REG8936_S1 : DFF_X1 port map( D => n3043, CK => CLK, Q => n30880, QN 
                           => n_1966);
   clk_r_REG8938_S1 : DFF_X1 port map( D => n3042, CK => CLK, Q => n30879, QN 
                           => n_1967);
   clk_r_REG8940_S1 : DFF_X1 port map( D => n3041, CK => CLK, Q => n30878, QN 
                           => n_1968);
   clk_r_REG8992_S1 : DFF_X1 port map( D => n3015, CK => CLK, Q => n30877, QN 
                           => n_1969);
   clk_r_REG9052_S1 : DFF_X1 port map( D => n2760, CK => CLK, Q => n30876, QN 
                           => n_1970);
   clk_r_REG9703_S1 : DFF_X1 port map( D => n2754, CK => CLK, Q => n30875, QN 
                           => n_1971);
   clk_r_REG9679_S1 : DFF_X1 port map( D => n2702, CK => CLK, Q => n30874, QN 
                           => n_1972);
   clk_r_REG9573_S1 : DFF_X1 port map( D => n2691, CK => CLK, Q => n30873, QN 
                           => n_1973);
   clk_r_REG9509_S1 : DFF_X1 port map( D => n2659, CK => CLK, Q => n30872, QN 
                           => n_1974);
   clk_r_REG9054_S1 : DFF_X1 port map( D => n2759, CK => CLK, Q => n30871, QN 
                           => n_1975);
   clk_r_REG7106_S1 : DFF_X1 port map( D => n2789, CK => CLK, Q => n30870, QN 
                           => n_1976);
   clk_r_REG8996_S1 : DFF_X1 port map( D => n2788, CK => CLK, Q => n30869, QN 
                           => n_1977);
   clk_r_REG8998_S1 : DFF_X1 port map( D => n2787, CK => CLK, Q => n30868, QN 
                           => n_1978);
   clk_r_REG9000_S1 : DFF_X1 port map( D => n2786, CK => CLK, Q => n30867, QN 
                           => n_1979);
   clk_r_REG9002_S1 : DFF_X1 port map( D => n2785, CK => CLK, Q => n30866, QN 
                           => n_1980);
   clk_r_REG9467_S1 : DFF_X1 port map( D => n2599, CK => CLK, Q => n30865, QN 
                           => n_1981);
   clk_r_REG9381_S1 : DFF_X1 port map( D => n2595, CK => CLK, Q => n30864, QN 
                           => n_1982);
   clk_r_REG9357_S1 : DFF_X1 port map( D => n2542, CK => CLK, Q => n30863, QN 
                           => n_1983);
   clk_r_REG8924_S1 : DFF_X1 port map( D => n2985, CK => CLK, Q => n30862, QN 
                           => n_1984);
   clk_r_REG8926_S1 : DFF_X1 port map( D => n2984, CK => CLK, Q => n30861, QN 
                           => n_1985);
   clk_r_REG8928_S1 : DFF_X1 port map( D => n2983, CK => CLK, Q => n30860, QN 
                           => n_1986);
   clk_r_REG7125_S1 : DFF_X1 port map( D => n3013, CK => CLK, Q => n30859, QN 
                           => n_1987);
   clk_r_REG8870_S1 : DFF_X1 port map( D => n3012, CK => CLK, Q => n30858, QN 
                           => n_1988);
   clk_r_REG8872_S1 : DFF_X1 port map( D => n3011, CK => CLK, Q => n30857, QN 
                           => n_1989);
   clk_r_REG7488_S1 : DFF_X1 port map( D => n3278, CK => CLK, Q => n30856, QN 
                           => n_1990);
   clk_r_REG8323_S1 : DFF_X1 port map( D => n3245, CK => CLK, Q => n30855, QN 
                           => n_1991);
   clk_r_REG8874_S1 : DFF_X1 port map( D => n3010, CK => CLK, Q => n30854, QN 
                           => n_1992);
   clk_r_REG8876_S1 : DFF_X1 port map( D => n3009, CK => CLK, Q => n30853, QN 
                           => n_1993);
   clk_r_REG8878_S1 : DFF_X1 port map( D => n3008, CK => CLK, Q => n30852, QN 
                           => n_1994);
   clk_r_REG8880_S1 : DFF_X1 port map( D => n3007, CK => CLK, Q => n30851, QN 
                           => n_1995);
   clk_r_REG8882_S1 : DFF_X1 port map( D => n3006, CK => CLK, Q => n30850, QN 
                           => n_1996);
   clk_r_REG8884_S1 : DFF_X1 port map( D => n3005, CK => CLK, Q => n30849, QN 
                           => n_1997);
   clk_r_REG7065_S1 : DFF_X1 port map( D => n3174, CK => CLK, Q => n30848, QN 
                           => n_1998);
   clk_r_REG8886_S1 : DFF_X1 port map( D => n3004, CK => CLK, Q => n30847, QN 
                           => n_1999);
   clk_r_REG9127_S1 : DFF_X1 port map( D => n3234, CK => CLK, Q => n30846, QN 
                           => n_2000);
   clk_r_REG9060_S1 : DFF_X1 port map( D => n3175, CK => CLK, Q => n30845, QN 
                           => n_2001);
   clk_r_REG8663_S1 : DFF_X1 port map( D => n3148, CK => CLK, Q => n30844, QN 
                           => n_2002);
   clk_r_REG8595_S1 : DFF_X1 port map( D => n3118, CK => CLK, Q => n30843, QN 
                           => n_2003);
   clk_r_REG9705_S1 : DFF_X1 port map( D => n2753, CK => CLK, Q => n30842, QN 
                           => n_2004);
   clk_r_REG8469_S1 : DFF_X1 port map( D => n3085, CK => CLK, Q => n30841, QN 
                           => n_2005);
   clk_r_REG8541_S1 : DFF_X1 port map( D => n3049, CK => CLK, Q => n30840, QN 
                           => n_2006);
   clk_r_REG8852_S1 : DFF_X1 port map( D => n2957, CK => CLK, Q => n30839, QN 
                           => n_2007);
   clk_r_REG8724_S1 : DFF_X1 port map( D => n2861, CK => CLK, Q => n30838, QN 
                           => n_2008);
   clk_r_REG8726_S1 : DFF_X1 port map( D => n2860, CK => CLK, Q => n30837, QN 
                           => n_2009);
   clk_r_REG8728_S1 : DFF_X1 port map( D => n2859, CK => CLK, Q => n30836, QN 
                           => n_2010);
   clk_r_REG8730_S1 : DFF_X1 port map( D => n2858, CK => CLK, Q => n30835, QN 
                           => n_2011);
   clk_r_REG8732_S1 : DFF_X1 port map( D => n2857, CK => CLK, Q => n30834, QN 
                           => n_2012);
   clk_r_REG8734_S1 : DFF_X1 port map( D => n2856, CK => CLK, Q => n30833, QN 
                           => n_2013);
   clk_r_REG8736_S1 : DFF_X1 port map( D => n2855, CK => CLK, Q => n30832, QN 
                           => n_2014);
   clk_r_REG8788_S1 : DFF_X1 port map( D => n2925, CK => CLK, Q => n30831, QN 
                           => n_2015);
   clk_r_REG9775_S1 : DFF_X1 port map( D => n2910, CK => CLK, Q => n30830, QN 
                           => n_2016);
   clk_r_REG9255_S1 : DFF_X1 port map( D => n2850, CK => CLK, Q => n30829, QN 
                           => n_2017);
   clk_r_REG9191_S1 : DFF_X1 port map( D => n2818, CK => CLK, Q => n30828, QN 
                           => n_2018);
   clk_r_REG7146_S1 : DFF_X1 port map( D => n2885, CK => CLK, Q => n30827, QN 
                           => n_2019);
   clk_r_REG8678_S1 : DFF_X1 port map( D => n2884, CK => CLK, Q => n30826, QN 
                           => n_2020);
   clk_r_REG8680_S1 : DFF_X1 port map( D => n2883, CK => CLK, Q => n30825, QN 
                           => n_2021);
   clk_r_REG8682_S1 : DFF_X1 port map( D => n2882, CK => CLK, Q => n30824, QN 
                           => n_2022);
   clk_r_REG8684_S1 : DFF_X1 port map( D => n2881, CK => CLK, Q => n30823, QN 
                           => n_2023);
   clk_r_REG8686_S1 : DFF_X1 port map( D => n2880, CK => CLK, Q => n30822, QN 
                           => n_2024);
   clk_r_REG9707_S1 : DFF_X1 port map( D => n2752, CK => CLK, Q => n30821, QN 
                           => n_2025);
   clk_r_REG9709_S1 : DFF_X1 port map( D => n2751, CK => CLK, Q => n30820, QN 
                           => n_2026);
   clk_r_REG9711_S1 : DFF_X1 port map( D => n2750, CK => CLK, Q => n30819, QN 
                           => n_2027);
   clk_r_REG9129_S1 : DFF_X1 port map( D => n3233, CK => CLK, Q => n30818, QN 
                           => n_2028);
   clk_r_REG8325_S1 : DFF_X1 port map( D => n3244, CK => CLK, Q => n30817, QN 
                           => n_2029);
   clk_r_REG7490_S1 : DFF_X1 port map( D => n3277, CK => CLK, Q => n30816, QN 
                           => n_2030);
   clk_r_REG9062_S1 : DFF_X1 port map( D => n3176, CK => CLK, Q => n30815, QN 
                           => n_2031);
   clk_r_REG8665_S1 : DFF_X1 port map( D => n3147, CK => CLK, Q => n30814, QN 
                           => n_2032);
   clk_r_REG8597_S1 : DFF_X1 port map( D => n3117, CK => CLK, Q => n30813, QN 
                           => n_2033);
   clk_r_REG8471_S1 : DFF_X1 port map( D => n3084, CK => CLK, Q => n30812, QN 
                           => n_2034);
   clk_r_REG8543_S1 : DFF_X1 port map( D => n3048, CK => CLK, Q => n30811, QN 
                           => n_2035);
   clk_r_REG8854_S1 : DFF_X1 port map( D => n2956, CK => CLK, Q => n30810, QN 
                           => n_2036);
   clk_r_REG8790_S1 : DFF_X1 port map( D => n2924, CK => CLK, Q => n30809, QN 
                           => n_2037);
   clk_r_REG9359_S1 : DFF_X1 port map( D => n2541, CK => CLK, Q => n30808, QN 
                           => n_2038);
   clk_r_REG9383_S1 : DFF_X1 port map( D => n2594, CK => CLK, Q => n30807, QN 
                           => n_2039);
   clk_r_REG9469_S1 : DFF_X1 port map( D => n2600, CK => CLK, Q => n30806, QN 
                           => n_2040);
   clk_r_REG9511_S1 : DFF_X1 port map( D => n2658, CK => CLK, Q => n30805, QN 
                           => n_2041);
   clk_r_REG9575_S1 : DFF_X1 port map( D => n2690, CK => CLK, Q => n30804, QN 
                           => n_2042);
   clk_r_REG9361_S1 : DFF_X1 port map( D => n2540, CK => CLK, Q => n30803, QN 
                           => n_2043);
   clk_r_REG9363_S1 : DFF_X1 port map( D => n2539, CK => CLK, Q => n30802, QN 
                           => n_2044);
   clk_r_REG9365_S1 : DFF_X1 port map( D => n2538, CK => CLK, Q => n30801, QN 
                           => n_2045);
   clk_r_REG9367_S1 : DFF_X1 port map( D => n2537, CK => CLK, Q => n30800, QN 
                           => n_2046);
   clk_r_REG9369_S1 : DFF_X1 port map( D => n2536, CK => CLK, Q => n30799, QN 
                           => n_2047);
   clk_r_REG9371_S1 : DFF_X1 port map( D => n2535, CK => CLK, Q => n30798, QN 
                           => n_2048);
   clk_r_REG7005_S1 : DFF_X1 port map( D => n2565, CK => CLK, Q => n30797, QN 
                           => n_2049);
   clk_r_REG9313_S1 : DFF_X1 port map( D => n2564, CK => CLK, Q => n30796, QN 
                           => n_2050);
   clk_r_REG9315_S1 : DFF_X1 port map( D => n2563, CK => CLK, Q => n30795, QN 
                           => n_2051);
   clk_r_REG9681_S1 : DFF_X1 port map( D => n2701, CK => CLK, Q => n30794, QN 
                           => n_2052);
   clk_r_REG9193_S1 : DFF_X1 port map( D => n2817, CK => CLK, Q => n30793, QN 
                           => n_2053);
   clk_r_REG9317_S1 : DFF_X1 port map( D => n2562, CK => CLK, Q => n30792, QN 
                           => n_2054);
   clk_r_REG9319_S1 : DFF_X1 port map( D => n2561, CK => CLK, Q => n30791, QN 
                           => n_2055);
   clk_r_REG9321_S1 : DFF_X1 port map( D => n2560, CK => CLK, Q => n30790, QN 
                           => n_2056);
   clk_r_REG9257_S1 : DFF_X1 port map( D => n2849, CK => CLK, Q => n30789, QN 
                           => n_2057);
   clk_r_REG9777_S1 : DFF_X1 port map( D => n2909, CK => CLK, Q => n30788, QN 
                           => n_2058);
   clk_r_REG8792_S1 : DFF_X1 port map( D => n2923, CK => CLK, Q => n30787, QN 
                           => n_2059);
   clk_r_REG8856_S1 : DFF_X1 port map( D => n2955, CK => CLK, Q => n30786, QN 
                           => n_2060);
   clk_r_REG8545_S1 : DFF_X1 port map( D => n3047, CK => CLK, Q => n30785, QN 
                           => n_2061);
   clk_r_REG8473_S1 : DFF_X1 port map( D => n3083, CK => CLK, Q => n30784, QN 
                           => n_2062);
   clk_r_REG9683_S1 : DFF_X1 port map( D => n2700, CK => CLK, Q => n30783, QN 
                           => n_2063);
   clk_r_REG9577_S1 : DFF_X1 port map( D => n2689, CK => CLK, Q => n30782, QN 
                           => n_2064);
   clk_r_REG9513_S1 : DFF_X1 port map( D => n2657, CK => CLK, Q => n30781, QN 
                           => n_2065);
   clk_r_REG9471_S1 : DFF_X1 port map( D => n2601, CK => CLK, Q => n30780, QN 
                           => n_2066);
   clk_r_REG9385_S1 : DFF_X1 port map( D => n2593, CK => CLK, Q => n30779, QN 
                           => n_2067);
   clk_r_REG8599_S1 : DFF_X1 port map( D => n3116, CK => CLK, Q => n30778, QN 
                           => n_2068);
   clk_r_REG8667_S1 : DFF_X1 port map( D => n3146, CK => CLK, Q => n30777, QN 
                           => n_2069);
   clk_r_REG9064_S1 : DFF_X1 port map( D => n3177, CK => CLK, Q => n30776, QN 
                           => n_2070);
   clk_r_REG7492_S1 : DFF_X1 port map( D => n3276, CK => CLK, Q => n30775, QN 
                           => n_2071);
   clk_r_REG8327_S1 : DFF_X1 port map( D => n3243, CK => CLK, Q => n30774, QN 
                           => n_2072);
   clk_r_REG9066_S1 : DFF_X1 port map( D => n3178, CK => CLK, Q => n30773, QN 
                           => n_2073);
   clk_r_REG9473_S1 : DFF_X1 port map( D => n2602, CK => CLK, Q => n30772, QN 
                           => n_2074);
   clk_r_REG9475_S1 : DFF_X1 port map( D => n2603, CK => CLK, Q => n30771, QN 
                           => n_2075);
   clk_r_REG8329_S1 : DFF_X1 port map( D => n3242, CK => CLK, Q => n30770, QN 
                           => n_2076);
   clk_r_REG7494_S1 : DFF_X1 port map( D => n3275, CK => CLK, Q => n30769, QN 
                           => n_2077);
   clk_r_REG8669_S1 : DFF_X1 port map( D => n3145, CK => CLK, Q => n30768, QN 
                           => n_2078);
   clk_r_REG8601_S1 : DFF_X1 port map( D => n3115, CK => CLK, Q => n30767, QN 
                           => n_2079);
   clk_r_REG9477_S1 : DFF_X1 port map( D => n2604, CK => CLK, Q => n30766, QN 
                           => n_2080);
   clk_r_REG9479_S1 : DFF_X1 port map( D => n2605, CK => CLK, Q => n30765, QN 
                           => n_2081);
   clk_r_REG8475_S1 : DFF_X1 port map( D => n3082, CK => CLK, Q => n30764, QN 
                           => n_2082);
   clk_r_REG6987_S1 : DFF_X1 port map( D => n2629, CK => CLK, Q => n30763, QN 
                           => n_2083);
   clk_r_REG9443_S1 : DFF_X1 port map( D => n2628, CK => CLK, Q => n30762, QN 
                           => n_2084);
   clk_r_REG9445_S1 : DFF_X1 port map( D => n2627, CK => CLK, Q => n30761, QN 
                           => n_2085);
   clk_r_REG9447_S1 : DFF_X1 port map( D => n2626, CK => CLK, Q => n30760, QN 
                           => n_2086);
   clk_r_REG9449_S1 : DFF_X1 port map( D => n2625, CK => CLK, Q => n30759, QN 
                           => n_2087);
   clk_r_REG9451_S1 : DFF_X1 port map( D => n2624, CK => CLK, Q => n30758, QN 
                           => n_2088);
   clk_r_REG7237_S1 : DFF_X1 port map( D => n3077, CK => CLK, Q => n30757, QN 
                           => n_2089);
   clk_r_REG8858_S1 : DFF_X1 port map( D => n2954, CK => CLK, Q => n30756, QN 
                           => n_2090);
   clk_r_REG8794_S1 : DFF_X1 port map( D => n2922, CK => CLK, Q => n30755, QN 
                           => n_2091);
   clk_r_REG9387_S1 : DFF_X1 port map( D => n2592, CK => CLK, Q => n30754, QN 
                           => n_2092);
   clk_r_REG9389_S1 : DFF_X1 port map( D => n2591, CK => CLK, Q => n30753, QN 
                           => n_2093);
   clk_r_REG9515_S1 : DFF_X1 port map( D => n2656, CK => CLK, Q => n30752, QN 
                           => n_2094);
   clk_r_REG9391_S1 : DFF_X1 port map( D => n2590, CK => CLK, Q => n30751, QN 
                           => n_2095);
   clk_r_REG9393_S1 : DFF_X1 port map( D => n2589, CK => CLK, Q => n30750, QN 
                           => n_2096);
   clk_r_REG9395_S1 : DFF_X1 port map( D => n2588, CK => CLK, Q => n30749, QN 
                           => n_2097);
   clk_r_REG9397_S1 : DFF_X1 port map( D => n2587, CK => CLK, Q => n30748, QN 
                           => n_2098);
   clk_r_REG9713_S1 : DFF_X1 port map( D => n2749, CK => CLK, Q => n30747, QN 
                           => n_2099);
   clk_r_REG9399_S1 : DFF_X1 port map( D => n2586, CK => CLK, Q => n30746, QN 
                           => n_2100);
   clk_r_REG9401_S1 : DFF_X1 port map( D => n2585, CK => CLK, Q => n30745, QN 
                           => n_2101);
   clk_r_REG9685_S1 : DFF_X1 port map( D => n2699, CK => CLK, Q => n30744, QN 
                           => n_2102);
   clk_r_REG9579_S1 : DFF_X1 port map( D => n2688, CK => CLK, Q => n30743, QN 
                           => n_2103);
   clk_r_REG9581_S1 : DFF_X1 port map( D => n2687, CK => CLK, Q => n30742, QN 
                           => n_2104);
   clk_r_REG9583_S1 : DFF_X1 port map( D => n2686, CK => CLK, Q => n30741, QN 
                           => n_2105);
   clk_r_REG9585_S1 : DFF_X1 port map( D => n2685, CK => CLK, Q => n30740, QN 
                           => n_2106);
   clk_r_REG9587_S1 : DFF_X1 port map( D => n2684, CK => CLK, Q => n30739, QN 
                           => n_2107);
   clk_r_REG9589_S1 : DFF_X1 port map( D => n2683, CK => CLK, Q => n30738, QN 
                           => n_2108);
   clk_r_REG9591_S1 : DFF_X1 port map( D => n2682, CK => CLK, Q => n30737, QN 
                           => n_2109);
   clk_r_REG9593_S1 : DFF_X1 port map( D => n2681, CK => CLK, Q => n30736, QN 
                           => n_2110);
   clk_r_REG9517_S1 : DFF_X1 port map( D => n2655, CK => CLK, Q => n30735, QN 
                           => n_2111);
   clk_r_REG7496_S1 : DFF_X1 port map( D => n3274, CK => CLK, Q => n30734, QN 
                           => n_2112);
   clk_r_REG9519_S1 : DFF_X1 port map( D => n2654, CK => CLK, Q => n30733, QN 
                           => n_2113);
   clk_r_REG8331_S1 : DFF_X1 port map( D => n3241, CK => CLK, Q => n30732, QN 
                           => n_2114);
   clk_r_REG9521_S1 : DFF_X1 port map( D => n2653, CK => CLK, Q => n30731, QN 
                           => n_2115);
   clk_r_REG9131_S1 : DFF_X1 port map( D => n3232, CK => CLK, Q => n30730, QN 
                           => n_2116);
   clk_r_REG9523_S1 : DFF_X1 port map( D => n2652, CK => CLK, Q => n30729, QN 
                           => n_2117);
   clk_r_REG9525_S1 : DFF_X1 port map( D => n2651, CK => CLK, Q => n30728, QN 
                           => n_2118);
   clk_r_REG9068_S1 : DFF_X1 port map( D => n3179, CK => CLK, Q => n30727, QN 
                           => n_2119);
   clk_r_REG8671_S1 : DFF_X1 port map( D => n3144, CK => CLK, Q => n30726, QN 
                           => n_2120);
   clk_r_REG8603_S1 : DFF_X1 port map( D => n3114, CK => CLK, Q => n30725, QN 
                           => n_2121);
   clk_r_REG8477_S1 : DFF_X1 port map( D => n3081, CK => CLK, Q => n30724, QN 
                           => n_2122);
   clk_r_REG9527_S1 : DFF_X1 port map( D => n2650, CK => CLK, Q => n30723, QN 
                           => n_2123);
   clk_r_REG9529_S1 : DFF_X1 port map( D => n2649, CK => CLK, Q => n30722, QN 
                           => n_2124);
   clk_r_REG8487_S1 : DFF_X1 port map( D => n3076, CK => CLK, Q => n30721, QN 
                           => n_2125);
   clk_r_REG8860_S1 : DFF_X1 port map( D => n2953, CK => CLK, Q => n30720, QN 
                           => n_2126);
   clk_r_REG9687_S1 : DFF_X1 port map( D => n2698, CK => CLK, Q => n30719, QN 
                           => n_2127);
   clk_r_REG8796_S1 : DFF_X1 port map( D => n2921, CK => CLK, Q => n30718, QN 
                           => n_2128);
   clk_r_REG9779_S1 : DFF_X1 port map( D => n2908, CK => CLK, Q => n30717, QN 
                           => n_2129);
   clk_r_REG9259_S1 : DFF_X1 port map( D => n2848, CK => CLK, Q => n30716, QN 
                           => n_2130);
   clk_r_REG9195_S1 : DFF_X1 port map( D => n2816, CK => CLK, Q => n30715, QN 
                           => n_2131);
   clk_r_REG9261_S1 : DFF_X1 port map( D => n2847, CK => CLK, Q => n30714, QN 
                           => n_2132);
   clk_r_REG9781_S1 : DFF_X1 port map( D => n2907, CK => CLK, Q => n30713, QN 
                           => n_2133);
   clk_r_REG8798_S1 : DFF_X1 port map( D => n2920, CK => CLK, Q => n30712, QN 
                           => n_2134);
   clk_r_REG9689_S1 : DFF_X1 port map( D => n2697, CK => CLK, Q => n30711, QN 
                           => n_2135);
   clk_r_REG9197_S1 : DFF_X1 port map( D => n2815, CK => CLK, Q => n30710, QN 
                           => n_2136);
   clk_r_REG9691_S1 : DFF_X1 port map( D => n2696, CK => CLK, Q => n30709, QN 
                           => n_2137);
   clk_r_REG9693_S1 : DFF_X1 port map( D => n2695, CK => CLK, Q => n30708, QN 
                           => n_2138);
   clk_r_REG6966_S1 : DFF_X1 port map( D => n2725, CK => CLK, Q => n30707, QN 
                           => n_2139);
   clk_r_REG9635_S1 : DFF_X1 port map( D => n2724, CK => CLK, Q => n30706, QN 
                           => n_2140);
   clk_r_REG9637_S1 : DFF_X1 port map( D => n2723, CK => CLK, Q => n30705, QN 
                           => n_2141);
   clk_r_REG9639_S1 : DFF_X1 port map( D => n2722, CK => CLK, Q => n30704, QN 
                           => n_2142);
   clk_r_REG9641_S1 : DFF_X1 port map( D => n2721, CK => CLK, Q => n30703, QN 
                           => n_2143);
   clk_r_REG8862_S1 : DFF_X1 port map( D => n2952, CK => CLK, Q => n30702, QN 
                           => n_2144);
   clk_r_REG8489_S1 : DFF_X1 port map( D => n3075, CK => CLK, Q => n30701, QN 
                           => n_2145);
   clk_r_REG9643_S1 : DFF_X1 port map( D => n2720, CK => CLK, Q => n30700, QN 
                           => n_2146);
   clk_r_REG8479_S1 : DFF_X1 port map( D => n3080, CK => CLK, Q => n30699, QN 
                           => n_2147);
   clk_r_REG8605_S1 : DFF_X1 port map( D => n3113, CK => CLK, Q => n30698, QN 
                           => n_2148);
   clk_r_REG8673_S1 : DFF_X1 port map( D => n3143, CK => CLK, Q => n30697, QN 
                           => n_2149);
   clk_r_REG9070_S1 : DFF_X1 port map( D => n3180, CK => CLK, Q => n30696, QN 
                           => n_2150);
   clk_r_REG9133_S1 : DFF_X1 port map( D => n3231, CK => CLK, Q => n30695, QN 
                           => n_2151);
   clk_r_REG8333_S1 : DFF_X1 port map( D => n3240, CK => CLK, Q => n30694, QN 
                           => n_2152);
   clk_r_REG7498_S1 : DFF_X1 port map( D => n3273, CK => CLK, Q => n30693, QN 
                           => n_2153);
   clk_r_REG9715_S1 : DFF_X1 port map( D => n2748, CK => CLK, Q => n30692, QN 
                           => n_2154);
   clk_r_REG9717_S1 : DFF_X1 port map( D => n2747, CK => CLK, Q => n30691, QN 
                           => n_2155);
   clk_r_REG9719_S1 : DFF_X1 port map( D => n2746, CK => CLK, Q => n30690, QN 
                           => n_2156);
   clk_r_REG9721_S1 : DFF_X1 port map( D => n2745, CK => CLK, Q => n30689, QN 
                           => n_2157);
   clk_r_REG8335_S1 : DFF_X1 port map( D => n3239, CK => CLK, Q => n30688, QN 
                           => n_2158);
   clk_r_REG9135_S1 : DFF_X1 port map( D => n3230, CK => CLK, Q => n30687, QN 
                           => n_2159);
   clk_r_REG9137_S1 : DFF_X1 port map( D => n3229, CK => CLK, Q => n30686, QN 
                           => n_2160);
   clk_r_REG9139_S1 : DFF_X1 port map( D => n3228, CK => CLK, Q => n30685, QN 
                           => n_2161);
   clk_r_REG9141_S1 : DFF_X1 port map( D => n3227, CK => CLK, Q => n30684, QN 
                           => n_2162);
   clk_r_REG9143_S1 : DFF_X1 port map( D => n3226, CK => CLK, Q => n30683, QN 
                           => n_2163);
   clk_r_REG9183_S1 : DFF_X1 port map( D => n3206, CK => CLK, Q => n30682, QN 
                           => n_2164);
   clk_r_REG7500_S1 : DFF_X1 port map( D => n3272, CK => CLK, Q => n30681, QN 
                           => n_2165);
   clk_r_REG8337_S1 : DFF_X1 port map( D => n3238, CK => CLK, Q => n30680, QN 
                           => n_2166);
   clk_r_REG9072_S1 : DFF_X1 port map( D => n3181, CK => CLK, Q => n30679, QN 
                           => n_2167);
   clk_r_REG9074_S1 : DFF_X1 port map( D => n3205, CK => CLK, Q => n30678, QN 
                           => n_2168);
   clk_r_REG9076_S1 : DFF_X1 port map( D => n3204, CK => CLK, Q => n30677, QN 
                           => n_2169);
   clk_r_REG9078_S1 : DFF_X1 port map( D => n3203, CK => CLK, Q => n30676, QN 
                           => n_2170);
   clk_r_REG9080_S1 : DFF_X1 port map( D => n3202, CK => CLK, Q => n30675, QN 
                           => n_2171);
   clk_r_REG9082_S1 : DFF_X1 port map( D => n3201, CK => CLK, Q => n30674, QN 
                           => n_2172);
   clk_r_REG9084_S1 : DFF_X1 port map( D => n3200, CK => CLK, Q => n30673, QN 
                           => n_2173);
   clk_r_REG8675_S1 : DFF_X1 port map( D => n3142, CK => CLK, Q => n30672, QN 
                           => n_2174);
   clk_r_REG8607_S1 : DFF_X1 port map( D => n3112, CK => CLK, Q => n30671, QN 
                           => n_2175);
   clk_r_REG8481_S1 : DFF_X1 port map( D => n3079, CK => CLK, Q => n30670, QN 
                           => n_2176);
   clk_r_REG8491_S1 : DFF_X1 port map( D => n3074, CK => CLK, Q => n30669, QN 
                           => n_2177);
   clk_r_REG8864_S1 : DFF_X1 port map( D => n2951, CK => CLK, Q => n30668, QN 
                           => n_2178);
   clk_r_REG8800_S1 : DFF_X1 port map( D => n2919, CK => CLK, Q => n30667, QN 
                           => n_2179);
   clk_r_REG9783_S1 : DFF_X1 port map( D => n2906, CK => CLK, Q => n30666, QN 
                           => n_2180);
   clk_r_REG9263_S1 : DFF_X1 port map( D => n2846, CK => CLK, Q => n30665, QN 
                           => n_2181);
   clk_r_REG7168_S1 : DFF_X1 port map( D => n3173, CK => CLK, Q => n30664, QN 
                           => n_2182);
   clk_r_REG8615_S1 : DFF_X1 port map( D => n3172, CK => CLK, Q => n30663, QN 
                           => n_2183);
   clk_r_REG8617_S1 : DFF_X1 port map( D => n3171, CK => CLK, Q => n30662, QN 
                           => n_2184);
   clk_r_REG8619_S1 : DFF_X1 port map( D => n3170, CK => CLK, Q => n30661, QN 
                           => n_2185);
   clk_r_REG8621_S1 : DFF_X1 port map( D => n3169, CK => CLK, Q => n30660, QN 
                           => n_2186);
   clk_r_REG8623_S1 : DFF_X1 port map( D => n3168, CK => CLK, Q => n30659, QN 
                           => n_2187);
   clk_r_REG9199_S1 : DFF_X1 port map( D => n2814, CK => CLK, Q => n30658, QN 
                           => n_2188);
   clk_r_REG7186_S1 : DFF_X1 port map( D => n3141, CK => CLK, Q => n30657, QN 
                           => n_2189);
   clk_r_REG8551_S1 : DFF_X1 port map( D => n3140, CK => CLK, Q => n30656, QN 
                           => n_2190);
   clk_r_REG8553_S1 : DFF_X1 port map( D => n3139, CK => CLK, Q => n30655, QN 
                           => n_2191);
   clk_r_REG8555_S1 : DFF_X1 port map( D => n3138, CK => CLK, Q => n30654, QN 
                           => n_2192);
   clk_r_REG8557_S1 : DFF_X1 port map( D => n3137, CK => CLK, Q => n30653, QN 
                           => n_2193);
   clk_r_REG8609_S1 : DFF_X1 port map( D => n3111, CK => CLK, Q => n30652, QN 
                           => n_2194);
   clk_r_REG7502_S1 : DFF_X1 port map( D => n3271, CK => CLK, Q => n30651, QN 
                           => n_2195);
   clk_r_REG7329_S1 : DFF_X1 port map( D => n3269, CK => CLK, Q => n30650, QN 
                           => n_2196);
   clk_r_REG7256_S1 : DFF_X1 port map( D => n3109, CK => CLK, Q => n30649, QN 
                           => n_2197);
   clk_r_REG8493_S1 : DFF_X1 port map( D => n3073, CK => CLK, Q => n30648, QN 
                           => n_2198);
   clk_r_REG8495_S1 : DFF_X1 port map( D => n3072, CK => CLK, Q => n30647, QN 
                           => n_2199);
   clk_r_REG8497_S1 : DFF_X1 port map( D => n3071, CK => CLK, Q => n30646, QN 
                           => n_2200);
   clk_r_REG8499_S1 : DFF_X1 port map( D => n3070, CK => CLK, Q => n30645, QN 
                           => n_2201);
   clk_r_REG8501_S1 : DFF_X1 port map( D => n3069, CK => CLK, Q => n30644, QN 
                           => n_2202);
   clk_r_REG8503_S1 : DFF_X1 port map( D => n3068, CK => CLK, Q => n30643, QN 
                           => n_2203);
   clk_r_REG9145_S1 : DFF_X1 port map( D => n3225, CK => CLK, Q => n30642, QN 
                           => n_2204);
   clk_r_REG8277_S1 : DFF_X1 port map( D => n3268, CK => CLK, Q => n30641, QN 
                           => n_2205);
   clk_r_REG8279_S1 : DFF_X1 port map( D => n3267, CK => CLK, Q => n30640, QN 
                           => n_2206);
   clk_r_REG8281_S1 : DFF_X1 port map( D => n3266, CK => CLK, Q => n30639, QN 
                           => n_2207);
   clk_r_REG8283_S1 : DFF_X1 port map( D => n3265, CK => CLK, Q => n30638, QN 
                           => n_2208);
   clk_r_REG8285_S1 : DFF_X1 port map( D => n3264, CK => CLK, Q => n30637, QN 
                           => n_2209);
   clk_r_REG9201_S1 : DFF_X1 port map( D => n2813, CK => CLK, Q => n30636, QN 
                           => n_2210);
   clk_r_REG9265_S1 : DFF_X1 port map( D => n2845, CK => CLK, Q => n30635, QN 
                           => n_2211);
   clk_r_REG9785_S1 : DFF_X1 port map( D => n2905, CK => CLK, Q => n30634, QN 
                           => n_2212);
   clk_r_REG7139_S1 : DFF_X1 port map( D => n2949, CK => CLK, Q => n30633, QN 
                           => n_2213);
   clk_r_REG7132_S1 : DFF_X1 port map( D => n2981, CK => CLK, Q => n30632, QN 
                           => n_2214);
   clk_r_REG7399_S1 : DFF_X1 port map( D => n3301, CK => CLK, Q => n30631, QN 
                           => n_2215);
   clk_r_REG7444_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n30630, QN 
                           => n_2216);
   clk_r_REG7446_S1 : DFF_X1 port map( D => n3299, CK => CLK, Q => n30629, QN 
                           => n_2217);
   clk_r_REG8423_S1 : DFF_X1 port map( D => n3108, CK => CLK, Q => n30628, QN 
                           => n_2218);
   clk_r_REG7448_S1 : DFF_X1 port map( D => n3298, CK => CLK, Q => n30627, QN 
                           => n_2219);
   clk_r_REG7450_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n30626, QN 
                           => n_2220);
   clk_r_REG7452_S1 : DFF_X1 port map( D => n3296, CK => CLK, Q => n30625, QN 
                           => n_2221);
   clk_r_REG9203_S1 : DFF_X1 port map( D => n2812, CK => CLK, Q => n30624, QN 
                           => n_2222);
   clk_r_REG9267_S1 : DFF_X1 port map( D => n2844, CK => CLK, Q => n30623, QN 
                           => n_2223);
   clk_r_REG9787_S1 : DFF_X1 port map( D => n2904, CK => CLK, Q => n30622, QN 
                           => n_2224);
   clk_r_REG8742_S1 : DFF_X1 port map( D => n2948, CK => CLK, Q => n30621, QN 
                           => n_2225);
   clk_r_REG8806_S1 : DFF_X1 port map( D => n2980, CK => CLK, Q => n30620, QN 
                           => n_2226);
   clk_r_REG8425_S1 : DFF_X1 port map( D => n3107, CK => CLK, Q => n30619, QN 
                           => n_2227);
   clk_r_REG9004_S1 : DFF_X1 port map( D => n2784, CK => CLK, Q => n30618, QN 
                           => n_2228);
   clk_r_REG9205_S1 : DFF_X1 port map( D => n2811, CK => CLK, Q => n30617, QN 
                           => n_2229);
   clk_r_REG9269_S1 : DFF_X1 port map( D => n2843, CK => CLK, Q => n30616, QN 
                           => n_2230);
   clk_r_REG9789_S1 : DFF_X1 port map( D => n2903, CK => CLK, Q => n30615, QN 
                           => n_2231);
   clk_r_REG8744_S1 : DFF_X1 port map( D => n2947, CK => CLK, Q => n30614, QN 
                           => n_2232);
   clk_r_REG8808_S1 : DFF_X1 port map( D => n2979, CK => CLK, Q => n30613, QN 
                           => n_2233);
   clk_r_REG8427_S1 : DFF_X1 port map( D => n3106, CK => CLK, Q => n30612, QN 
                           => n_2234);
   clk_r_REG8810_S1 : DFF_X1 port map( D => n2978, CK => CLK, Q => n30611, QN 
                           => n_2235);
   clk_r_REG8812_S1 : DFF_X1 port map( D => n2977, CK => CLK, Q => n30610, QN 
                           => n_2236);
   clk_r_REG8814_S1 : DFF_X1 port map( D => n2976, CK => CLK, Q => n30609, QN 
                           => n_2237);
   clk_r_REG9271_S1 : DFF_X1 port map( D => n2842, CK => CLK, Q => n30608, QN 
                           => n_2238);
   clk_r_REG9273_S1 : DFF_X1 port map( D => n2841, CK => CLK, Q => n30607, QN 
                           => n_2239);
   clk_r_REG9275_S1 : DFF_X1 port map( D => n2840, CK => CLK, Q => n30606, QN 
                           => n_2240);
   clk_r_REG9207_S1 : DFF_X1 port map( D => n2810, CK => CLK, Q => n30605, QN 
                           => n_2241);
   clk_r_REG9209_S1 : DFF_X1 port map( D => n2809, CK => CLK, Q => n30604, QN 
                           => n_2242);
   clk_r_REG9211_S1 : DFF_X1 port map( D => n2808, CK => CLK, Q => n30603, QN 
                           => n_2243);
   clk_r_REG9791_S1 : DFF_X1 port map( D => n2902, CK => CLK, Q => n30602, QN 
                           => n_2244);
   clk_r_REG8746_S1 : DFF_X1 port map( D => n2946, CK => CLK, Q => n30601, QN 
                           => n_2245);
   clk_r_REG8748_S1 : DFF_X1 port map( D => n2945, CK => CLK, Q => n30600, QN 
                           => n_2246);
   clk_r_REG8750_S1 : DFF_X1 port map( D => n2944, CK => CLK, Q => n30599, QN 
                           => n_2247);
   clk_r_REG8429_S1 : DFF_X1 port map( D => n3105, CK => CLK, Q => n30598, QN 
                           => n_2248);
   clk_r_REG9793_S1 : DFF_X1 port map( D => n2901, CK => CLK, Q => n30597, QN 
                           => n_2249);
   clk_r_REG9795_S1 : DFF_X1 port map( D => n2900, CK => CLK, Q => n30596, QN 
                           => n_2250);
   clk_r_REG8431_S1 : DFF_X1 port map( D => n3104, CK => CLK, Q => n30595, QN 
                           => n_2251);
   clk_r_REG8433_S1 : DFF_X1 port map( D => n3103, CK => CLK, Q => n30594, QN 
                           => n_2252);
   clk_r_REG9323_S1 : DFF_X1 port map( D => n2559, CK => CLK, Q => n30593, QN 
                           => n_2253);
   clk_r_REG8287_S1 : DFF_X1 port map( D => n3263, CK => CLK, Q => n30592, QN 
                           => n_2254);
   clk_r_REG9213_S1 : DFF_X1 port map( D => n2807, CK => CLK, Q => n30591, QN 
                           => n_2255);
   clk_r_REG7454_S1 : DFF_X1 port map( D => n3295, CK => CLK, Q => n30590, QN 
                           => n_2256);
   clk_r_REG9531_S1 : DFF_X1 port map( D => n2648, CK => CLK, Q => n30589, QN 
                           => n_2257);
   clk_r_REG8816_S1 : DFF_X1 port map( D => n2975, CK => CLK, Q => n30588, QN 
                           => n_2258);
   clk_r_REG8559_S1 : DFF_X1 port map( D => n3136, CK => CLK, Q => n30587, QN 
                           => n_2259);
   clk_r_REG8942_S1 : DFF_X1 port map( D => n3040, CK => CLK, Q => n30586, QN 
                           => n_2260);
   clk_r_REG9645_S1 : DFF_X1 port map( D => n2719, CK => CLK, Q => n30585, QN 
                           => n_2261);
   clk_r_REG9006_S1 : DFF_X1 port map( D => n2783, CK => CLK, Q => n30584, QN 
                           => n_2262);
   clk_r_REG9277_S1 : DFF_X1 port map( D => n2839, CK => CLK, Q => n30583, QN 
                           => n_2263);
   clk_r_REG9147_S1 : DFF_X1 port map( D => n3224, CK => CLK, Q => n30582, QN 
                           => n_2264);
   clk_r_REG8688_S1 : DFF_X1 port map( D => n2879, CK => CLK, Q => n30581, QN 
                           => n_2265);
   clk_r_REG9086_S1 : DFF_X1 port map( D => n3199, CK => CLK, Q => n30580, QN 
                           => n_2266);
   clk_r_REG8625_S1 : DFF_X1 port map( D => n3167, CK => CLK, Q => n30579, QN 
                           => n_2267);
   clk_r_REG9723_S1 : DFF_X1 port map( D => n2744, CK => CLK, Q => n30578, QN 
                           => n_2268);
   clk_r_REG9453_S1 : DFF_X1 port map( D => n2623, CK => CLK, Q => n30577, QN 
                           => n_2269);
   clk_r_REG8752_S1 : DFF_X1 port map( D => n2943, CK => CLK, Q => n30576, QN 
                           => n_2270);
   clk_r_REG9595_S1 : DFF_X1 port map( D => n2680, CK => CLK, Q => n30575, QN 
                           => n_2271);
   clk_r_REG9403_S1 : DFF_X1 port map( D => n2584, CK => CLK, Q => n30574, QN 
                           => n_2272);
   clk_r_REG9405_S1 : DFF_X1 port map( D => n2583, CK => CLK, Q => n30573, QN 
                           => n_2273);
   clk_r_REG9759_S1 : DFF_X1 port map( D => n2726, CK => CLK, Q => n30572, QN 
                           => n_2274);
   clk_r_REG9797_S1 : DFF_X1 port map( D => n2899, CK => CLK, Q => n30571, QN 
                           => n_2275);
   clk_r_REG9799_S1 : DFF_X1 port map( D => n2898, CK => CLK, Q => n30570, QN 
                           => n_2276);
   clk_r_REG9801_S1 : DFF_X1 port map( D => n2897, CK => CLK, Q => n30569, QN 
                           => n_2277);
   clk_r_REG9407_S1 : DFF_X1 port map( D => n2582, CK => CLK, Q => n30568, QN 
                           => n_2278);
   clk_r_REG9725_S1 : DFF_X1 port map( D => n2743, CK => CLK, Q => n30567, QN 
                           => n_2279);
   clk_r_REG9597_S1 : DFF_X1 port map( D => n2679, CK => CLK, Q => n30566, QN 
                           => n_2280);
   clk_r_REG9215_S1 : DFF_X1 port map( D => n2806, CK => CLK, Q => n30565, QN 
                           => n_2281);
   clk_r_REG9533_S1 : DFF_X1 port map( D => n2647, CK => CLK, Q => n30564, QN 
                           => n_2282);
   clk_r_REG9217_S1 : DFF_X1 port map( D => n2805, CK => CLK, Q => n30563, QN 
                           => n_2283);
   clk_r_REG9219_S1 : DFF_X1 port map( D => n2804, CK => CLK, Q => n30562, QN 
                           => n_2284);
   clk_r_REG9409_S1 : DFF_X1 port map( D => n2581, CK => CLK, Q => n30561, QN 
                           => n_2285);
   clk_r_REG9727_S1 : DFF_X1 port map( D => n2742, CK => CLK, Q => n30560, QN 
                           => n_2286);
   clk_r_REG9279_S1 : DFF_X1 port map( D => n2838, CK => CLK, Q => n30559, QN 
                           => n_2287);
   clk_r_REG9535_S1 : DFF_X1 port map( D => n2646, CK => CLK, Q => n30558, QN 
                           => n_2288);
   clk_r_REG9411_S1 : DFF_X1 port map( D => n2580, CK => CLK, Q => n30557, QN 
                           => n_2289);
   clk_r_REG9803_S1 : DFF_X1 port map( D => n2896, CK => CLK, Q => n30556, QN 
                           => n_2290);
   clk_r_REG9599_S1 : DFF_X1 port map( D => n2678, CK => CLK, Q => n30555, QN 
                           => n_2291);
   clk_r_REG9537_S1 : DFF_X1 port map( D => n2645, CK => CLK, Q => n30554, QN 
                           => n_2292);
   clk_r_REG9539_S1 : DFF_X1 port map( D => n2644, CK => CLK, Q => n30553, QN 
                           => n_2293);
   clk_r_REG9281_S1 : DFF_X1 port map( D => n2837, CK => CLK, Q => n30552, QN 
                           => n_2294);
   clk_r_REG9221_S1 : DFF_X1 port map( D => n2803, CK => CLK, Q => n30551, QN 
                           => n_2295);
   clk_r_REG9729_S1 : DFF_X1 port map( D => n2741, CK => CLK, Q => n30550, QN 
                           => n_2296);
   clk_r_REG9601_S1 : DFF_X1 port map( D => n2677, CK => CLK, Q => n30549, QN 
                           => n_2297);
   clk_r_REG9731_S1 : DFF_X1 port map( D => n2740, CK => CLK, Q => n30548, QN 
                           => n_2298);
   clk_r_REG9603_S1 : DFF_X1 port map( D => n2676, CK => CLK, Q => n30547, QN 
                           => n_2299);
   clk_r_REG9541_S1 : DFF_X1 port map( D => n2643, CK => CLK, Q => n30546, QN 
                           => n_2300);
   clk_r_REG9413_S1 : DFF_X1 port map( D => n2579, CK => CLK, Q => n30545, QN 
                           => n_2301);
   clk_r_REG9805_S1 : DFF_X1 port map( D => n2895, CK => CLK, Q => n30544, QN 
                           => n_2302);
   clk_r_REG9283_S1 : DFF_X1 port map( D => n2836, CK => CLK, Q => n30543, QN 
                           => n_2303);
   clk_r_REG9285_S1 : DFF_X1 port map( D => n2835, CK => CLK, Q => n30542, QN 
                           => n_2304);
   clk_r_REG9605_S1 : DFF_X1 port map( D => n2675, CK => CLK, Q => n30541, QN 
                           => n_2305);
   clk_r_REG9543_S1 : DFF_X1 port map( D => n2642, CK => CLK, Q => n30540, QN 
                           => n_2306);
   clk_r_REG9733_S1 : DFF_X1 port map( D => n2739, CK => CLK, Q => n30539, QN 
                           => n_2307);
   clk_r_REG9607_S1 : DFF_X1 port map( D => n2674, CK => CLK, Q => n30538, QN 
                           => n_2308);
   clk_r_REG9545_S1 : DFF_X1 port map( D => n2641, CK => CLK, Q => n30537, QN 
                           => n_2309);
   clk_r_REG9415_S1 : DFF_X1 port map( D => n2578, CK => CLK, Q => n30536, QN 
                           => n_2310);
   clk_r_REG9735_S1 : DFF_X1 port map( D => n2738, CK => CLK, Q => n30535, QN 
                           => n_2311);
   clk_r_REG9609_S1 : DFF_X1 port map( D => n2673, CK => CLK, Q => n30534, QN 
                           => n_2312);
   clk_r_REG9547_S1 : DFF_X1 port map( D => n2640, CK => CLK, Q => n30533, QN 
                           => n_2313);
   clk_r_REG9417_S1 : DFF_X1 port map( D => n2577, CK => CLK, Q => n30532, QN 
                           => n_2314);
   clk_r_REG9807_S1 : DFF_X1 port map( D => n2894, CK => CLK, Q => n30531, QN 
                           => n_2315);
   clk_r_REG9287_S1 : DFF_X1 port map( D => n2834, CK => CLK, Q => n30530, QN 
                           => n_2316);
   clk_r_REG9289_S1 : DFF_X1 port map( D => n2833, CK => CLK, Q => n30529, QN 
                           => n_2317);
   clk_r_REG9223_S1 : DFF_X1 port map( D => n2802, CK => CLK, Q => n30528, QN 
                           => n_2318);
   clk_r_REG9737_S1 : DFF_X1 port map( D => n2737, CK => CLK, Q => n30527, QN 
                           => n_2319);
   clk_r_REG9611_S1 : DFF_X1 port map( D => n2672, CK => CLK, Q => n30526, QN 
                           => n_2320);
   clk_r_REG9549_S1 : DFF_X1 port map( D => n2639, CK => CLK, Q => n30525, QN 
                           => n_2321);
   clk_r_REG9419_S1 : DFF_X1 port map( D => n2576, CK => CLK, Q => n30524, QN 
                           => n_2322);
   clk_r_REG9225_S1 : DFF_X1 port map( D => n2801, CK => CLK, Q => n30523, QN 
                           => n_2323);
   clk_r_REG9291_S1 : DFF_X1 port map( D => n2832, CK => CLK, Q => n30522, QN 
                           => n_2324);
   clk_r_REG9227_S1 : DFF_X1 port map( D => n2800, CK => CLK, Q => n30521, QN 
                           => n_2325);
   clk_r_REG9739_S1 : DFF_X1 port map( D => n2736, CK => CLK, Q => n30520, QN 
                           => n_2326);
   clk_r_REG9613_S1 : DFF_X1 port map( D => n2671, CK => CLK, Q => n30519, QN 
                           => n_2327);
   clk_r_REG9551_S1 : DFF_X1 port map( D => n2638, CK => CLK, Q => n30518, QN 
                           => n_2328);
   clk_r_REG9421_S1 : DFF_X1 port map( D => n2575, CK => CLK, Q => n30517, QN 
                           => n_2329);
   clk_r_REG9293_S1 : DFF_X1 port map( D => n2831, CK => CLK, Q => n30516, QN 
                           => n_2330);
   clk_r_REG9229_S1 : DFF_X1 port map( D => n2799, CK => CLK, Q => n30515, QN 
                           => n_2331);
   clk_r_REG9295_S1 : DFF_X1 port map( D => n2830, CK => CLK, Q => n30514, QN 
                           => n_2332);
   clk_r_REG9741_S1 : DFF_X1 port map( D => n2735, CK => CLK, Q => n30513, QN 
                           => n_2333);
   clk_r_REG9231_S1 : DFF_X1 port map( D => n2798, CK => CLK, Q => n30512, QN 
                           => n_2334);
   clk_r_REG9615_S1 : DFF_X1 port map( D => n2670, CK => CLK, Q => n30511, QN 
                           => n_2335);
   clk_r_REG9423_S1 : DFF_X1 port map( D => n2574, CK => CLK, Q => n30510, QN 
                           => n_2336);
   clk_r_REG7602_S1 : DFF_X1 port map( D => n3315, CK => CLK, Q => n30509, QN 
                           => n_2337);
   clk_r_REG7604_S1 : DFF_X1 port map( D => n3314, CK => CLK, Q => n30508, QN 
                           => n_2338);
   clk_r_REG7606_S1 : DFF_X1 port map( D => n3313, CK => CLK, Q => n30507, QN 
                           => n_2339);
   clk_r_REG7608_S1 : DFF_X1 port map( D => n3312, CK => CLK, Q => n30506, QN 
                           => n_2340);
   clk_r_REG7610_S1 : DFF_X1 port map( D => n3311, CK => CLK, Q => n30505, QN 
                           => n_2341);
   clk_r_REG7612_S1 : DFF_X1 port map( D => n3310, CK => CLK, Q => n30504, QN 
                           => n_2342);
   clk_r_REG8627_S1 : DFF_X1 port map( D => n3166, CK => CLK, Q => n30503, QN 
                           => n_2343);
   clk_r_REG8629_S1 : DFF_X1 port map( D => n3165, CK => CLK, Q => n30502, QN 
                           => n_2344);
   clk_r_REG8690_S1 : DFF_X1 port map( D => n2878, CK => CLK, Q => n30501, QN 
                           => n_2345);
   clk_r_REG8435_S1 : DFF_X1 port map( D => n3102, CK => CLK, Q => n30500, QN 
                           => n_2346);
   clk_r_REG7456_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n30499, QN 
                           => n_2347);
   clk_r_REG8437_S1 : DFF_X1 port map( D => n3101, CK => CLK, Q => n30498, QN 
                           => n_2348);
   clk_r_REG9325_S1 : DFF_X1 port map( D => n2558, CK => CLK, Q => n30497, QN 
                           => n_2349);
   clk_r_REG9149_S1 : DFF_X1 port map( D => n3223, CK => CLK, Q => n30496, QN 
                           => n_2350);
   clk_r_REG8289_S1 : DFF_X1 port map( D => n3262, CK => CLK, Q => n30495, QN 
                           => n_2351);
   clk_r_REG7458_S1 : DFF_X1 port map( D => n3293, CK => CLK, Q => n30494, QN 
                           => n_2352);
   clk_r_REG8818_S1 : DFF_X1 port map( D => n2974, CK => CLK, Q => n30493, QN 
                           => n_2353);
   clk_r_REG8994_S1 : DFF_X1 port map( D => n3014, CK => CLK, Q => n30492, QN 
                           => n_2354);
   clk_r_REG9647_S1 : DFF_X1 port map( D => n2718, CK => CLK, Q => n30491, QN 
                           => n_2355);
   clk_r_REG9649_S1 : DFF_X1 port map( D => n2717, CK => CLK, Q => n30490, QN 
                           => n_2356);
   clk_r_REG9088_S1 : DFF_X1 port map( D => n3198, CK => CLK, Q => n30489, QN 
                           => n_2357);
   clk_r_REG9008_S1 : DFF_X1 port map( D => n2782, CK => CLK, Q => n30488, QN 
                           => n_2358);
   clk_r_REG8754_S1 : DFF_X1 port map( D => n2942, CK => CLK, Q => n30487, QN 
                           => n_2359);
   clk_r_REG9151_S1 : DFF_X1 port map( D => n3222, CK => CLK, Q => n30486, QN 
                           => n_2360);
   clk_r_REG8692_S1 : DFF_X1 port map( D => n2877, CK => CLK, Q => n30485, QN 
                           => n_2361);
   clk_r_REG8756_S1 : DFF_X1 port map( D => n2941, CK => CLK, Q => n30484, QN 
                           => n_2362);
   clk_r_REG8820_S1 : DFF_X1 port map( D => n2973, CK => CLK, Q => n30483, QN 
                           => n_2363);
   clk_r_REG8758_S1 : DFF_X1 port map( D => n2940, CK => CLK, Q => n30482, QN 
                           => n_2364);
   clk_r_REG8611_S1 : DFF_X1 port map( D => n3110, CK => CLK, Q => n30481, QN 
                           => n_2365);
   clk_r_REG9010_S1 : DFF_X1 port map( D => n2781, CK => CLK, Q => n30480, QN 
                           => n_2366);
   clk_r_REG8944_S1 : DFF_X1 port map( D => n3039, CK => CLK, Q => n30479, QN 
                           => n_2367);
   clk_r_REG9327_S1 : DFF_X1 port map( D => n2557, CK => CLK, Q => n30478, QN 
                           => n_2368);
   clk_r_REG8439_S1 : DFF_X1 port map( D => n3100, CK => CLK, Q => n30477, QN 
                           => n_2369);
   clk_r_REG9455_S1 : DFF_X1 port map( D => n2622, CK => CLK, Q => n30476, QN 
                           => n_2370);
   clk_r_REG8946_S1 : DFF_X1 port map( D => n3038, CK => CLK, Q => n30475, QN 
                           => n_2371);
   clk_r_REG8694_S1 : DFF_X1 port map( D => n2876, CK => CLK, Q => n30474, QN 
                           => n_2372);
   clk_r_REG8631_S1 : DFF_X1 port map( D => n3164, CK => CLK, Q => n30473, QN 
                           => n_2373);
   clk_r_REG9090_S1 : DFF_X1 port map( D => n3197, CK => CLK, Q => n30472, QN 
                           => n_2374);
   clk_r_REG8561_S1 : DFF_X1 port map( D => n3135, CK => CLK, Q => n30471, QN 
                           => n_2375);
   clk_r_REG8291_S1 : DFF_X1 port map( D => n3261, CK => CLK, Q => n30470, QN 
                           => n_2376);
   clk_r_REG9092_S1 : DFF_X1 port map( D => n3196, CK => CLK, Q => n30469, QN 
                           => n_2377);
   clk_r_REG9651_S1 : DFF_X1 port map( D => n2716, CK => CLK, Q => n30468, QN 
                           => n_2378);
   clk_r_REG7460_S1 : DFF_X1 port map( D => n3292, CK => CLK, Q => n30467, QN 
                           => n_2379);
   clk_r_REG9457_S1 : DFF_X1 port map( D => n2621, CK => CLK, Q => n30466, QN 
                           => n_2380);
   clk_r_REG9459_S1 : DFF_X1 port map( D => n2620, CK => CLK, Q => n30465, QN 
                           => n_2381);
   clk_r_REG8563_S1 : DFF_X1 port map( D => n3134, CK => CLK, Q => n30464, QN 
                           => n_2382);
   clk_r_REG8822_S1 : DFF_X1 port map( D => n2972, CK => CLK, Q => n30463, QN 
                           => n_2383);
   clk_r_REG9153_S1 : DFF_X1 port map( D => n3221, CK => CLK, Q => n30462, QN 
                           => n_2384);
   clk_r_REG8293_S1 : DFF_X1 port map( D => n3260, CK => CLK, Q => n30461, QN 
                           => n_2385);
   clk_r_REG9012_S1 : DFF_X1 port map( D => n2780, CK => CLK, Q => n30460, QN 
                           => n_2386);
   clk_r_REG9329_S1 : DFF_X1 port map( D => n2556, CK => CLK, Q => n30459, QN 
                           => n_2387);
   clk_r_REG9155_S1 : DFF_X1 port map( D => n3220, CK => CLK, Q => n30458, QN 
                           => n_2388);
   clk_r_REG9157_S1 : DFF_X1 port map( D => n3219, CK => CLK, Q => n30457, QN 
                           => n_2389);
   clk_r_REG9159_S1 : DFF_X1 port map( D => n3218, CK => CLK, Q => n30456, QN 
                           => n_2390);
   clk_r_REG9161_S1 : DFF_X1 port map( D => n3217, CK => CLK, Q => n30455, QN 
                           => n_2391);
   clk_r_REG9163_S1 : DFF_X1 port map( D => n3216, CK => CLK, Q => n30454, QN 
                           => n_2392);
   clk_r_REG9165_S1 : DFF_X1 port map( D => n3215, CK => CLK, Q => n30453, QN 
                           => n_2393);
   clk_r_REG8233_S1 : DFF_X1 port map( D => n3483, CK => CLK, Q => n30452, QN 
                           => n_2394);
   clk_r_REG9848_S1 : DFF_X1 port map( D => n3451, CK => CLK, Q => n30451, QN 
                           => n_2395);
   clk_r_REG8373_S1 : DFF_X1 port map( D => n3515, CK => CLK, Q => n30450, QN 
                           => n_2396);
   clk_r_REG7974_S1 : DFF_X1 port map( D => n3387, CK => CLK, Q => n30449, QN 
                           => n_2397);
   clk_r_REG9850_S1 : DFF_X1 port map( D => n3450, CK => CLK, Q => n30448, QN 
                           => n_2398);
   clk_r_REG8235_S1 : DFF_X1 port map( D => n3482, CK => CLK, Q => n30447, QN 
                           => n_2399);
   clk_r_REG7678_S1 : DFF_X1 port map( D => n3355, CK => CLK, Q => n30446, QN 
                           => n_2400);
   clk_r_REG9890_S1 : DFF_X1 port map( D => n3430, CK => CLK, Q => n30445, QN 
                           => n_2401);
   clk_r_REG7680_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n30444, QN 
                           => n_2402);
   clk_r_REG7892_S1 : DFF_X1 port map( D => n3419, CK => CLK, Q => n30443, QN 
                           => n_2403);
   clk_r_REG7894_S1 : DFF_X1 port map( D => n3418, CK => CLK, Q => n30442, QN 
                           => n_2404);
   clk_r_REG8275_S1 : DFF_X1 port map( D => n3462, CK => CLK, Q => n30441, QN 
                           => n_2405);
   clk_r_REG7976_S1 : DFF_X1 port map( D => n3386, CK => CLK, Q => n30440, QN 
                           => n_2406);
   clk_r_REG7934_S1 : DFF_X1 port map( D => n3398, CK => CLK, Q => n30439, QN 
                           => n_2407);
   clk_r_REG8016_S1 : DFF_X1 port map( D => n3366, CK => CLK, Q => n30438, QN 
                           => n_2408);
   clk_r_REG7896_S1 : DFF_X1 port map( D => n3417, CK => CLK, Q => n30437, QN 
                           => n_2409);
   clk_r_REG7720_S1 : DFF_X1 port map( D => n3334, CK => CLK, Q => n30436, QN 
                           => n_2410);
   clk_r_REG7978_S1 : DFF_X1 port map( D => n3385, CK => CLK, Q => n30435, QN 
                           => n_2411);
   clk_r_REG7898_S1 : DFF_X1 port map( D => n3416, CK => CLK, Q => n30434, QN 
                           => n_2412);
   clk_r_REG8375_S1 : DFF_X1 port map( D => n3514, CK => CLK, Q => n30433, QN 
                           => n_2413);
   clk_r_REG9852_S1 : DFF_X1 port map( D => n3449, CK => CLK, Q => n30432, QN 
                           => n_2414);
   clk_r_REG8237_S1 : DFF_X1 port map( D => n3481, CK => CLK, Q => n30431, QN 
                           => n_2415);
   clk_r_REG8415_S1 : DFF_X1 port map( D => n3494, CK => CLK, Q => n30430, QN 
                           => n_2416);
   clk_r_REG8239_S1 : DFF_X1 port map( D => n3480, CK => CLK, Q => n30429, QN 
                           => n_2417);
   clk_r_REG7682_S1 : DFF_X1 port map( D => n3353, CK => CLK, Q => n30428, QN 
                           => n_2418);
   clk_r_REG7684_S1 : DFF_X1 port map( D => n3352, CK => CLK, Q => n30427, QN 
                           => n_2419);
   clk_r_REG8377_S1 : DFF_X1 port map( D => n3513, CK => CLK, Q => n30426, QN 
                           => n_2420);
   clk_r_REG8379_S1 : DFF_X1 port map( D => n3512, CK => CLK, Q => n30425, QN 
                           => n_2421);
   clk_r_REG8241_S1 : DFF_X1 port map( D => n3479, CK => CLK, Q => n30424, QN 
                           => n_2422);
   clk_r_REG9854_S1 : DFF_X1 port map( D => n3448, CK => CLK, Q => n30423, QN 
                           => n_2423);
   clk_r_REG7900_S1 : DFF_X1 port map( D => n3415, CK => CLK, Q => n30422, QN 
                           => n_2424);
   clk_r_REG7980_S1 : DFF_X1 port map( D => n3384, CK => CLK, Q => n30421, QN 
                           => n_2425);
   clk_r_REG7982_S1 : DFF_X1 port map( D => n3383, CK => CLK, Q => n30420, QN 
                           => n_2426);
   clk_r_REG8381_S1 : DFF_X1 port map( D => n3511, CK => CLK, Q => n30419, QN 
                           => n_2427);
   clk_r_REG7686_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n30418, QN 
                           => n_2428);
   clk_r_REG9856_S1 : DFF_X1 port map( D => n3447, CK => CLK, Q => n30417, QN 
                           => n_2429);
   clk_r_REG9937_S1 : DFF_X1 port map( D => n3547, CK => CLK, Q => n30416, QN 
                           => n_2430);
   clk_r_REG9939_S1 : DFF_X1 port map( D => n3546, CK => CLK, Q => n30415, QN 
                           => n_2431);
   clk_r_REG9979_S1 : DFF_X1 port map( D => n3526, CK => CLK, Q => n30414, QN 
                           => n_2432);
   clk_r_REG9941_S1 : DFF_X1 port map( D => n3545, CK => CLK, Q => n30413, QN 
                           => n_2433);
   clk_r_REG9943_S1 : DFF_X1 port map( D => n3544, CK => CLK, Q => n30412, QN 
                           => n_2434);
   clk_r_REG9945_S1 : DFF_X1 port map( D => n3543, CK => CLK, Q => n30411, QN 
                           => n_2435);
   clk_r_REG9947_S1 : DFF_X1 port map( D => n3542, CK => CLK, Q => n30410, QN 
                           => n_2436);
   clk_r_REG9949_S1 : DFF_X1 port map( D => n3541, CK => CLK, Q => n30409, QN 
                           => n_2437);
   clk_r_REG8888_S1 : DFF_X1 port map( D => n3003, CK => CLK, Q => n30408, QN 
                           => n_2438);
   clk_r_REG8890_S1 : DFF_X1 port map( D => n3002, CK => CLK, Q => n30407, QN 
                           => n_2439);
   clk_r_REG8930_S1 : DFF_X1 port map( D => n2982, CK => CLK, Q => n30406, QN 
                           => n_2440);
   clk_r_REG8383_S1 : DFF_X1 port map( D => n3510, CK => CLK, Q => n30405, QN 
                           => n_2441);
   clk_r_REG8892_S1 : DFF_X1 port map( D => n3001, CK => CLK, Q => n30404, QN 
                           => n_2442);
   clk_r_REG8948_S1 : DFF_X1 port map( D => n3037, CK => CLK, Q => n30403, QN 
                           => n_2443);
   clk_r_REG8894_S1 : DFF_X1 port map( D => n3000, CK => CLK, Q => n30402, QN 
                           => n_2444);
   clk_r_REG7902_S1 : DFF_X1 port map( D => n3414, CK => CLK, Q => n30401, QN 
                           => n_2445);
   clk_r_REG8896_S1 : DFF_X1 port map( D => n2999, CK => CLK, Q => n30400, QN 
                           => n_2446);
   clk_r_REG8385_S1 : DFF_X1 port map( D => n3509, CK => CLK, Q => n30399, QN 
                           => n_2447);
   clk_r_REG8898_S1 : DFF_X1 port map( D => n2998, CK => CLK, Q => n30398, QN 
                           => n_2448);
   clk_r_REG7904_S1 : DFF_X1 port map( D => n3413, CK => CLK, Q => n30397, QN 
                           => n_2449);
   clk_r_REG8243_S1 : DFF_X1 port map( D => n3478, CK => CLK, Q => n30396, QN 
                           => n_2450);
   clk_r_REG8245_S1 : DFF_X1 port map( D => n3477, CK => CLK, Q => n30395, QN 
                           => n_2451);
   clk_r_REG8441_S1 : DFF_X1 port map( D => n3099, CK => CLK, Q => n30394, QN 
                           => n_2452);
   clk_r_REG8247_S1 : DFF_X1 port map( D => n3476, CK => CLK, Q => n30393, QN 
                           => n_2453);
   clk_r_REG8387_S1 : DFF_X1 port map( D => n3508, CK => CLK, Q => n30392, QN 
                           => n_2454);
   clk_r_REG8389_S1 : DFF_X1 port map( D => n3507, CK => CLK, Q => n30391, QN 
                           => n_2455);
   clk_r_REG8391_S1 : DFF_X1 port map( D => n3506, CK => CLK, Q => n30390, QN 
                           => n_2456);
   clk_r_REG8393_S1 : DFF_X1 port map( D => n3505, CK => CLK, Q => n30389, QN 
                           => n_2457);
   clk_r_REG7688_S1 : DFF_X1 port map( D => n3350, CK => CLK, Q => n30388, QN 
                           => n_2458);
   clk_r_REG7906_S1 : DFF_X1 port map( D => n3412, CK => CLK, Q => n30387, QN 
                           => n_2459);
   clk_r_REG8395_S1 : DFF_X1 port map( D => n3504, CK => CLK, Q => n30386, QN 
                           => n_2460);
   clk_r_REG9858_S1 : DFF_X1 port map( D => n3446, CK => CLK, Q => n30385, QN 
                           => n_2461);
   clk_r_REG8249_S1 : DFF_X1 port map( D => n3475, CK => CLK, Q => n30384, QN 
                           => n_2462);
   clk_r_REG8251_S1 : DFF_X1 port map( D => n3474, CK => CLK, Q => n30383, QN 
                           => n_2463);
   clk_r_REG8397_S1 : DFF_X1 port map( D => n3503, CK => CLK, Q => n30382, QN 
                           => n_2464);
   clk_r_REG7908_S1 : DFF_X1 port map( D => n3411, CK => CLK, Q => n30381, QN 
                           => n_2465);
   clk_r_REG7910_S1 : DFF_X1 port map( D => n3410, CK => CLK, Q => n30380, QN 
                           => n_2466);
   clk_r_REG9860_S1 : DFF_X1 port map( D => n3445, CK => CLK, Q => n30379, QN 
                           => n_2467);
   clk_r_REG9862_S1 : DFF_X1 port map( D => n3444, CK => CLK, Q => n30378, QN 
                           => n_2468);
   clk_r_REG9864_S1 : DFF_X1 port map( D => n3443, CK => CLK, Q => n30377, QN 
                           => n_2469);
   clk_r_REG9866_S1 : DFF_X1 port map( D => n3442, CK => CLK, Q => n30376, QN 
                           => n_2470);
   clk_r_REG8253_S1 : DFF_X1 port map( D => n3473, CK => CLK, Q => n30375, QN 
                           => n_2471);
   clk_r_REG7912_S1 : DFF_X1 port map( D => n3409, CK => CLK, Q => n30374, QN 
                           => n_2472);
   clk_r_REG8505_S1 : DFF_X1 port map( D => n3067, CK => CLK, Q => n30373, QN 
                           => n_2473);
   clk_r_REG8255_S1 : DFF_X1 port map( D => n3472, CK => CLK, Q => n30372, QN 
                           => n_2474);
   clk_r_REG8257_S1 : DFF_X1 port map( D => n3471, CK => CLK, Q => n30371, QN 
                           => n_2475);
   clk_r_REG7914_S1 : DFF_X1 port map( D => n3408, CK => CLK, Q => n30370, QN 
                           => n_2476);
   clk_r_REG7916_S1 : DFF_X1 port map( D => n3407, CK => CLK, Q => n30369, QN 
                           => n_2477);
   clk_r_REG9868_S1 : DFF_X1 port map( D => n3441, CK => CLK, Q => n30368, QN 
                           => n_2478);
   clk_r_REG7690_S1 : DFF_X1 port map( D => n3349, CK => CLK, Q => n30367, QN 
                           => n_2479);
   clk_r_REG7984_S1 : DFF_X1 port map( D => n3382, CK => CLK, Q => n30366, QN 
                           => n_2480);
   clk_r_REG9870_S1 : DFF_X1 port map( D => n3440, CK => CLK, Q => n30365, QN 
                           => n_2481);
   clk_r_REG9872_S1 : DFF_X1 port map( D => n3439, CK => CLK, Q => n30364, QN 
                           => n_2482);
   clk_r_REG7986_S1 : DFF_X1 port map( D => n3381, CK => CLK, Q => n30363, QN 
                           => n_2483);
   clk_r_REG8507_S1 : DFF_X1 port map( D => n3066, CK => CLK, Q => n30362, QN 
                           => n_2484);
   clk_r_REG8547_S1 : DFF_X1 port map( D => n3046, CK => CLK, Q => n30361, QN 
                           => n_2485);
   clk_r_REG8509_S1 : DFF_X1 port map( D => n3065, CK => CLK, Q => n30360, QN 
                           => n_2486);
   clk_r_REG7692_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n30359, QN 
                           => n_2487);
   clk_r_REG7988_S1 : DFF_X1 port map( D => n3380, CK => CLK, Q => n30358, QN 
                           => n_2488);
   clk_r_REG8511_S1 : DFF_X1 port map( D => n3064, CK => CLK, Q => n30357, QN 
                           => n_2489);
   clk_r_REG8513_S1 : DFF_X1 port map( D => n3063, CK => CLK, Q => n30356, QN 
                           => n_2490);
   clk_r_REG7990_S1 : DFF_X1 port map( D => n3379, CK => CLK, Q => n30355, QN 
                           => n_2491);
   clk_r_REG7694_S1 : DFF_X1 port map( D => n3347, CK => CLK, Q => n30354, QN 
                           => n_2492);
   clk_r_REG7696_S1 : DFF_X1 port map( D => n3346, CK => CLK, Q => n30353, QN 
                           => n_2493);
   clk_r_REG7698_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n30352, QN 
                           => n_2494);
   clk_r_REG8515_S1 : DFF_X1 port map( D => n3062, CK => CLK, Q => n30351, QN 
                           => n_2495);
   clk_r_REG7700_S1 : DFF_X1 port map( D => n3344, CK => CLK, Q => n30350, QN 
                           => n_2496);
   clk_r_REG7702_S1 : DFF_X1 port map( D => n3343, CK => CLK, Q => n30349, QN 
                           => n_2497);
   clk_r_REG7992_S1 : DFF_X1 port map( D => n3378, CK => CLK, Q => n30348, QN 
                           => n_2498);
   clk_r_REG7994_S1 : DFF_X1 port map( D => n3377, CK => CLK, Q => n30347, QN 
                           => n_2499);
   clk_r_REG7996_S1 : DFF_X1 port map( D => n3376, CK => CLK, Q => n30346, QN 
                           => n_2500);
   clk_r_REG7998_S1 : DFF_X1 port map( D => n3375, CK => CLK, Q => n30345, QN 
                           => n_2501);
   clk_r_REG9951_S1 : DFF_X1 port map( D => n3540, CK => CLK, Q => n30344, QN 
                           => n_2502);
   clk_r_REG9953_S1 : DFF_X1 port map( D => n3539, CK => CLK, Q => n30343, QN 
                           => n_2503);
   clk_r_REG9955_S1 : DFF_X1 port map( D => n3538, CK => CLK, Q => n30342, QN 
                           => n_2504);
   clk_r_REG9957_S1 : DFF_X1 port map( D => n3537, CK => CLK, Q => n30341, QN 
                           => n_2505);
   clk_r_REG9959_S1 : DFF_X1 port map( D => n3536, CK => CLK, Q => n30340, QN 
                           => n_2506);
   clk_r_REG9961_S1 : DFF_X1 port map( D => n3535, CK => CLK, Q => n30339, QN 
                           => n_2507);
   clk_r_REG8760_S1 : DFF_X1 port map( D => n2939, CK => CLK, Q => n30338, QN 
                           => n_2508);
   clk_r_REG8762_S1 : DFF_X1 port map( D => n2938, CK => CLK, Q => n30337, QN 
                           => n_2509);
   clk_r_REG8802_S1 : DFF_X1 port map( D => n2918, CK => CLK, Q => n30336, QN 
                           => n_2510);
   clk_r_REG8764_S1 : DFF_X1 port map( D => n2937, CK => CLK, Q => n30335, QN 
                           => n_2511);
   clk_r_REG8766_S1 : DFF_X1 port map( D => n2936, CK => CLK, Q => n30334, QN 
                           => n_2512);
   clk_r_REG8824_S1 : DFF_X1 port map( D => n2971, CK => CLK, Q => n30333, QN 
                           => n_2513);
   clk_r_REG8826_S1 : DFF_X1 port map( D => n2970, CK => CLK, Q => n30332, QN 
                           => n_2514);
   clk_r_REG8866_S1 : DFF_X1 port map( D => n2950, CK => CLK, Q => n30331, QN 
                           => n_2515);
   clk_r_REG8828_S1 : DFF_X1 port map( D => n2969, CK => CLK, Q => n30330, QN 
                           => n_2516);
   clk_r_REG8830_S1 : DFF_X1 port map( D => n2968, CK => CLK, Q => n30329, QN 
                           => n_2517);
   clk_r_REG8832_S1 : DFF_X1 port map( D => n2967, CK => CLK, Q => n30328, QN 
                           => n_2518);
   clk_r_REG8834_S1 : DFF_X1 port map( D => n2966, CK => CLK, Q => n30327, QN 
                           => n_2519);
   clk_r_REG8696_S1 : DFF_X1 port map( D => n2875, CK => CLK, Q => n30326, QN 
                           => n_2520);
   clk_r_REG8698_S1 : DFF_X1 port map( D => n2874, CK => CLK, Q => n30325, QN 
                           => n_2521);
   clk_r_REG8738_S1 : DFF_X1 port map( D => n2854, CK => CLK, Q => n30324, QN 
                           => n_2522);
   clk_r_REG8700_S1 : DFF_X1 port map( D => n2873, CK => CLK, Q => n30323, QN 
                           => n_2523);
   clk_r_REG8702_S1 : DFF_X1 port map( D => n2872, CK => CLK, Q => n30322, QN 
                           => n_2524);
   clk_r_REG8768_S1 : DFF_X1 port map( D => n2935, CK => CLK, Q => n30321, QN 
                           => n_2525);
   clk_r_REG8704_S1 : DFF_X1 port map( D => n2871, CK => CLK, Q => n30320, QN 
                           => n_2526);
   clk_r_REG8706_S1 : DFF_X1 port map( D => n2870, CK => CLK, Q => n30319, QN 
                           => n_2527);
   clk_r_REG8770_S1 : DFF_X1 port map( D => n2934, CK => CLK, Q => n30318, QN 
                           => n_2528);
   clk_r_REG8708_S1 : DFF_X1 port map( D => n2869, CK => CLK, Q => n30317, QN 
                           => n_2529);
   clk_r_REG8950_S1 : DFF_X1 port map( D => n3036, CK => CLK, Q => n30316, QN 
                           => n_2530);
   clk_r_REG9094_S1 : DFF_X1 port map( D => n3195, CK => CLK, Q => n30315, QN 
                           => n_2531);
   clk_r_REG8952_S1 : DFF_X1 port map( D => n3035, CK => CLK, Q => n30314, QN 
                           => n_2532);
   clk_r_REG8954_S1 : DFF_X1 port map( D => n3034, CK => CLK, Q => n30313, QN 
                           => n_2533);
   clk_r_REG8956_S1 : DFF_X1 port map( D => n3033, CK => CLK, Q => n30312, QN 
                           => n_2534);
   clk_r_REG8958_S1 : DFF_X1 port map( D => n3032, CK => CLK, Q => n30311, QN 
                           => n_2535);
   clk_r_REG8960_S1 : DFF_X1 port map( D => n3031, CK => CLK, Q => n30310, QN 
                           => n_2536);
   clk_r_REG8962_S1 : DFF_X1 port map( D => n3030, CK => CLK, Q => n30309, QN 
                           => n_2537);
   clk_r_REG9096_S1 : DFF_X1 port map( D => n3194, CK => CLK, Q => n30308, QN 
                           => n_2538);
   clk_r_REG9098_S1 : DFF_X1 port map( D => n3193, CK => CLK, Q => n30307, QN 
                           => n_2539);
   clk_r_REG8772_S1 : DFF_X1 port map( D => n2933, CK => CLK, Q => n30306, QN 
                           => n_2540);
   clk_r_REG9100_S1 : DFF_X1 port map( D => n3192, CK => CLK, Q => n30305, QN 
                           => n_2541);
   clk_r_REG9102_S1 : DFF_X1 port map( D => n3191, CK => CLK, Q => n30304, QN 
                           => n_2542);
   clk_r_REG9104_S1 : DFF_X1 port map( D => n3190, CK => CLK, Q => n30303, QN 
                           => n_2543);
   clk_r_REG9106_S1 : DFF_X1 port map( D => n3189, CK => CLK, Q => n30302, QN 
                           => n_2544);
   clk_r_REG9108_S1 : DFF_X1 port map( D => n3188, CK => CLK, Q => n30301, QN 
                           => n_2545);
   clk_r_REG9331_S1 : DFF_X1 port map( D => n2555, CK => CLK, Q => n30300, QN 
                           => n_2546);
   clk_r_REG8900_S1 : DFF_X1 port map( D => n2997, CK => CLK, Q => n30299, QN 
                           => n_2547);
   clk_r_REG8633_S1 : DFF_X1 port map( D => n3163, CK => CLK, Q => n30298, QN 
                           => n_2548);
   clk_r_REG8635_S1 : DFF_X1 port map( D => n3162, CK => CLK, Q => n30297, QN 
                           => n_2549);
   clk_r_REG8637_S1 : DFF_X1 port map( D => n3161, CK => CLK, Q => n30296, QN 
                           => n_2550);
   clk_r_REG8639_S1 : DFF_X1 port map( D => n3160, CK => CLK, Q => n30295, QN 
                           => n_2551);
   clk_r_REG8641_S1 : DFF_X1 port map( D => n3159, CK => CLK, Q => n30294, QN 
                           => n_2552);
   clk_r_REG8643_S1 : DFF_X1 port map( D => n3158, CK => CLK, Q => n30293, QN 
                           => n_2553);
   clk_r_REG9333_S1 : DFF_X1 port map( D => n2554, CK => CLK, Q => n30292, QN 
                           => n_2554);
   clk_r_REG8836_S1 : DFF_X1 port map( D => n2965, CK => CLK, Q => n30291, QN 
                           => n_2555);
   clk_r_REG8645_S1 : DFF_X1 port map( D => n3157, CK => CLK, Q => n30290, QN 
                           => n_2556);
   clk_r_REG8647_S1 : DFF_X1 port map( D => n3156, CK => CLK, Q => n30289, QN 
                           => n_2557);
   clk_r_REG8565_S1 : DFF_X1 port map( D => n3133, CK => CLK, Q => n30288, QN 
                           => n_2558);
   clk_r_REG8567_S1 : DFF_X1 port map( D => n3132, CK => CLK, Q => n30287, QN 
                           => n_2559);
   clk_r_REG8569_S1 : DFF_X1 port map( D => n3131, CK => CLK, Q => n30286, QN 
                           => n_2560);
   clk_r_REG8571_S1 : DFF_X1 port map( D => n3130, CK => CLK, Q => n30285, QN 
                           => n_2561);
   clk_r_REG8573_S1 : DFF_X1 port map( D => n3129, CK => CLK, Q => n30284, QN 
                           => n_2562);
   clk_r_REG9461_S1 : DFF_X1 port map( D => n2619, CK => CLK, Q => n30283, QN 
                           => n_2563);
   clk_r_REG9653_S1 : DFF_X1 port map( D => n2715, CK => CLK, Q => n30282, QN 
                           => n_2564);
   clk_r_REG9373_S1 : DFF_X1 port map( D => n2534, CK => CLK, Q => n30281, QN 
                           => n_2565);
   clk_r_REG8575_S1 : DFF_X1 port map( D => n3128, CK => CLK, Q => n30280, QN 
                           => n_2566);
   clk_r_REG8577_S1 : DFF_X1 port map( D => n3127, CK => CLK, Q => n30279, QN 
                           => n_2567);
   clk_r_REG8579_S1 : DFF_X1 port map( D => n3126, CK => CLK, Q => n30278, QN 
                           => n_2568);
   clk_r_REG9335_S1 : DFF_X1 port map( D => n2553, CK => CLK, Q => n30277, QN 
                           => n_2569);
   clk_r_REG9655_S1 : DFF_X1 port map( D => n2714, CK => CLK, Q => n30276, QN 
                           => n_2570);
   clk_r_REG9695_S1 : DFF_X1 port map( D => n2694, CK => CLK, Q => n30275, QN 
                           => n_2571);
   clk_r_REG9657_S1 : DFF_X1 port map( D => n2713, CK => CLK, Q => n30274, QN 
                           => n_2572);
   clk_r_REG9659_S1 : DFF_X1 port map( D => n2712, CK => CLK, Q => n30273, QN 
                           => n_2573);
   clk_r_REG9337_S1 : DFF_X1 port map( D => n2552, CK => CLK, Q => n30272, QN 
                           => n_2574);
   clk_r_REG8443_S1 : DFF_X1 port map( D => n3098, CK => CLK, Q => n30271, QN 
                           => n_2575);
   clk_r_REG8483_S1 : DFF_X1 port map( D => n3078, CK => CLK, Q => n30270, QN 
                           => n_2576);
   clk_r_REG8445_S1 : DFF_X1 port map( D => n3097, CK => CLK, Q => n30269, QN 
                           => n_2577);
   clk_r_REG8517_S1 : DFF_X1 port map( D => n3061, CK => CLK, Q => n30268, QN 
                           => n_2578);
   clk_r_REG8447_S1 : DFF_X1 port map( D => n3096, CK => CLK, Q => n30267, QN 
                           => n_2579);
   clk_r_REG8449_S1 : DFF_X1 port map( D => n3095, CK => CLK, Q => n30266, QN 
                           => n_2580);
   clk_r_REG8451_S1 : DFF_X1 port map( D => n3094, CK => CLK, Q => n30265, QN 
                           => n_2581);
   clk_r_REG8453_S1 : DFF_X1 port map( D => n3093, CK => CLK, Q => n30264, QN 
                           => n_2582);
   clk_r_REG9661_S1 : DFF_X1 port map( D => n2711, CK => CLK, Q => n30263, QN 
                           => n_2583);
   clk_r_REG9663_S1 : DFF_X1 port map( D => n2710, CK => CLK, Q => n30262, QN 
                           => n_2584);
   clk_r_REG9463_S1 : DFF_X1 port map( D => n2618, CK => CLK, Q => n30261, QN 
                           => n_2585);
   clk_r_REG9481_S1 : DFF_X1 port map( D => n2606, CK => CLK, Q => n30260, QN 
                           => n_2586);
   clk_r_REG9483_S1 : DFF_X1 port map( D => n2617, CK => CLK, Q => n30259, QN 
                           => n_2587);
   clk_r_REG9339_S1 : DFF_X1 port map( D => n2551, CK => CLK, Q => n30258, QN 
                           => n_2588);
   clk_r_REG9485_S1 : DFF_X1 port map( D => n2616, CK => CLK, Q => n30257, QN 
                           => n_2589);
   clk_r_REG9487_S1 : DFF_X1 port map( D => n2615, CK => CLK, Q => n30256, QN 
                           => n_2590);
   clk_r_REG9489_S1 : DFF_X1 port map( D => n2614, CK => CLK, Q => n30255, QN 
                           => n_2591);
   clk_r_REG7462_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n30254, QN 
                           => n_2592);
   clk_r_REG7464_S1 : DFF_X1 port map( D => n3290, CK => CLK, Q => n30253, QN 
                           => n_2593);
   clk_r_REG7504_S1 : DFF_X1 port map( D => n3270, CK => CLK, Q => n30252, QN 
                           => n_2594);
   clk_r_REG7466_S1 : DFF_X1 port map( D => n3289, CK => CLK, Q => n30251, QN 
                           => n_2595);
   clk_r_REG7468_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n30250, QN 
                           => n_2596);
   clk_r_REG7470_S1 : DFF_X1 port map( D => n3287, CK => CLK, Q => n30249, QN 
                           => n_2597);
   clk_r_REG7472_S1 : DFF_X1 port map( D => n3286, CK => CLK, Q => n30248, QN 
                           => n_2598);
   clk_r_REG7474_S1 : DFF_X1 port map( D => n3285, CK => CLK, Q => n30247, QN 
                           => n_2599);
   clk_r_REG9014_S1 : DFF_X1 port map( D => n2779, CK => CLK, Q => n30246, QN 
                           => n_2600);
   clk_r_REG9016_S1 : DFF_X1 port map( D => n2778, CK => CLK, Q => n30245, QN 
                           => n_2601);
   clk_r_REG9056_S1 : DFF_X1 port map( D => n2758, CK => CLK, Q => n30244, QN 
                           => n_2602);
   clk_r_REG9018_S1 : DFF_X1 port map( D => n2777, CK => CLK, Q => n30243, QN 
                           => n_2603);
   clk_r_REG9020_S1 : DFF_X1 port map( D => n2776, CK => CLK, Q => n30242, QN 
                           => n_2604);
   clk_r_REG9022_S1 : DFF_X1 port map( D => n2775, CK => CLK, Q => n30241, QN 
                           => n_2605);
   clk_r_REG9024_S1 : DFF_X1 port map( D => n2774, CK => CLK, Q => n30240, QN 
                           => n_2606);
   clk_r_REG8295_S1 : DFF_X1 port map( D => n3259, CK => CLK, Q => n30239, QN 
                           => n_2607);
   clk_r_REG8297_S1 : DFF_X1 port map( D => n3258, CK => CLK, Q => n30238, QN 
                           => n_2608);
   clk_r_REG8299_S1 : DFF_X1 port map( D => n3257, CK => CLK, Q => n30237, QN 
                           => n_2609);
   clk_r_REG8301_S1 : DFF_X1 port map( D => n3256, CK => CLK, Q => n30236, QN 
                           => n_2610);
   clk_r_REG8303_S1 : DFF_X1 port map( D => n3255, CK => CLK, Q => n30235, QN 
                           => n_2611);
   clk_r_REG8305_S1 : DFF_X1 port map( D => n3254, CK => CLK, Q => n30234, QN 
                           => n_2612);
   clk_r_REG8307_S1 : DFF_X1 port map( D => n3253, CK => CLK, Q => n30233, QN 
                           => n_2613);
   clk_r_REG8309_S1 : DFF_X1 port map( D => n3252, CK => CLK, Q => n30232, QN 
                           => n_2614);
   clk_r_REG8581_S1 : DFF_X1 port map( D => n3125, CK => CLK, Q => n30231, QN 
                           => n_2615);
   clk_r_REG8455_S1 : DFF_X1 port map( D => n3092, CK => CLK, Q => n30230, QN 
                           => n_2616);
   clk_r_REG9110_S1 : DFF_X1 port map( D => n3187, CK => CLK, Q => n30229, QN 
                           => n_2617);
   clk_r_REG9491_S1 : DFF_X1 port map( D => n2613, CK => CLK, Q => n30228, QN 
                           => n_2618);
   clk_r_REG9665_S1 : DFF_X1 port map( D => n2709, CK => CLK, Q => n30227, QN 
                           => n_2619);
   clk_r_REG8710_S1 : DFF_X1 port map( D => n2868, CK => CLK, Q => n30226, QN 
                           => n_2620);
   clk_r_REG8649_S1 : DFF_X1 port map( D => n3155, CK => CLK, Q => n30225, QN 
                           => n_2621);
   clk_r_REG7476_S1 : DFF_X1 port map( D => n3284, CK => CLK, Q => n30224, QN 
                           => n_2622);
   clk_r_REG8964_S1 : DFF_X1 port map( D => n3029, CK => CLK, Q => n30223, QN 
                           => n_2623);
   clk_r_REG8311_S1 : DFF_X1 port map( D => n3251, CK => CLK, Q => n30222, QN 
                           => n_2624);
   clk_r_REG9112_S1 : DFF_X1 port map( D => n3186, CK => CLK, Q => n30221, QN 
                           => n_2625);
   clk_r_REG9026_S1 : DFF_X1 port map( D => n2773, CK => CLK, Q => n30220, QN 
                           => n_2626);
   clk_r_REG8774_S1 : DFF_X1 port map( D => n2932, CK => CLK, Q => n30219, QN 
                           => n_2627);
   clk_r_REG8519_S1 : DFF_X1 port map( D => n3060, CK => CLK, Q => n30218, QN 
                           => n_2628);
   clk_r_REG8651_S1 : DFF_X1 port map( D => n3154, CK => CLK, Q => n30217, QN 
                           => n_2629);
   clk_r_REG8838_S1 : DFF_X1 port map( D => n2964, CK => CLK, Q => n30216, QN 
                           => n_2630);
   clk_r_REG9493_S1 : DFF_X1 port map( D => n2612, CK => CLK, Q => n30215, QN 
                           => n_2631);
   clk_r_REG8583_S1 : DFF_X1 port map( D => n3124, CK => CLK, Q => n30214, QN 
                           => n_2632);
   clk_r_REG8653_S1 : DFF_X1 port map( D => n3153, CK => CLK, Q => n30213, QN 
                           => n_2633);
   clk_r_REG9028_S1 : DFF_X1 port map( D => n2772, CK => CLK, Q => n30212, QN 
                           => n_2634);
   clk_r_REG8585_S1 : DFF_X1 port map( D => n3123, CK => CLK, Q => n30211, QN 
                           => n_2635);
   clk_r_REG8313_S1 : DFF_X1 port map( D => n3250, CK => CLK, Q => n30210, QN 
                           => n_2636);
   clk_r_REG8457_S1 : DFF_X1 port map( D => n3091, CK => CLK, Q => n30209, QN 
                           => n_2637);
   clk_r_REG9667_S1 : DFF_X1 port map( D => n2708, CK => CLK, Q => n30208, QN 
                           => n_2638);
   clk_r_REG8521_S1 : DFF_X1 port map( D => n3059, CK => CLK, Q => n30207, QN 
                           => n_2639);
   clk_r_REG8712_S1 : DFF_X1 port map( D => n2867, CK => CLK, Q => n30206, QN 
                           => n_2640);
   clk_r_REG8966_S1 : DFF_X1 port map( D => n3028, CK => CLK, Q => n30205, QN 
                           => n_2641);
   clk_r_REG7478_S1 : DFF_X1 port map( D => n3283, CK => CLK, Q => n30204, QN 
                           => n_2642);
   clk_r_REG8902_S1 : DFF_X1 port map( D => n2996, CK => CLK, Q => n30203, QN 
                           => n_2643);
   clk_r_REG8315_S1 : DFF_X1 port map( D => n3249, CK => CLK, Q => n30202, QN 
                           => n_2644);
   clk_r_REG9114_S1 : DFF_X1 port map( D => n3185, CK => CLK, Q => n30201, QN 
                           => n_2645);
   clk_r_REG8776_S1 : DFF_X1 port map( D => n2931, CK => CLK, Q => n30200, QN 
                           => n_2646);
   clk_r_REG7480_S1 : DFF_X1 port map( D => n3282, CK => CLK, Q => n30199, QN 
                           => n_2647);
   clk_r_REG8840_S1 : DFF_X1 port map( D => n2963, CK => CLK, Q => n30198, QN 
                           => n_2648);
   clk_r_REG8968_S1 : DFF_X1 port map( D => n3027, CK => CLK, Q => n30197, QN 
                           => n_2649);
   clk_r_REG8904_S1 : DFF_X1 port map( D => n2995, CK => CLK, Q => n30196, QN 
                           => n_2650);
   clk_r_REG8970_S1 : DFF_X1 port map( D => n3026, CK => CLK, Q => n30195, QN 
                           => n_2651);
   clk_r_REG8523_S1 : DFF_X1 port map( D => n3058, CK => CLK, Q => n30194, QN 
                           => n_2652);
   clk_r_REG8842_S1 : DFF_X1 port map( D => n2962, CK => CLK, Q => n30193, QN 
                           => n_2653);
   clk_r_REG8778_S1 : DFF_X1 port map( D => n2930, CK => CLK, Q => n30192, QN 
                           => n_2654);
   clk_r_REG8714_S1 : DFF_X1 port map( D => n2866, CK => CLK, Q => n30191, QN 
                           => n_2655);
   clk_r_REG9030_S1 : DFF_X1 port map( D => n2771, CK => CLK, Q => n30190, QN 
                           => n_2656);
   clk_r_REG9669_S1 : DFF_X1 port map( D => n2707, CK => CLK, Q => n30189, QN 
                           => n_2657);
   clk_r_REG9495_S1 : DFF_X1 port map( D => n2611, CK => CLK, Q => n30188, QN 
                           => n_2658);
   clk_r_REG7482_S1 : DFF_X1 port map( D => n3281, CK => CLK, Q => n30187, QN 
                           => n_2659);
   clk_r_REG8459_S1 : DFF_X1 port map( D => n3090, CK => CLK, Q => n30186, QN 
                           => n_2660);
   clk_r_REG8587_S1 : DFF_X1 port map( D => n3122, CK => CLK, Q => n30185, QN 
                           => n_2661);
   clk_r_REG8716_S1 : DFF_X1 port map( D => n2865, CK => CLK, Q => n30184, QN 
                           => n_2662);
   clk_r_REG8655_S1 : DFF_X1 port map( D => n3152, CK => CLK, Q => n30183, QN 
                           => n_2663);
   clk_r_REG9116_S1 : DFF_X1 port map( D => n3184, CK => CLK, Q => n30182, QN 
                           => n_2664);
   clk_r_REG8780_S1 : DFF_X1 port map( D => n2929, CK => CLK, Q => n30181, QN 
                           => n_2665);
   clk_r_REG8317_S1 : DFF_X1 port map( D => n3248, CK => CLK, Q => n30180, QN 
                           => n_2666);
   clk_r_REG7484_S1 : DFF_X1 port map( D => n3280, CK => CLK, Q => n30179, QN 
                           => n_2667);
   clk_r_REG8319_S1 : DFF_X1 port map( D => n3247, CK => CLK, Q => n30178, QN 
                           => n_2668);
   clk_r_REG8844_S1 : DFF_X1 port map( D => n2961, CK => CLK, Q => n30177, QN 
                           => n_2669);
   clk_r_REG9118_S1 : DFF_X1 port map( D => n3183, CK => CLK, Q => n30176, QN 
                           => n_2670);
   clk_r_REG8657_S1 : DFF_X1 port map( D => n3151, CK => CLK, Q => n30175, QN 
                           => n_2671);
   clk_r_REG8589_S1 : DFF_X1 port map( D => n3121, CK => CLK, Q => n30174, QN 
                           => n_2672);
   clk_r_REG8718_S1 : DFF_X1 port map( D => n2864, CK => CLK, Q => n30173, QN 
                           => n_2673);
   clk_r_REG8461_S1 : DFF_X1 port map( D => n3089, CK => CLK, Q => n30172, QN 
                           => n_2674);
   clk_r_REG8906_S1 : DFF_X1 port map( D => n2994, CK => CLK, Q => n30171, QN 
                           => n_2675);
   clk_r_REG8525_S1 : DFF_X1 port map( D => n3057, CK => CLK, Q => n30170, QN 
                           => n_2676);
   clk_r_REG8782_S1 : DFF_X1 port map( D => n2928, CK => CLK, Q => n30169, QN 
                           => n_2677);
   clk_r_REG8846_S1 : DFF_X1 port map( D => n2960, CK => CLK, Q => n30168, QN 
                           => n_2678);
   clk_r_REG8908_S1 : DFF_X1 port map( D => n2993, CK => CLK, Q => n30167, QN 
                           => n_2679);
   clk_r_REG8972_S1 : DFF_X1 port map( D => n3025, CK => CLK, Q => n30166, QN 
                           => n_2680);
   clk_r_REG8527_S1 : DFF_X1 port map( D => n3056, CK => CLK, Q => n30165, QN 
                           => n_2681);
   clk_r_REG8910_S1 : DFF_X1 port map( D => n2992, CK => CLK, Q => n30164, QN 
                           => n_2682);
   clk_r_REG9497_S1 : DFF_X1 port map( D => n2610, CK => CLK, Q => n30163, QN 
                           => n_2683);
   clk_r_REG8463_S1 : DFF_X1 port map( D => n3088, CK => CLK, Q => n30162, QN 
                           => n_2684);
   clk_r_REG8591_S1 : DFF_X1 port map( D => n3120, CK => CLK, Q => n30161, QN 
                           => n_2685);
   clk_r_REG8659_S1 : DFF_X1 port map( D => n3150, CK => CLK, Q => n30160, QN 
                           => n_2686);
   clk_r_REG9120_S1 : DFF_X1 port map( D => n3182, CK => CLK, Q => n30159, QN 
                           => n_2687);
   clk_r_REG8321_S1 : DFF_X1 port map( D => n3246, CK => CLK, Q => n30158, QN 
                           => n_2688);
   clk_r_REG7486_S1 : DFF_X1 port map( D => n3279, CK => CLK, Q => n30157, QN 
                           => n_2689);
   clk_r_REG9671_S1 : DFF_X1 port map( D => n2706, CK => CLK, Q => n30156, QN 
                           => n_2690);
   clk_r_REG9032_S1 : DFF_X1 port map( D => n2770, CK => CLK, Q => n30155, QN 
                           => n_2691);
   clk_r_REG8720_S1 : DFF_X1 port map( D => n2863, CK => CLK, Q => n30154, QN 
                           => n_2692);
   clk_r_REG8465_S1 : DFF_X1 port map( D => n3087, CK => CLK, Q => n30153, QN 
                           => n_2693);
   clk_r_REG8784_S1 : DFF_X1 port map( D => n2927, CK => CLK, Q => n30152, QN 
                           => n_2694);
   clk_r_REG9499_S1 : DFF_X1 port map( D => n2609, CK => CLK, Q => n30151, QN 
                           => n_2695);
   clk_r_REG9673_S1 : DFF_X1 port map( D => n2705, CK => CLK, Q => n30150, QN 
                           => n_2696);
   clk_r_REG8848_S1 : DFF_X1 port map( D => n2959, CK => CLK, Q => n30149, QN 
                           => n_2697);
   clk_r_REG9034_S1 : DFF_X1 port map( D => n2769, CK => CLK, Q => n30148, QN 
                           => n_2698);
   clk_r_REG8912_S1 : DFF_X1 port map( D => n2991, CK => CLK, Q => n30147, QN 
                           => n_2699);
   clk_r_REG8529_S1 : DFF_X1 port map( D => n3055, CK => CLK, Q => n30146, QN 
                           => n_2700);
   clk_r_REG9341_S1 : DFF_X1 port map( D => n2550, CK => CLK, Q => n30145, QN 
                           => n_2701);
   clk_r_REG9675_S1 : DFF_X1 port map( D => n2704, CK => CLK, Q => n30144, QN 
                           => n_2702);
   clk_r_REG9036_S1 : DFF_X1 port map( D => n2768, CK => CLK, Q => n30143, QN 
                           => n_2703);
   clk_r_REG9343_S1 : DFF_X1 port map( D => n2549, CK => CLK, Q => n30142, QN 
                           => n_2704);
   clk_r_REG9345_S1 : DFF_X1 port map( D => n2548, CK => CLK, Q => n30141, QN 
                           => n_2705);
   clk_r_REG9347_S1 : DFF_X1 port map( D => n2547, CK => CLK, Q => n30140, QN 
                           => n_2706);
   clk_r_REG9349_S1 : DFF_X1 port map( D => n2546, CK => CLK, Q => n30139, QN 
                           => n_2707);
   clk_r_REG9501_S1 : DFF_X1 port map( D => n2608, CK => CLK, Q => n30138, QN 
                           => n_2708);
   clk_r_REG9503_S1 : DFF_X1 port map( D => n2607, CK => CLK, Q => n30137, QN 
                           => n_2709);
   clk_r_REG9677_S1 : DFF_X1 port map( D => n2703, CK => CLK, Q => n30136, QN 
                           => n_2710);
   clk_r_REG9351_S1 : DFF_X1 port map( D => n2545, CK => CLK, Q => n30135, QN 
                           => n_2711);
   clk_r_REG9353_S1 : DFF_X1 port map( D => n2544, CK => CLK, Q => n30134, QN 
                           => n_2712);
   clk_r_REG9355_S1 : DFF_X1 port map( D => n2543, CK => CLK, Q => n30133, QN 
                           => n_2713);
   clk_r_REG10248_S7 : DFFS_X1 port map( D => n3569, CK => CLK, SN => RESET_BAR
                           , Q => n30132, QN => n_2714);
   clk_r_REG10290_S7 : DFFS_X1 port map( D => n3560, CK => CLK, SN => RESET_BAR
                           , Q => n30131, QN => n_2715);
   clk_r_REG10061_S4 : DFFR_X1 port map( D => n35760, CK => CLK, RN => 
                           RESET_BAR, Q => n30130, QN => n_2716);
   clk_r_REG10057_S4 : DFFR_X1 port map( D => n35759, CK => CLK, RN => 
                           RESET_BAR, Q => n30129, QN => n_2717);
   clk_r_REG10034_S3 : DFFR_X1 port map( D => n18358, CK => CLK, RN => 
                           RESET_BAR, Q => n30122, QN => n_2718);
   clk_r_REG10035_S4 : DFFR_X1 port map( D => n30122, CK => CLK, RN => 
                           RESET_BAR, Q => n30121, QN => n_2719);
   clk_r_REG10032_S3 : DFFR_X1 port map( D => n18356, CK => CLK, RN => 
                           RESET_BAR, Q => n30119, QN => n_2720);
   clk_r_REG10033_S4 : DFFR_X1 port map( D => n30119, CK => CLK, RN => 
                           RESET_BAR, Q => n30118, QN => n_2721);
   clk_r_REG10026_S3 : DFFR_X1 port map( D => n18352, CK => CLK, RN => 
                           RESET_BAR, Q => n30114, QN => n_2722);
   clk_r_REG10027_S4 : DFFR_X1 port map( D => n30114, CK => CLK, RN => 
                           RESET_BAR, Q => n30113, QN => n_2723);
   clk_r_REG10024_S3 : DFFR_X1 port map( D => n18350, CK => CLK, RN => 
                           RESET_BAR, Q => n30111, QN => n_2724);
   clk_r_REG10025_S4 : DFFR_X1 port map( D => n30111, CK => CLK, RN => 
                           RESET_BAR, Q => n30110, QN => n_2725);
   clk_r_REG10231_S7 : DFFR_X1 port map( D => n18324, CK => CLK, RN => 
                           RESET_BAR, Q => n30084, QN => n_2726);
   clk_r_REG10224_S7 : DFFR_X1 port map( D => n18323, CK => CLK, RN => 
                           RESET_BAR, Q => n30083, QN => n_2727);
   clk_r_REG10218_S7 : DFFR_X1 port map( D => n18322, CK => CLK, RN => 
                           RESET_BAR, Q => n30082, QN => n_2728);
   clk_r_REG10210_S7 : DFFR_X1 port map( D => n18321, CK => CLK, RN => 
                           RESET_BAR, Q => n30081, QN => n_2729);
   clk_r_REG10216_S7 : DFFR_X1 port map( D => n18320, CK => CLK, RN => 
                           RESET_BAR, Q => n30080, QN => n_2730);
   clk_r_REG10203_S7 : DFFR_X1 port map( D => n18319, CK => CLK, RN => 
                           RESET_BAR, Q => n30079, QN => n_2731);
   clk_r_REG10196_S7 : DFFR_X1 port map( D => n18318, CK => CLK, RN => 
                           RESET_BAR, Q => n30078, QN => n_2732);
   clk_r_REG10208_S7 : DFFR_X1 port map( D => n18317, CK => CLK, RN => 
                           RESET_BAR, Q => n30077, QN => n_2733);
   clk_r_REG10238_S7 : DFFR_X1 port map( D => n18316, CK => CLK, RN => 
                           RESET_BAR, Q => n30076, QN => n_2734);
   clk_r_REG10229_S7 : DFFR_X1 port map( D => n18315, CK => CLK, RN => 
                           RESET_BAR, Q => n30075, QN => n_2735);
   clk_r_REG10236_S7 : DFFR_X1 port map( D => n18314, CK => CLK, RN => 
                           RESET_BAR, Q => n30074, QN => n_2736);
   clk_r_REG10189_S7 : DFFR_X1 port map( D => n18313, CK => CLK, RN => 
                           RESET_BAR, Q => n30073, QN => n_2737);
   clk_r_REG10187_S7 : DFFR_X1 port map( D => n18312, CK => CLK, RN => 
                           RESET_BAR, Q => n30072, QN => n_2738);
   clk_r_REG10201_S7 : DFFR_X1 port map( D => n18311, CK => CLK, RN => 
                           RESET_BAR, Q => n30071, QN => n_2739);
   clk_r_REG10222_S7 : DFFR_X1 port map( D => n18310, CK => CLK, RN => 
                           RESET_BAR, Q => n30070, QN => n_2740);
   clk_r_REG10194_S7 : DFFR_X1 port map( D => n18309, CK => CLK, RN => 
                           RESET_BAR, Q => n30069, QN => n_2741);
   clk_r_REG10147_S7 : DFFR_X1 port map( D => n18308, CK => CLK, RN => 
                           RESET_BAR, Q => n30068, QN => n_2742);
   clk_r_REG10132_S7 : DFFR_X1 port map( D => n18307, CK => CLK, RN => 
                           RESET_BAR, Q => n30067, QN => n_2743);
   clk_r_REG10145_S7 : DFFR_X1 port map( D => n18306, CK => CLK, RN => 
                           RESET_BAR, Q => n30066, QN => n_2744);
   clk_r_REG10161_S7 : DFFR_X1 port map( D => n18305, CK => CLK, RN => 
                           RESET_BAR, Q => n30065, QN => n_2745);
   clk_r_REG10168_S7 : DFFR_X1 port map( D => n18304, CK => CLK, RN => 
                           RESET_BAR, Q => n30064, QN => n_2746);
   clk_r_REG10175_S7 : DFFR_X1 port map( D => n18303, CK => CLK, RN => 
                           RESET_BAR, Q => n30063, QN => n_2747);
   clk_r_REG10154_S7 : DFFR_X1 port map( D => n18302, CK => CLK, RN => 
                           RESET_BAR, Q => n30062, QN => n_2748);
   clk_r_REG10159_S7 : DFFR_X1 port map( D => n18301, CK => CLK, RN => 
                           RESET_BAR, Q => n30061, QN => n_2749);
   clk_r_REG10130_S7 : DFFR_X1 port map( D => n18300, CK => CLK, RN => 
                           RESET_BAR, Q => n30060, QN => n_2750);
   clk_r_REG10173_S7 : DFFR_X1 port map( D => n18299, CK => CLK, RN => 
                           RESET_BAR, Q => n30059, QN => n_2751);
   clk_r_REG10181_S7 : DFFR_X1 port map( D => n18298, CK => CLK, RN => 
                           RESET_BAR, Q => n30058, QN => n_2752);
   clk_r_REG10179_S7 : DFFR_X1 port map( D => n18297, CK => CLK, RN => 
                           RESET_BAR, Q => n30057, QN => n_2753);
   clk_r_REG10140_S7 : DFFR_X1 port map( D => n18296, CK => CLK, RN => 
                           RESET_BAR, Q => n30056, QN => n_2754);
   clk_r_REG10152_S7 : DFFR_X1 port map( D => n18295, CK => CLK, RN => 
                           RESET_BAR, Q => n30055, QN => n_2755);
   clk_r_REG10166_S7 : DFFR_X1 port map( D => n18294, CK => CLK, RN => 
                           RESET_BAR, Q => n30054, QN => n_2756);
   clk_r_REG10138_S7 : DFFR_X1 port map( D => n18293, CK => CLK, RN => 
                           RESET_BAR, Q => n30053, QN => n_2757);
   clk_r_REG10038_S3 : DFFS_X1 port map( D => n18284, CK => CLK, SN => 
                           RESET_BAR, Q => n30049, QN => n_2758);
   clk_r_REG10039_S4 : DFFS_X1 port map( D => n30049, CK => CLK, SN => 
                           RESET_BAR, Q => n30048, QN => n_2759);
   clk_r_REG10036_S3 : DFFR_X1 port map( D => n18283, CK => CLK, RN => 
                           RESET_BAR, Q => n30047, QN => n_2760);
   clk_r_REG10037_S4 : DFFR_X1 port map( D => n30047, CK => CLK, RN => 
                           RESET_BAR, Q => n30046, QN => n_2761);
   clk_r_REG10030_S3 : DFFR_X1 port map( D => n18282, CK => CLK, RN => 
                           RESET_BAR, Q => n30045, QN => n_2762);
   clk_r_REG10031_S4 : DFFR_X1 port map( D => n30045, CK => CLK, RN => 
                           RESET_BAR, Q => n30044, QN => n_2763);
   clk_r_REG10028_S3 : DFFR_X1 port map( D => n18281, CK => CLK, RN => 
                           RESET_BAR, Q => n30043, QN => n_2764);
   clk_r_REG10029_S4 : DFFR_X1 port map( D => n30043, CK => CLK, RN => 
                           RESET_BAR, Q => n30042, QN => n_2765);
   clk_r_REG9354_S1 : DFF_X1 port map( D => n2543, CK => CLK, Q => n_2766, QN 
                           => n30041);
   clk_r_REG9352_S1 : DFF_X1 port map( D => n2544, CK => CLK, Q => n_2767, QN 
                           => n30040);
   clk_r_REG9350_S1 : DFF_X1 port map( D => n2545, CK => CLK, Q => n_2768, QN 
                           => n30039);
   clk_r_REG9037_S1 : DFF_X1 port map( D => n2767, CK => CLK, Q => n_2769, QN 
                           => n30038);
   clk_r_REG9676_S1 : DFF_X1 port map( D => n2703, CK => CLK, Q => n_2770, QN 
                           => n30037);
   clk_r_REG9502_S1 : DFF_X1 port map( D => n2607, CK => CLK, Q => n_2771, QN 
                           => n30036);
   clk_r_REG9500_S1 : DFF_X1 port map( D => n2608, CK => CLK, Q => n_2772, QN 
                           => n30035);
   clk_r_REG9348_S1 : DFF_X1 port map( D => n2546, CK => CLK, Q => n_2773, QN 
                           => n30034);
   clk_r_REG9346_S1 : DFF_X1 port map( D => n2547, CK => CLK, Q => n_2774, QN 
                           => n30033);
   clk_r_REG9344_S1 : DFF_X1 port map( D => n2548, CK => CLK, Q => n_2775, QN 
                           => n30032);
   clk_r_REG9342_S1 : DFF_X1 port map( D => n2549, CK => CLK, Q => n_2776, QN 
                           => n30031);
   clk_r_REG9035_S1 : DFF_X1 port map( D => n2768, CK => CLK, Q => n_2777, QN 
                           => n30030);
   clk_r_REG9674_S1 : DFF_X1 port map( D => n2704, CK => CLK, Q => n_2778, QN 
                           => n30029);
   clk_r_REG9340_S1 : DFF_X1 port map( D => n2550, CK => CLK, Q => n_2779, QN 
                           => n30028);
   clk_r_REG8528_S1 : DFF_X1 port map( D => n3055, CK => CLK, Q => n_2780, QN 
                           => n30027);
   clk_r_REG8911_S1 : DFF_X1 port map( D => n2991, CK => CLK, Q => n_2781, QN 
                           => n30026);
   clk_r_REG9033_S1 : DFF_X1 port map( D => n2769, CK => CLK, Q => n_2782, QN 
                           => n30025);
   clk_r_REG8847_S1 : DFF_X1 port map( D => n2959, CK => CLK, Q => n_2783, QN 
                           => n30024);
   clk_r_REG9672_S1 : DFF_X1 port map( D => n2705, CK => CLK, Q => n_2784, QN 
                           => n30023);
   clk_r_REG9498_S1 : DFF_X1 port map( D => n2609, CK => CLK, Q => n_2785, QN 
                           => n30022);
   clk_r_REG8783_S1 : DFF_X1 port map( D => n2927, CK => CLK, Q => n_2786, QN 
                           => n30021);
   clk_r_REG8464_S1 : DFF_X1 port map( D => n3087, CK => CLK, Q => n_2787, QN 
                           => n30020);
   clk_r_REG8719_S1 : DFF_X1 port map( D => n2863, CK => CLK, Q => n_2788, QN 
                           => n30019);
   clk_r_REG9031_S1 : DFF_X1 port map( D => n2770, CK => CLK, Q => n_2789, QN 
                           => n30018);
   clk_r_REG9670_S1 : DFF_X1 port map( D => n2706, CK => CLK, Q => n_2790, QN 
                           => n30017);
   clk_r_REG7485_S1 : DFF_X1 port map( D => n3279, CK => CLK, Q => n_2791, QN 
                           => n30016);
   clk_r_REG8320_S1 : DFF_X1 port map( D => n3246, CK => CLK, Q => n_2792, QN 
                           => n30015);
   clk_r_REG9119_S1 : DFF_X1 port map( D => n3182, CK => CLK, Q => n_2793, QN 
                           => n30014);
   clk_r_REG8658_S1 : DFF_X1 port map( D => n3150, CK => CLK, Q => n_2794, QN 
                           => n30013);
   clk_r_REG8590_S1 : DFF_X1 port map( D => n3120, CK => CLK, Q => n_2795, QN 
                           => n30012);
   clk_r_REG8462_S1 : DFF_X1 port map( D => n3088, CK => CLK, Q => n_2796, QN 
                           => n30011);
   clk_r_REG9496_S1 : DFF_X1 port map( D => n2610, CK => CLK, Q => n_2797, QN 
                           => n30010);
   clk_r_REG8973_S1 : DFF_X1 port map( D => n3024, CK => CLK, Q => n_2798, QN 
                           => n30009);
   clk_r_REG8909_S1 : DFF_X1 port map( D => n2992, CK => CLK, Q => n_2799, QN 
                           => n30008);
   clk_r_REG8526_S1 : DFF_X1 port map( D => n3056, CK => CLK, Q => n_2800, QN 
                           => n30007);
   clk_r_REG8971_S1 : DFF_X1 port map( D => n3025, CK => CLK, Q => n_2801, QN 
                           => n30006);
   clk_r_REG8907_S1 : DFF_X1 port map( D => n2993, CK => CLK, Q => n_2802, QN 
                           => n30005);
   clk_r_REG8845_S1 : DFF_X1 port map( D => n2960, CK => CLK, Q => n_2803, QN 
                           => n30004);
   clk_r_REG8781_S1 : DFF_X1 port map( D => n2928, CK => CLK, Q => n_2804, QN 
                           => n30003);
   clk_r_REG8524_S1 : DFF_X1 port map( D => n3057, CK => CLK, Q => n_2805, QN 
                           => n30002);
   clk_r_REG8905_S1 : DFF_X1 port map( D => n2994, CK => CLK, Q => n_2806, QN 
                           => n30001);
   clk_r_REG8460_S1 : DFF_X1 port map( D => n3089, CK => CLK, Q => n_2807, QN 
                           => n30000);
   clk_r_REG8717_S1 : DFF_X1 port map( D => n2864, CK => CLK, Q => n_2808, QN 
                           => n29999);
   clk_r_REG8588_S1 : DFF_X1 port map( D => n3121, CK => CLK, Q => n_2809, QN 
                           => n29998);
   clk_r_REG8656_S1 : DFF_X1 port map( D => n3151, CK => CLK, Q => n_2810, QN 
                           => n29997);
   clk_r_REG9117_S1 : DFF_X1 port map( D => n3183, CK => CLK, Q => n_2811, QN 
                           => n29996);
   clk_r_REG8843_S1 : DFF_X1 port map( D => n2961, CK => CLK, Q => n_2812, QN 
                           => n29995);
   clk_r_REG8318_S1 : DFF_X1 port map( D => n3247, CK => CLK, Q => n_2813, QN 
                           => n29994);
   clk_r_REG7483_S1 : DFF_X1 port map( D => n3280, CK => CLK, Q => n_2814, QN 
                           => n29993);
   clk_r_REG8316_S1 : DFF_X1 port map( D => n3248, CK => CLK, Q => n_2815, QN 
                           => n29992);
   clk_r_REG8779_S1 : DFF_X1 port map( D => n2929, CK => CLK, Q => n_2816, QN 
                           => n29991);
   clk_r_REG9115_S1 : DFF_X1 port map( D => n3184, CK => CLK, Q => n_2817, QN 
                           => n29990);
   clk_r_REG8654_S1 : DFF_X1 port map( D => n3152, CK => CLK, Q => n_2818, QN 
                           => n29989);
   clk_r_REG8715_S1 : DFF_X1 port map( D => n2865, CK => CLK, Q => n_2819, QN 
                           => n29988);
   clk_r_REG8586_S1 : DFF_X1 port map( D => n3122, CK => CLK, Q => n_2820, QN 
                           => n29987);
   clk_r_REG8458_S1 : DFF_X1 port map( D => n3090, CK => CLK, Q => n_2821, QN 
                           => n29986);
   clk_r_REG7481_S1 : DFF_X1 port map( D => n3281, CK => CLK, Q => n_2822, QN 
                           => n29985);
   clk_r_REG9494_S1 : DFF_X1 port map( D => n2611, CK => CLK, Q => n_2823, QN 
                           => n29984);
   clk_r_REG9668_S1 : DFF_X1 port map( D => n2707, CK => CLK, Q => n_2824, QN 
                           => n29983);
   clk_r_REG9029_S1 : DFF_X1 port map( D => n2771, CK => CLK, Q => n_2825, QN 
                           => n29982);
   clk_r_REG8713_S1 : DFF_X1 port map( D => n2866, CK => CLK, Q => n_2826, QN 
                           => n29981);
   clk_r_REG8777_S1 : DFF_X1 port map( D => n2930, CK => CLK, Q => n_2827, QN 
                           => n29980);
   clk_r_REG8841_S1 : DFF_X1 port map( D => n2962, CK => CLK, Q => n_2828, QN 
                           => n29979);
   clk_r_REG8522_S1 : DFF_X1 port map( D => n3058, CK => CLK, Q => n_2829, QN 
                           => n29978);
   clk_r_REG8969_S1 : DFF_X1 port map( D => n3026, CK => CLK, Q => n_2830, QN 
                           => n29977);
   clk_r_REG8903_S1 : DFF_X1 port map( D => n2995, CK => CLK, Q => n_2831, QN 
                           => n29976);
   clk_r_REG8967_S1 : DFF_X1 port map( D => n3027, CK => CLK, Q => n_2832, QN 
                           => n29975);
   clk_r_REG8839_S1 : DFF_X1 port map( D => n2963, CK => CLK, Q => n_2833, QN 
                           => n29974);
   clk_r_REG7479_S1 : DFF_X1 port map( D => n3282, CK => CLK, Q => n_2834, QN 
                           => n29973);
   clk_r_REG8775_S1 : DFF_X1 port map( D => n2931, CK => CLK, Q => n_2835, QN 
                           => n29972);
   clk_r_REG9113_S1 : DFF_X1 port map( D => n3185, CK => CLK, Q => n_2836, QN 
                           => n29971);
   clk_r_REG8314_S1 : DFF_X1 port map( D => n3249, CK => CLK, Q => n_2837, QN 
                           => n29970);
   clk_r_REG8901_S1 : DFF_X1 port map( D => n2996, CK => CLK, Q => n_2838, QN 
                           => n29969);
   clk_r_REG7477_S1 : DFF_X1 port map( D => n3283, CK => CLK, Q => n_2839, QN 
                           => n29968);
   clk_r_REG8965_S1 : DFF_X1 port map( D => n3028, CK => CLK, Q => n_2840, QN 
                           => n29967);
   clk_r_REG8711_S1 : DFF_X1 port map( D => n2867, CK => CLK, Q => n_2841, QN 
                           => n29966);
   clk_r_REG8520_S1 : DFF_X1 port map( D => n3059, CK => CLK, Q => n_2842, QN 
                           => n29965);
   clk_r_REG9666_S1 : DFF_X1 port map( D => n2708, CK => CLK, Q => n_2843, QN 
                           => n29964);
   clk_r_REG8456_S1 : DFF_X1 port map( D => n3091, CK => CLK, Q => n_2844, QN 
                           => n29963);
   clk_r_REG8312_S1 : DFF_X1 port map( D => n3250, CK => CLK, Q => n_2845, QN 
                           => n29962);
   clk_r_REG8584_S1 : DFF_X1 port map( D => n3123, CK => CLK, Q => n_2846, QN 
                           => n29961);
   clk_r_REG9027_S1 : DFF_X1 port map( D => n2772, CK => CLK, Q => n_2847, QN 
                           => n29960);
   clk_r_REG8652_S1 : DFF_X1 port map( D => n3153, CK => CLK, Q => n_2848, QN 
                           => n29959);
   clk_r_REG8582_S1 : DFF_X1 port map( D => n3124, CK => CLK, Q => n_2849, QN 
                           => n29958);
   clk_r_REG9492_S1 : DFF_X1 port map( D => n2612, CK => CLK, Q => n_2850, QN 
                           => n29957);
   clk_r_REG8837_S1 : DFF_X1 port map( D => n2964, CK => CLK, Q => n_2851, QN 
                           => n29956);
   clk_r_REG8650_S1 : DFF_X1 port map( D => n3154, CK => CLK, Q => n_2852, QN 
                           => n29955);
   clk_r_REG8518_S1 : DFF_X1 port map( D => n3060, CK => CLK, Q => n_2853, QN 
                           => n29954);
   clk_r_REG8773_S1 : DFF_X1 port map( D => n2932, CK => CLK, Q => n_2854, QN 
                           => n29953);
   clk_r_REG9025_S1 : DFF_X1 port map( D => n2773, CK => CLK, Q => n_2855, QN 
                           => n29952);
   clk_r_REG9111_S1 : DFF_X1 port map( D => n3186, CK => CLK, Q => n_2856, QN 
                           => n29951);
   clk_r_REG8310_S1 : DFF_X1 port map( D => n3251, CK => CLK, Q => n_2857, QN 
                           => n29950);
   clk_r_REG8963_S1 : DFF_X1 port map( D => n3029, CK => CLK, Q => n_2858, QN 
                           => n29949);
   clk_r_REG7475_S1 : DFF_X1 port map( D => n3284, CK => CLK, Q => n_2859, QN 
                           => n29948);
   clk_r_REG8648_S1 : DFF_X1 port map( D => n3155, CK => CLK, Q => n_2860, QN 
                           => n29947);
   clk_r_REG8709_S1 : DFF_X1 port map( D => n2868, CK => CLK, Q => n_2861, QN 
                           => n29946);
   clk_r_REG9664_S1 : DFF_X1 port map( D => n2709, CK => CLK, Q => n_2862, QN 
                           => n29945);
   clk_r_REG9490_S1 : DFF_X1 port map( D => n2613, CK => CLK, Q => n_2863, QN 
                           => n29944);
   clk_r_REG9109_S1 : DFF_X1 port map( D => n3187, CK => CLK, Q => n_2864, QN 
                           => n29943);
   clk_r_REG8454_S1 : DFF_X1 port map( D => n3092, CK => CLK, Q => n_2865, QN 
                           => n29942);
   clk_r_REG8580_S1 : DFF_X1 port map( D => n3125, CK => CLK, Q => n_2866, QN 
                           => n29941);
   clk_r_REG8308_S1 : DFF_X1 port map( D => n3252, CK => CLK, Q => n_2867, QN 
                           => n29940);
   clk_r_REG8306_S1 : DFF_X1 port map( D => n3253, CK => CLK, Q => n_2868, QN 
                           => n29939);
   clk_r_REG8304_S1 : DFF_X1 port map( D => n3254, CK => CLK, Q => n_2869, QN 
                           => n29938);
   clk_r_REG8302_S1 : DFF_X1 port map( D => n3255, CK => CLK, Q => n_2870, QN 
                           => n29937);
   clk_r_REG8300_S1 : DFF_X1 port map( D => n3256, CK => CLK, Q => n_2871, QN 
                           => n29936);
   clk_r_REG8298_S1 : DFF_X1 port map( D => n3257, CK => CLK, Q => n_2872, QN 
                           => n29935);
   clk_r_REG8296_S1 : DFF_X1 port map( D => n3258, CK => CLK, Q => n_2873, QN 
                           => n29934);
   clk_r_REG8294_S1 : DFF_X1 port map( D => n3259, CK => CLK, Q => n_2874, QN 
                           => n29933);
   clk_r_REG9023_S1 : DFF_X1 port map( D => n2774, CK => CLK, Q => n_2875, QN 
                           => n29932);
   clk_r_REG9021_S1 : DFF_X1 port map( D => n2775, CK => CLK, Q => n_2876, QN 
                           => n29931);
   clk_r_REG9019_S1 : DFF_X1 port map( D => n2776, CK => CLK, Q => n_2877, QN 
                           => n29930);
   clk_r_REG9017_S1 : DFF_X1 port map( D => n2777, CK => CLK, Q => n_2878, QN 
                           => n29929);
   clk_r_REG9055_S1 : DFF_X1 port map( D => n2758, CK => CLK, Q => n_2879, QN 
                           => n29928);
   clk_r_REG9015_S1 : DFF_X1 port map( D => n2778, CK => CLK, Q => n_2880, QN 
                           => n29927);
   clk_r_REG9013_S1 : DFF_X1 port map( D => n2779, CK => CLK, Q => n_2881, QN 
                           => n29926);
   clk_r_REG7473_S1 : DFF_X1 port map( D => n3285, CK => CLK, Q => n_2882, QN 
                           => n29925);
   clk_r_REG7471_S1 : DFF_X1 port map( D => n3286, CK => CLK, Q => n_2883, QN 
                           => n29924);
   clk_r_REG7469_S1 : DFF_X1 port map( D => n3287, CK => CLK, Q => n_2884, QN 
                           => n29923);
   clk_r_REG7467_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n_2885, QN 
                           => n29922);
   clk_r_REG7465_S1 : DFF_X1 port map( D => n3289, CK => CLK, Q => n_2886, QN 
                           => n29921);
   clk_r_REG7503_S1 : DFF_X1 port map( D => n3270, CK => CLK, Q => n_2887, QN 
                           => n29920);
   clk_r_REG7463_S1 : DFF_X1 port map( D => n3290, CK => CLK, Q => n_2888, QN 
                           => n29919);
   clk_r_REG7461_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n_2889, QN 
                           => n29918);
   clk_r_REG9488_S1 : DFF_X1 port map( D => n2614, CK => CLK, Q => n_2890, QN 
                           => n29917);
   clk_r_REG9486_S1 : DFF_X1 port map( D => n2615, CK => CLK, Q => n_2891, QN 
                           => n29916);
   clk_r_REG9484_S1 : DFF_X1 port map( D => n2616, CK => CLK, Q => n_2892, QN 
                           => n29915);
   clk_r_REG9338_S1 : DFF_X1 port map( D => n2551, CK => CLK, Q => n_2893, QN 
                           => n29914);
   clk_r_REG9482_S1 : DFF_X1 port map( D => n2617, CK => CLK, Q => n_2894, QN 
                           => n29913);
   clk_r_REG9480_S1 : DFF_X1 port map( D => n2606, CK => CLK, Q => n_2895, QN 
                           => n29912);
   clk_r_REG9462_S1 : DFF_X1 port map( D => n2618, CK => CLK, Q => n_2896, QN 
                           => n29911);
   clk_r_REG9662_S1 : DFF_X1 port map( D => n2710, CK => CLK, Q => n_2897, QN 
                           => n29910);
   clk_r_REG9660_S1 : DFF_X1 port map( D => n2711, CK => CLK, Q => n_2898, QN 
                           => n29909);
   clk_r_REG8452_S1 : DFF_X1 port map( D => n3093, CK => CLK, Q => n_2899, QN 
                           => n29908);
   clk_r_REG8450_S1 : DFF_X1 port map( D => n3094, CK => CLK, Q => n_2900, QN 
                           => n29907);
   clk_r_REG8448_S1 : DFF_X1 port map( D => n3095, CK => CLK, Q => n_2901, QN 
                           => n29906);
   clk_r_REG8446_S1 : DFF_X1 port map( D => n3096, CK => CLK, Q => n_2902, QN 
                           => n29905);
   clk_r_REG8516_S1 : DFF_X1 port map( D => n3061, CK => CLK, Q => n_2903, QN 
                           => n29904);
   clk_r_REG8444_S1 : DFF_X1 port map( D => n3097, CK => CLK, Q => n_2904, QN 
                           => n29903);
   clk_r_REG8482_S1 : DFF_X1 port map( D => n3078, CK => CLK, Q => n_2905, QN 
                           => n29902);
   clk_r_REG8442_S1 : DFF_X1 port map( D => n3098, CK => CLK, Q => n_2906, QN 
                           => n29901);
   clk_r_REG9336_S1 : DFF_X1 port map( D => n2552, CK => CLK, Q => n_2907, QN 
                           => n29900);
   clk_r_REG9658_S1 : DFF_X1 port map( D => n2712, CK => CLK, Q => n_2908, QN 
                           => n29899);
   clk_r_REG9656_S1 : DFF_X1 port map( D => n2713, CK => CLK, Q => n_2909, QN 
                           => n29898);
   clk_r_REG9694_S1 : DFF_X1 port map( D => n2694, CK => CLK, Q => n_2910, QN 
                           => n29897);
   clk_r_REG9654_S1 : DFF_X1 port map( D => n2714, CK => CLK, Q => n_2911, QN 
                           => n29896);
   clk_r_REG9334_S1 : DFF_X1 port map( D => n2553, CK => CLK, Q => n_2912, QN 
                           => n29895);
   clk_r_REG8578_S1 : DFF_X1 port map( D => n3126, CK => CLK, Q => n_2913, QN 
                           => n29894);
   clk_r_REG8576_S1 : DFF_X1 port map( D => n3127, CK => CLK, Q => n_2914, QN 
                           => n29893);
   clk_r_REG8574_S1 : DFF_X1 port map( D => n3128, CK => CLK, Q => n_2915, QN 
                           => n29892);
   clk_r_REG9372_S1 : DFF_X1 port map( D => n2534, CK => CLK, Q => n_2916, QN 
                           => n29891);
   clk_r_REG9652_S1 : DFF_X1 port map( D => n2715, CK => CLK, Q => n_2917, QN 
                           => n29890);
   clk_r_REG9460_S1 : DFF_X1 port map( D => n2619, CK => CLK, Q => n_2918, QN 
                           => n29889);
   clk_r_REG8572_S1 : DFF_X1 port map( D => n3129, CK => CLK, Q => n_2919, QN 
                           => n29888);
   clk_r_REG8570_S1 : DFF_X1 port map( D => n3130, CK => CLK, Q => n_2920, QN 
                           => n29887);
   clk_r_REG8568_S1 : DFF_X1 port map( D => n3131, CK => CLK, Q => n_2921, QN 
                           => n29886);
   clk_r_REG8566_S1 : DFF_X1 port map( D => n3132, CK => CLK, Q => n_2922, QN 
                           => n29885);
   clk_r_REG8564_S1 : DFF_X1 port map( D => n3133, CK => CLK, Q => n_2923, QN 
                           => n29884);
   clk_r_REG8646_S1 : DFF_X1 port map( D => n3156, CK => CLK, Q => n_2924, QN 
                           => n29883);
   clk_r_REG8644_S1 : DFF_X1 port map( D => n3157, CK => CLK, Q => n_2925, QN 
                           => n29882);
   clk_r_REG8835_S1 : DFF_X1 port map( D => n2965, CK => CLK, Q => n_2926, QN 
                           => n29881);
   clk_r_REG9332_S1 : DFF_X1 port map( D => n2554, CK => CLK, Q => n_2927, QN 
                           => n29880);
   clk_r_REG8642_S1 : DFF_X1 port map( D => n3158, CK => CLK, Q => n_2928, QN 
                           => n29879);
   clk_r_REG8640_S1 : DFF_X1 port map( D => n3159, CK => CLK, Q => n_2929, QN 
                           => n29878);
   clk_r_REG8638_S1 : DFF_X1 port map( D => n3160, CK => CLK, Q => n_2930, QN 
                           => n29877);
   clk_r_REG8636_S1 : DFF_X1 port map( D => n3161, CK => CLK, Q => n_2931, QN 
                           => n29876);
   clk_r_REG8634_S1 : DFF_X1 port map( D => n3162, CK => CLK, Q => n_2932, QN 
                           => n29875);
   clk_r_REG8632_S1 : DFF_X1 port map( D => n3163, CK => CLK, Q => n_2933, QN 
                           => n29874);
   clk_r_REG8899_S1 : DFF_X1 port map( D => n2997, CK => CLK, Q => n_2934, QN 
                           => n29873);
   clk_r_REG9330_S1 : DFF_X1 port map( D => n2555, CK => CLK, Q => n_2935, QN 
                           => n29872);
   clk_r_REG9107_S1 : DFF_X1 port map( D => n3188, CK => CLK, Q => n_2936, QN 
                           => n29871);
   clk_r_REG9105_S1 : DFF_X1 port map( D => n3189, CK => CLK, Q => n_2937, QN 
                           => n29870);
   clk_r_REG9103_S1 : DFF_X1 port map( D => n3190, CK => CLK, Q => n_2938, QN 
                           => n29869);
   clk_r_REG9101_S1 : DFF_X1 port map( D => n3191, CK => CLK, Q => n_2939, QN 
                           => n29868);
   clk_r_REG9099_S1 : DFF_X1 port map( D => n3192, CK => CLK, Q => n_2940, QN 
                           => n29867);
   clk_r_REG8771_S1 : DFF_X1 port map( D => n2933, CK => CLK, Q => n_2941, QN 
                           => n29866);
   clk_r_REG9097_S1 : DFF_X1 port map( D => n3193, CK => CLK, Q => n_2942, QN 
                           => n29865);
   clk_r_REG9095_S1 : DFF_X1 port map( D => n3194, CK => CLK, Q => n_2943, QN 
                           => n29864);
   clk_r_REG8961_S1 : DFF_X1 port map( D => n3030, CK => CLK, Q => n_2944, QN 
                           => n29863);
   clk_r_REG8959_S1 : DFF_X1 port map( D => n3031, CK => CLK, Q => n_2945, QN 
                           => n29862);
   clk_r_REG8957_S1 : DFF_X1 port map( D => n3032, CK => CLK, Q => n_2946, QN 
                           => n29861);
   clk_r_REG8955_S1 : DFF_X1 port map( D => n3033, CK => CLK, Q => n_2947, QN 
                           => n29860);
   clk_r_REG8953_S1 : DFF_X1 port map( D => n3034, CK => CLK, Q => n_2948, QN 
                           => n29859);
   clk_r_REG8951_S1 : DFF_X1 port map( D => n3035, CK => CLK, Q => n_2949, QN 
                           => n29858);
   clk_r_REG9093_S1 : DFF_X1 port map( D => n3195, CK => CLK, Q => n_2950, QN 
                           => n29857);
   clk_r_REG8949_S1 : DFF_X1 port map( D => n3036, CK => CLK, Q => n_2951, QN 
                           => n29856);
   clk_r_REG8707_S1 : DFF_X1 port map( D => n2869, CK => CLK, Q => n_2952, QN 
                           => n29855);
   clk_r_REG8769_S1 : DFF_X1 port map( D => n2934, CK => CLK, Q => n_2953, QN 
                           => n29854);
   clk_r_REG8705_S1 : DFF_X1 port map( D => n2870, CK => CLK, Q => n_2954, QN 
                           => n29853);
   clk_r_REG8703_S1 : DFF_X1 port map( D => n2871, CK => CLK, Q => n_2955, QN 
                           => n29852);
   clk_r_REG8767_S1 : DFF_X1 port map( D => n2935, CK => CLK, Q => n_2956, QN 
                           => n29851);
   clk_r_REG8701_S1 : DFF_X1 port map( D => n2872, CK => CLK, Q => n_2957, QN 
                           => n29850);
   clk_r_REG8699_S1 : DFF_X1 port map( D => n2873, CK => CLK, Q => n_2958, QN 
                           => n29849);
   clk_r_REG8737_S1 : DFF_X1 port map( D => n2854, CK => CLK, Q => n_2959, QN 
                           => n29848);
   clk_r_REG8697_S1 : DFF_X1 port map( D => n2874, CK => CLK, Q => n_2960, QN 
                           => n29847);
   clk_r_REG8695_S1 : DFF_X1 port map( D => n2875, CK => CLK, Q => n_2961, QN 
                           => n29846);
   clk_r_REG8833_S1 : DFF_X1 port map( D => n2966, CK => CLK, Q => n_2962, QN 
                           => n29845);
   clk_r_REG8831_S1 : DFF_X1 port map( D => n2967, CK => CLK, Q => n_2963, QN 
                           => n29844);
   clk_r_REG8829_S1 : DFF_X1 port map( D => n2968, CK => CLK, Q => n_2964, QN 
                           => n29843);
   clk_r_REG8827_S1 : DFF_X1 port map( D => n2969, CK => CLK, Q => n_2965, QN 
                           => n29842);
   clk_r_REG8865_S1 : DFF_X1 port map( D => n2950, CK => CLK, Q => n_2966, QN 
                           => n29841);
   clk_r_REG8825_S1 : DFF_X1 port map( D => n2970, CK => CLK, Q => n_2967, QN 
                           => n29840);
   clk_r_REG8823_S1 : DFF_X1 port map( D => n2971, CK => CLK, Q => n_2968, QN 
                           => n29839);
   clk_r_REG8765_S1 : DFF_X1 port map( D => n2936, CK => CLK, Q => n_2969, QN 
                           => n29838);
   clk_r_REG8763_S1 : DFF_X1 port map( D => n2937, CK => CLK, Q => n_2970, QN 
                           => n29837);
   clk_r_REG8801_S1 : DFF_X1 port map( D => n2918, CK => CLK, Q => n_2971, QN 
                           => n29836);
   clk_r_REG8761_S1 : DFF_X1 port map( D => n2938, CK => CLK, Q => n_2972, QN 
                           => n29835);
   clk_r_REG8759_S1 : DFF_X1 port map( D => n2939, CK => CLK, Q => n_2973, QN 
                           => n29834);
   clk_r_REG9960_S1 : DFF_X1 port map( D => n3535, CK => CLK, Q => n_2974, QN 
                           => n29833);
   clk_r_REG9958_S1 : DFF_X1 port map( D => n3536, CK => CLK, Q => n_2975, QN 
                           => n29832);
   clk_r_REG9956_S1 : DFF_X1 port map( D => n3537, CK => CLK, Q => n_2976, QN 
                           => n29831);
   clk_r_REG9954_S1 : DFF_X1 port map( D => n3538, CK => CLK, Q => n_2977, QN 
                           => n29830);
   clk_r_REG9952_S1 : DFF_X1 port map( D => n3539, CK => CLK, Q => n_2978, QN 
                           => n29829);
   clk_r_REG9950_S1 : DFF_X1 port map( D => n3540, CK => CLK, Q => n_2979, QN 
                           => n29828);
   clk_r_REG7997_S1 : DFF_X1 port map( D => n3375, CK => CLK, Q => n_2980, QN 
                           => n29827);
   clk_r_REG7995_S1 : DFF_X1 port map( D => n3376, CK => CLK, Q => n_2981, QN 
                           => n29826);
   clk_r_REG7993_S1 : DFF_X1 port map( D => n3377, CK => CLK, Q => n_2982, QN 
                           => n29825);
   clk_r_REG7991_S1 : DFF_X1 port map( D => n3378, CK => CLK, Q => n_2983, QN 
                           => n29824);
   clk_r_REG7701_S1 : DFF_X1 port map( D => n3343, CK => CLK, Q => n_2984, QN 
                           => n29823);
   clk_r_REG7699_S1 : DFF_X1 port map( D => n3344, CK => CLK, Q => n_2985, QN 
                           => n29822);
   clk_r_REG8514_S1 : DFF_X1 port map( D => n3062, CK => CLK, Q => n_2986, QN 
                           => n29821);
   clk_r_REG7697_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n_2987, QN 
                           => n29820);
   clk_r_REG7695_S1 : DFF_X1 port map( D => n3346, CK => CLK, Q => n_2988, QN 
                           => n29819);
   clk_r_REG7693_S1 : DFF_X1 port map( D => n3347, CK => CLK, Q => n_2989, QN 
                           => n29818);
   clk_r_REG7989_S1 : DFF_X1 port map( D => n3379, CK => CLK, Q => n_2990, QN 
                           => n29817);
   clk_r_REG8512_S1 : DFF_X1 port map( D => n3063, CK => CLK, Q => n_2991, QN 
                           => n29816);
   clk_r_REG8510_S1 : DFF_X1 port map( D => n3064, CK => CLK, Q => n_2992, QN 
                           => n29815);
   clk_r_REG7987_S1 : DFF_X1 port map( D => n3380, CK => CLK, Q => n_2993, QN 
                           => n29814);
   clk_r_REG7691_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n_2994, QN 
                           => n29813);
   clk_r_REG8508_S1 : DFF_X1 port map( D => n3065, CK => CLK, Q => n_2995, QN 
                           => n29812);
   clk_r_REG8546_S1 : DFF_X1 port map( D => n3046, CK => CLK, Q => n_2996, QN 
                           => n29811);
   clk_r_REG8506_S1 : DFF_X1 port map( D => n3066, CK => CLK, Q => n_2997, QN 
                           => n29810);
   clk_r_REG7985_S1 : DFF_X1 port map( D => n3381, CK => CLK, Q => n_2998, QN 
                           => n29809);
   clk_r_REG9871_S1 : DFF_X1 port map( D => n3439, CK => CLK, Q => n_2999, QN 
                           => n29808);
   clk_r_REG9869_S1 : DFF_X1 port map( D => n3440, CK => CLK, Q => n_3000, QN 
                           => n29807);
   clk_r_REG7983_S1 : DFF_X1 port map( D => n3382, CK => CLK, Q => n_3001, QN 
                           => n29806);
   clk_r_REG7689_S1 : DFF_X1 port map( D => n3349, CK => CLK, Q => n_3002, QN 
                           => n29805);
   clk_r_REG9867_S1 : DFF_X1 port map( D => n3441, CK => CLK, Q => n_3003, QN 
                           => n29804);
   clk_r_REG7915_S1 : DFF_X1 port map( D => n3407, CK => CLK, Q => n_3004, QN 
                           => n29803);
   clk_r_REG7913_S1 : DFF_X1 port map( D => n3408, CK => CLK, Q => n_3005, QN 
                           => n29802);
   clk_r_REG8256_S1 : DFF_X1 port map( D => n3471, CK => CLK, Q => n_3006, QN 
                           => n29801);
   clk_r_REG8254_S1 : DFF_X1 port map( D => n3472, CK => CLK, Q => n_3007, QN 
                           => n29800);
   clk_r_REG8504_S1 : DFF_X1 port map( D => n3067, CK => CLK, Q => n_3008, QN 
                           => n29799);
   clk_r_REG7911_S1 : DFF_X1 port map( D => n3409, CK => CLK, Q => n_3009, QN 
                           => n29798);
   clk_r_REG8252_S1 : DFF_X1 port map( D => n3473, CK => CLK, Q => n_3010, QN 
                           => n29797);
   clk_r_REG9865_S1 : DFF_X1 port map( D => n3442, CK => CLK, Q => n_3011, QN 
                           => n29796);
   clk_r_REG9863_S1 : DFF_X1 port map( D => n3443, CK => CLK, Q => n_3012, QN 
                           => n29795);
   clk_r_REG9861_S1 : DFF_X1 port map( D => n3444, CK => CLK, Q => n_3013, QN 
                           => n29794);
   clk_r_REG9859_S1 : DFF_X1 port map( D => n3445, CK => CLK, Q => n_3014, QN 
                           => n29793);
   clk_r_REG7909_S1 : DFF_X1 port map( D => n3410, CK => CLK, Q => n_3015, QN 
                           => n29792);
   clk_r_REG7907_S1 : DFF_X1 port map( D => n3411, CK => CLK, Q => n_3016, QN 
                           => n29791);
   clk_r_REG8396_S1 : DFF_X1 port map( D => n3503, CK => CLK, Q => n_3017, QN 
                           => n29790);
   clk_r_REG8250_S1 : DFF_X1 port map( D => n3474, CK => CLK, Q => n_3018, QN 
                           => n29789);
   clk_r_REG8248_S1 : DFF_X1 port map( D => n3475, CK => CLK, Q => n_3019, QN 
                           => n29788);
   clk_r_REG9857_S1 : DFF_X1 port map( D => n3446, CK => CLK, Q => n_3020, QN 
                           => n29787);
   clk_r_REG8394_S1 : DFF_X1 port map( D => n3504, CK => CLK, Q => n_3021, QN 
                           => n29786);
   clk_r_REG7905_S1 : DFF_X1 port map( D => n3412, CK => CLK, Q => n_3022, QN 
                           => n29785);
   clk_r_REG7687_S1 : DFF_X1 port map( D => n3350, CK => CLK, Q => n_3023, QN 
                           => n29784);
   clk_r_REG8392_S1 : DFF_X1 port map( D => n3505, CK => CLK, Q => n_3024, QN 
                           => n29783);
   clk_r_REG8390_S1 : DFF_X1 port map( D => n3506, CK => CLK, Q => n_3025, QN 
                           => n29782);
   clk_r_REG8388_S1 : DFF_X1 port map( D => n3507, CK => CLK, Q => n_3026, QN 
                           => n29781);
   clk_r_REG8386_S1 : DFF_X1 port map( D => n3508, CK => CLK, Q => n_3027, QN 
                           => n29780);
   clk_r_REG8246_S1 : DFF_X1 port map( D => n3476, CK => CLK, Q => n_3028, QN 
                           => n29779);
   clk_r_REG8440_S1 : DFF_X1 port map( D => n3099, CK => CLK, Q => n_3029, QN 
                           => n29778);
   clk_r_REG8244_S1 : DFF_X1 port map( D => n3477, CK => CLK, Q => n_3030, QN 
                           => n29777);
   clk_r_REG8242_S1 : DFF_X1 port map( D => n3478, CK => CLK, Q => n_3031, QN 
                           => n29776);
   clk_r_REG7903_S1 : DFF_X1 port map( D => n3413, CK => CLK, Q => n_3032, QN 
                           => n29775);
   clk_r_REG8897_S1 : DFF_X1 port map( D => n2998, CK => CLK, Q => n_3033, QN 
                           => n29774);
   clk_r_REG8384_S1 : DFF_X1 port map( D => n3509, CK => CLK, Q => n_3034, QN 
                           => n29773);
   clk_r_REG8895_S1 : DFF_X1 port map( D => n2999, CK => CLK, Q => n_3035, QN 
                           => n29772);
   clk_r_REG7901_S1 : DFF_X1 port map( D => n3414, CK => CLK, Q => n_3036, QN 
                           => n29771);
   clk_r_REG8893_S1 : DFF_X1 port map( D => n3000, CK => CLK, Q => n_3037, QN 
                           => n29770);
   clk_r_REG8947_S1 : DFF_X1 port map( D => n3037, CK => CLK, Q => n_3038, QN 
                           => n29769);
   clk_r_REG8891_S1 : DFF_X1 port map( D => n3001, CK => CLK, Q => n_3039, QN 
                           => n29768);
   clk_r_REG8382_S1 : DFF_X1 port map( D => n3510, CK => CLK, Q => n_3040, QN 
                           => n29767);
   clk_r_REG8929_S1 : DFF_X1 port map( D => n2982, CK => CLK, Q => n_3041, QN 
                           => n29766);
   clk_r_REG8889_S1 : DFF_X1 port map( D => n3002, CK => CLK, Q => n_3042, QN 
                           => n29765);
   clk_r_REG8887_S1 : DFF_X1 port map( D => n3003, CK => CLK, Q => n_3043, QN 
                           => n29764);
   clk_r_REG9948_S1 : DFF_X1 port map( D => n3541, CK => CLK, Q => n_3044, QN 
                           => n29763);
   clk_r_REG9946_S1 : DFF_X1 port map( D => n3542, CK => CLK, Q => n_3045, QN 
                           => n29762);
   clk_r_REG9944_S1 : DFF_X1 port map( D => n3543, CK => CLK, Q => n_3046, QN 
                           => n29761);
   clk_r_REG9942_S1 : DFF_X1 port map( D => n3544, CK => CLK, Q => n_3047, QN 
                           => n29760);
   clk_r_REG9940_S1 : DFF_X1 port map( D => n3545, CK => CLK, Q => n_3048, QN 
                           => n29759);
   clk_r_REG9978_S1 : DFF_X1 port map( D => n3526, CK => CLK, Q => n_3049, QN 
                           => n29758);
   clk_r_REG9938_S1 : DFF_X1 port map( D => n3546, CK => CLK, Q => n_3050, QN 
                           => n29757);
   clk_r_REG9936_S1 : DFF_X1 port map( D => n3547, CK => CLK, Q => n_3051, QN 
                           => n29756);
   clk_r_REG9855_S1 : DFF_X1 port map( D => n3447, CK => CLK, Q => n_3052, QN 
                           => n29755);
   clk_r_REG7685_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n_3053, QN 
                           => n29754);
   clk_r_REG8380_S1 : DFF_X1 port map( D => n3511, CK => CLK, Q => n_3054, QN 
                           => n29753);
   clk_r_REG7981_S1 : DFF_X1 port map( D => n3383, CK => CLK, Q => n_3055, QN 
                           => n29752);
   clk_r_REG7979_S1 : DFF_X1 port map( D => n3384, CK => CLK, Q => n_3056, QN 
                           => n29751);
   clk_r_REG7899_S1 : DFF_X1 port map( D => n3415, CK => CLK, Q => n_3057, QN 
                           => n29750);
   clk_r_REG9853_S1 : DFF_X1 port map( D => n3448, CK => CLK, Q => n_3058, QN 
                           => n29749);
   clk_r_REG8240_S1 : DFF_X1 port map( D => n3479, CK => CLK, Q => n_3059, QN 
                           => n29748);
   clk_r_REG8378_S1 : DFF_X1 port map( D => n3512, CK => CLK, Q => n_3060, QN 
                           => n29747);
   clk_r_REG8376_S1 : DFF_X1 port map( D => n3513, CK => CLK, Q => n_3061, QN 
                           => n29746);
   clk_r_REG7683_S1 : DFF_X1 port map( D => n3352, CK => CLK, Q => n_3062, QN 
                           => n29745);
   clk_r_REG7681_S1 : DFF_X1 port map( D => n3353, CK => CLK, Q => n_3063, QN 
                           => n29744);
   clk_r_REG8238_S1 : DFF_X1 port map( D => n3480, CK => CLK, Q => n_3064, QN 
                           => n29743);
   clk_r_REG8414_S1 : DFF_X1 port map( D => n3494, CK => CLK, Q => n_3065, QN 
                           => n29742);
   clk_r_REG8236_S1 : DFF_X1 port map( D => n3481, CK => CLK, Q => n_3066, QN 
                           => n29741);
   clk_r_REG9851_S1 : DFF_X1 port map( D => n3449, CK => CLK, Q => n_3067, QN 
                           => n29740);
   clk_r_REG8374_S1 : DFF_X1 port map( D => n3514, CK => CLK, Q => n_3068, QN 
                           => n29739);
   clk_r_REG7897_S1 : DFF_X1 port map( D => n3416, CK => CLK, Q => n_3069, QN 
                           => n29738);
   clk_r_REG7977_S1 : DFF_X1 port map( D => n3385, CK => CLK, Q => n_3070, QN 
                           => n29737);
   clk_r_REG7719_S1 : DFF_X1 port map( D => n3334, CK => CLK, Q => n_3071, QN 
                           => n29736);
   clk_r_REG7895_S1 : DFF_X1 port map( D => n3417, CK => CLK, Q => n_3072, QN 
                           => n29735);
   clk_r_REG8015_S1 : DFF_X1 port map( D => n3366, CK => CLK, Q => n_3073, QN 
                           => n29734);
   clk_r_REG7933_S1 : DFF_X1 port map( D => n3398, CK => CLK, Q => n_3074, QN 
                           => n29733);
   clk_r_REG7975_S1 : DFF_X1 port map( D => n3386, CK => CLK, Q => n_3075, QN 
                           => n29732);
   clk_r_REG8274_S1 : DFF_X1 port map( D => n3462, CK => CLK, Q => n_3076, QN 
                           => n29731);
   clk_r_REG7893_S1 : DFF_X1 port map( D => n3418, CK => CLK, Q => n_3077, QN 
                           => n29730);
   clk_r_REG7891_S1 : DFF_X1 port map( D => n3419, CK => CLK, Q => n_3078, QN 
                           => n29729);
   clk_r_REG7679_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n_3079, QN 
                           => n29728);
   clk_r_REG9889_S1 : DFF_X1 port map( D => n3430, CK => CLK, Q => n_3080, QN 
                           => n29727);
   clk_r_REG7677_S1 : DFF_X1 port map( D => n3355, CK => CLK, Q => n_3081, QN 
                           => n29726);
   clk_r_REG8234_S1 : DFF_X1 port map( D => n3482, CK => CLK, Q => n_3082, QN 
                           => n29725);
   clk_r_REG9849_S1 : DFF_X1 port map( D => n3450, CK => CLK, Q => n_3083, QN 
                           => n29724);
   clk_r_REG7973_S1 : DFF_X1 port map( D => n3387, CK => CLK, Q => n_3084, QN 
                           => n29723);
   clk_r_REG8372_S1 : DFF_X1 port map( D => n3515, CK => CLK, Q => n_3085, QN 
                           => n29722);
   clk_r_REG9847_S1 : DFF_X1 port map( D => n3451, CK => CLK, Q => n_3086, QN 
                           => n29721);
   clk_r_REG8232_S1 : DFF_X1 port map( D => n3483, CK => CLK, Q => n_3087, QN 
                           => n29720);
   clk_r_REG9164_S1 : DFF_X1 port map( D => n3215, CK => CLK, Q => n_3088, QN 
                           => n29719);
   clk_r_REG9162_S1 : DFF_X1 port map( D => n3216, CK => CLK, Q => n_3089, QN 
                           => n29718);
   clk_r_REG9160_S1 : DFF_X1 port map( D => n3217, CK => CLK, Q => n_3090, QN 
                           => n29717);
   clk_r_REG9158_S1 : DFF_X1 port map( D => n3218, CK => CLK, Q => n_3091, QN 
                           => n29716);
   clk_r_REG9156_S1 : DFF_X1 port map( D => n3219, CK => CLK, Q => n_3092, QN 
                           => n29715);
   clk_r_REG9154_S1 : DFF_X1 port map( D => n3220, CK => CLK, Q => n_3093, QN 
                           => n29714);
   clk_r_REG9328_S1 : DFF_X1 port map( D => n2556, CK => CLK, Q => n_3094, QN 
                           => n29713);
   clk_r_REG9011_S1 : DFF_X1 port map( D => n2780, CK => CLK, Q => n_3095, QN 
                           => n29712);
   clk_r_REG8292_S1 : DFF_X1 port map( D => n3260, CK => CLK, Q => n_3096, QN 
                           => n29711);
   clk_r_REG9152_S1 : DFF_X1 port map( D => n3221, CK => CLK, Q => n_3097, QN 
                           => n29710);
   clk_r_REG8821_S1 : DFF_X1 port map( D => n2972, CK => CLK, Q => n_3098, QN 
                           => n29709);
   clk_r_REG8562_S1 : DFF_X1 port map( D => n3134, CK => CLK, Q => n_3099, QN 
                           => n29708);
   clk_r_REG9458_S1 : DFF_X1 port map( D => n2620, CK => CLK, Q => n_3100, QN 
                           => n29707);
   clk_r_REG9456_S1 : DFF_X1 port map( D => n2621, CK => CLK, Q => n_3101, QN 
                           => n29706);
   clk_r_REG7459_S1 : DFF_X1 port map( D => n3292, CK => CLK, Q => n_3102, QN 
                           => n29705);
   clk_r_REG9650_S1 : DFF_X1 port map( D => n2716, CK => CLK, Q => n_3103, QN 
                           => n29704);
   clk_r_REG9091_S1 : DFF_X1 port map( D => n3196, CK => CLK, Q => n_3104, QN 
                           => n29703);
   clk_r_REG8290_S1 : DFF_X1 port map( D => n3261, CK => CLK, Q => n_3105, QN 
                           => n29702);
   clk_r_REG8560_S1 : DFF_X1 port map( D => n3135, CK => CLK, Q => n_3106, QN 
                           => n29701);
   clk_r_REG9089_S1 : DFF_X1 port map( D => n3197, CK => CLK, Q => n_3107, QN 
                           => n29700);
   clk_r_REG8630_S1 : DFF_X1 port map( D => n3164, CK => CLK, Q => n_3108, QN 
                           => n29699);
   clk_r_REG8693_S1 : DFF_X1 port map( D => n2876, CK => CLK, Q => n_3109, QN 
                           => n29698);
   clk_r_REG8945_S1 : DFF_X1 port map( D => n3038, CK => CLK, Q => n_3110, QN 
                           => n29697);
   clk_r_REG9454_S1 : DFF_X1 port map( D => n2622, CK => CLK, Q => n_3111, QN 
                           => n29696);
   clk_r_REG8438_S1 : DFF_X1 port map( D => n3100, CK => CLK, Q => n_3112, QN 
                           => n29695);
   clk_r_REG9326_S1 : DFF_X1 port map( D => n2557, CK => CLK, Q => n_3113, QN 
                           => n29694);
   clk_r_REG8943_S1 : DFF_X1 port map( D => n3039, CK => CLK, Q => n_3114, QN 
                           => n29693);
   clk_r_REG9009_S1 : DFF_X1 port map( D => n2781, CK => CLK, Q => n_3115, QN 
                           => n29692);
   clk_r_REG8610_S1 : DFF_X1 port map( D => n3110, CK => CLK, Q => n_3116, QN 
                           => n29691);
   clk_r_REG8757_S1 : DFF_X1 port map( D => n2940, CK => CLK, Q => n_3117, QN 
                           => n29690);
   clk_r_REG8819_S1 : DFF_X1 port map( D => n2973, CK => CLK, Q => n_3118, QN 
                           => n29689);
   clk_r_REG8755_S1 : DFF_X1 port map( D => n2941, CK => CLK, Q => n_3119, QN 
                           => n29688);
   clk_r_REG8691_S1 : DFF_X1 port map( D => n2877, CK => CLK, Q => n_3120, QN 
                           => n29687);
   clk_r_REG9150_S1 : DFF_X1 port map( D => n3222, CK => CLK, Q => n_3121, QN 
                           => n29686);
   clk_r_REG8753_S1 : DFF_X1 port map( D => n2942, CK => CLK, Q => n_3122, QN 
                           => n29685);
   clk_r_REG9007_S1 : DFF_X1 port map( D => n2782, CK => CLK, Q => n_3123, QN 
                           => n29684);
   clk_r_REG9087_S1 : DFF_X1 port map( D => n3198, CK => CLK, Q => n_3124, QN 
                           => n29683);
   clk_r_REG9648_S1 : DFF_X1 port map( D => n2717, CK => CLK, Q => n_3125, QN 
                           => n29682);
   clk_r_REG9646_S1 : DFF_X1 port map( D => n2718, CK => CLK, Q => n_3126, QN 
                           => n29681);
   clk_r_REG8993_S1 : DFF_X1 port map( D => n3014, CK => CLK, Q => n_3127, QN 
                           => n29680);
   clk_r_REG8817_S1 : DFF_X1 port map( D => n2974, CK => CLK, Q => n_3128, QN 
                           => n29679);
   clk_r_REG7457_S1 : DFF_X1 port map( D => n3293, CK => CLK, Q => n_3129, QN 
                           => n29678);
   clk_r_REG8288_S1 : DFF_X1 port map( D => n3262, CK => CLK, Q => n_3130, QN 
                           => n29677);
   clk_r_REG9148_S1 : DFF_X1 port map( D => n3223, CK => CLK, Q => n_3131, QN 
                           => n29676);
   clk_r_REG9324_S1 : DFF_X1 port map( D => n2558, CK => CLK, Q => n_3132, QN 
                           => n29675);
   clk_r_REG8436_S1 : DFF_X1 port map( D => n3101, CK => CLK, Q => n_3133, QN 
                           => n29674);
   clk_r_REG7455_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n_3134, QN 
                           => n29673);
   clk_r_REG8434_S1 : DFF_X1 port map( D => n3102, CK => CLK, Q => n_3135, QN 
                           => n29672);
   clk_r_REG8689_S1 : DFF_X1 port map( D => n2878, CK => CLK, Q => n_3136, QN 
                           => n29671);
   clk_r_REG8628_S1 : DFF_X1 port map( D => n3165, CK => CLK, Q => n_3137, QN 
                           => n29670);
   clk_r_REG8626_S1 : DFF_X1 port map( D => n3166, CK => CLK, Q => n_3138, QN 
                           => n29669);
   clk_r_REG7611_S1 : DFF_X1 port map( D => n3310, CK => CLK, Q => n_3139, QN 
                           => n29668);
   clk_r_REG7609_S1 : DFF_X1 port map( D => n3311, CK => CLK, Q => n_3140, QN 
                           => n29667);
   clk_r_REG7607_S1 : DFF_X1 port map( D => n3312, CK => CLK, Q => n_3141, QN 
                           => n29666);
   clk_r_REG7605_S1 : DFF_X1 port map( D => n3313, CK => CLK, Q => n_3142, QN 
                           => n29665);
   clk_r_REG7603_S1 : DFF_X1 port map( D => n3314, CK => CLK, Q => n_3143, QN 
                           => n29664);
   clk_r_REG7601_S1 : DFF_X1 port map( D => n3315, CK => CLK, Q => n_3144, QN 
                           => n29663);
   clk_r_REG9422_S1 : DFF_X1 port map( D => n2574, CK => CLK, Q => n_3145, QN 
                           => n29662);
   clk_r_REG9614_S1 : DFF_X1 port map( D => n2670, CK => CLK, Q => n_3146, QN 
                           => n29661);
   clk_r_REG9230_S1 : DFF_X1 port map( D => n2798, CK => CLK, Q => n_3147, QN 
                           => n29660);
   clk_r_REG9740_S1 : DFF_X1 port map( D => n2735, CK => CLK, Q => n_3148, QN 
                           => n29659);
   clk_r_REG9294_S1 : DFF_X1 port map( D => n2830, CK => CLK, Q => n_3149, QN 
                           => n29658);
   clk_r_REG9228_S1 : DFF_X1 port map( D => n2799, CK => CLK, Q => n_3150, QN 
                           => n29657);
   clk_r_REG9292_S1 : DFF_X1 port map( D => n2831, CK => CLK, Q => n_3151, QN 
                           => n29656);
   clk_r_REG9420_S1 : DFF_X1 port map( D => n2575, CK => CLK, Q => n_3152, QN 
                           => n29655);
   clk_r_REG9550_S1 : DFF_X1 port map( D => n2638, CK => CLK, Q => n_3153, QN 
                           => n29654);
   clk_r_REG9612_S1 : DFF_X1 port map( D => n2671, CK => CLK, Q => n_3154, QN 
                           => n29653);
   clk_r_REG9738_S1 : DFF_X1 port map( D => n2736, CK => CLK, Q => n_3155, QN 
                           => n29652);
   clk_r_REG9226_S1 : DFF_X1 port map( D => n2800, CK => CLK, Q => n_3156, QN 
                           => n29651);
   clk_r_REG9290_S1 : DFF_X1 port map( D => n2832, CK => CLK, Q => n_3157, QN 
                           => n29650);
   clk_r_REG9224_S1 : DFF_X1 port map( D => n2801, CK => CLK, Q => n_3158, QN 
                           => n29649);
   clk_r_REG9418_S1 : DFF_X1 port map( D => n2576, CK => CLK, Q => n_3159, QN 
                           => n29648);
   clk_r_REG9548_S1 : DFF_X1 port map( D => n2639, CK => CLK, Q => n_3160, QN 
                           => n29647);
   clk_r_REG9610_S1 : DFF_X1 port map( D => n2672, CK => CLK, Q => n_3161, QN 
                           => n29646);
   clk_r_REG9736_S1 : DFF_X1 port map( D => n2737, CK => CLK, Q => n_3162, QN 
                           => n29645);
   clk_r_REG9222_S1 : DFF_X1 port map( D => n2802, CK => CLK, Q => n_3163, QN 
                           => n29644);
   clk_r_REG9288_S1 : DFF_X1 port map( D => n2833, CK => CLK, Q => n_3164, QN 
                           => n29643);
   clk_r_REG9286_S1 : DFF_X1 port map( D => n2834, CK => CLK, Q => n_3165, QN 
                           => n29642);
   clk_r_REG9806_S1 : DFF_X1 port map( D => n2894, CK => CLK, Q => n_3166, QN 
                           => n29641);
   clk_r_REG9416_S1 : DFF_X1 port map( D => n2577, CK => CLK, Q => n_3167, QN 
                           => n29640);
   clk_r_REG9546_S1 : DFF_X1 port map( D => n2640, CK => CLK, Q => n_3168, QN 
                           => n29639);
   clk_r_REG9608_S1 : DFF_X1 port map( D => n2673, CK => CLK, Q => n_3169, QN 
                           => n29638);
   clk_r_REG9734_S1 : DFF_X1 port map( D => n2738, CK => CLK, Q => n_3170, QN 
                           => n29637);
   clk_r_REG9414_S1 : DFF_X1 port map( D => n2578, CK => CLK, Q => n_3171, QN 
                           => n29636);
   clk_r_REG9544_S1 : DFF_X1 port map( D => n2641, CK => CLK, Q => n_3172, QN 
                           => n29635);
   clk_r_REG9606_S1 : DFF_X1 port map( D => n2674, CK => CLK, Q => n_3173, QN 
                           => n29634);
   clk_r_REG9732_S1 : DFF_X1 port map( D => n2739, CK => CLK, Q => n_3174, QN 
                           => n29633);
   clk_r_REG9542_S1 : DFF_X1 port map( D => n2642, CK => CLK, Q => n_3175, QN 
                           => n29632);
   clk_r_REG9604_S1 : DFF_X1 port map( D => n2675, CK => CLK, Q => n_3176, QN 
                           => n29631);
   clk_r_REG9284_S1 : DFF_X1 port map( D => n2835, CK => CLK, Q => n_3177, QN 
                           => n29630);
   clk_r_REG9282_S1 : DFF_X1 port map( D => n2836, CK => CLK, Q => n_3178, QN 
                           => n29629);
   clk_r_REG9804_S1 : DFF_X1 port map( D => n2895, CK => CLK, Q => n_3179, QN 
                           => n29628);
   clk_r_REG9412_S1 : DFF_X1 port map( D => n2579, CK => CLK, Q => n_3180, QN 
                           => n29627);
   clk_r_REG9540_S1 : DFF_X1 port map( D => n2643, CK => CLK, Q => n_3181, QN 
                           => n29626);
   clk_r_REG9602_S1 : DFF_X1 port map( D => n2676, CK => CLK, Q => n_3182, QN 
                           => n29625);
   clk_r_REG9730_S1 : DFF_X1 port map( D => n2740, CK => CLK, Q => n_3183, QN 
                           => n29624);
   clk_r_REG9600_S1 : DFF_X1 port map( D => n2677, CK => CLK, Q => n_3184, QN 
                           => n29623);
   clk_r_REG9728_S1 : DFF_X1 port map( D => n2741, CK => CLK, Q => n_3185, QN 
                           => n29622);
   clk_r_REG9220_S1 : DFF_X1 port map( D => n2803, CK => CLK, Q => n_3186, QN 
                           => n29621);
   clk_r_REG9280_S1 : DFF_X1 port map( D => n2837, CK => CLK, Q => n_3187, QN 
                           => n29620);
   clk_r_REG9538_S1 : DFF_X1 port map( D => n2644, CK => CLK, Q => n_3188, QN 
                           => n29619);
   clk_r_REG9536_S1 : DFF_X1 port map( D => n2645, CK => CLK, Q => n_3189, QN 
                           => n29618);
   clk_r_REG9598_S1 : DFF_X1 port map( D => n2678, CK => CLK, Q => n_3190, QN 
                           => n29617);
   clk_r_REG9802_S1 : DFF_X1 port map( D => n2896, CK => CLK, Q => n_3191, QN 
                           => n29616);
   clk_r_REG9410_S1 : DFF_X1 port map( D => n2580, CK => CLK, Q => n_3192, QN 
                           => n29615);
   clk_r_REG9534_S1 : DFF_X1 port map( D => n2646, CK => CLK, Q => n_3193, QN 
                           => n29614);
   clk_r_REG9278_S1 : DFF_X1 port map( D => n2838, CK => CLK, Q => n_3194, QN 
                           => n29613);
   clk_r_REG9726_S1 : DFF_X1 port map( D => n2742, CK => CLK, Q => n_3195, QN 
                           => n29612);
   clk_r_REG9408_S1 : DFF_X1 port map( D => n2581, CK => CLK, Q => n_3196, QN 
                           => n29611);
   clk_r_REG9218_S1 : DFF_X1 port map( D => n2804, CK => CLK, Q => n_3197, QN 
                           => n29610);
   clk_r_REG9216_S1 : DFF_X1 port map( D => n2805, CK => CLK, Q => n_3198, QN 
                           => n29609);
   clk_r_REG9532_S1 : DFF_X1 port map( D => n2647, CK => CLK, Q => n_3199, QN 
                           => n29608);
   clk_r_REG9214_S1 : DFF_X1 port map( D => n2806, CK => CLK, Q => n_3200, QN 
                           => n29607);
   clk_r_REG9596_S1 : DFF_X1 port map( D => n2679, CK => CLK, Q => n_3201, QN 
                           => n29606);
   clk_r_REG9724_S1 : DFF_X1 port map( D => n2743, CK => CLK, Q => n_3202, QN 
                           => n29605);
   clk_r_REG9406_S1 : DFF_X1 port map( D => n2582, CK => CLK, Q => n_3203, QN 
                           => n29604);
   clk_r_REG9800_S1 : DFF_X1 port map( D => n2897, CK => CLK, Q => n_3204, QN 
                           => n29603);
   clk_r_REG9798_S1 : DFF_X1 port map( D => n2898, CK => CLK, Q => n_3205, QN 
                           => n29602);
   clk_r_REG9796_S1 : DFF_X1 port map( D => n2899, CK => CLK, Q => n_3206, QN 
                           => n29601);
   clk_r_REG9758_S1 : DFF_X1 port map( D => n2726, CK => CLK, Q => n_3207, QN 
                           => n29600);
   clk_r_REG9404_S1 : DFF_X1 port map( D => n2583, CK => CLK, Q => n_3208, QN 
                           => n29599);
   clk_r_REG9402_S1 : DFF_X1 port map( D => n2584, CK => CLK, Q => n_3209, QN 
                           => n29598);
   clk_r_REG9594_S1 : DFF_X1 port map( D => n2680, CK => CLK, Q => n_3210, QN 
                           => n29597);
   clk_r_REG8751_S1 : DFF_X1 port map( D => n2943, CK => CLK, Q => n_3211, QN 
                           => n29596);
   clk_r_REG9452_S1 : DFF_X1 port map( D => n2623, CK => CLK, Q => n_3212, QN 
                           => n29595);
   clk_r_REG9722_S1 : DFF_X1 port map( D => n2744, CK => CLK, Q => n_3213, QN 
                           => n29594);
   clk_r_REG8624_S1 : DFF_X1 port map( D => n3167, CK => CLK, Q => n_3214, QN 
                           => n29593);
   clk_r_REG9085_S1 : DFF_X1 port map( D => n3199, CK => CLK, Q => n_3215, QN 
                           => n29592);
   clk_r_REG8687_S1 : DFF_X1 port map( D => n2879, CK => CLK, Q => n_3216, QN 
                           => n29591);
   clk_r_REG9146_S1 : DFF_X1 port map( D => n3224, CK => CLK, Q => n_3217, QN 
                           => n29590);
   clk_r_REG9276_S1 : DFF_X1 port map( D => n2839, CK => CLK, Q => n_3218, QN 
                           => n29589);
   clk_r_REG9005_S1 : DFF_X1 port map( D => n2783, CK => CLK, Q => n_3219, QN 
                           => n29588);
   clk_r_REG9644_S1 : DFF_X1 port map( D => n2719, CK => CLK, Q => n_3220, QN 
                           => n29587);
   clk_r_REG8941_S1 : DFF_X1 port map( D => n3040, CK => CLK, Q => n_3221, QN 
                           => n29586);
   clk_r_REG8558_S1 : DFF_X1 port map( D => n3136, CK => CLK, Q => n_3222, QN 
                           => n29585);
   clk_r_REG8815_S1 : DFF_X1 port map( D => n2975, CK => CLK, Q => n_3223, QN 
                           => n29584);
   clk_r_REG9530_S1 : DFF_X1 port map( D => n2648, CK => CLK, Q => n_3224, QN 
                           => n29583);
   clk_r_REG7453_S1 : DFF_X1 port map( D => n3295, CK => CLK, Q => n_3225, QN 
                           => n29582);
   clk_r_REG9212_S1 : DFF_X1 port map( D => n2807, CK => CLK, Q => n_3226, QN 
                           => n29581);
   clk_r_REG8286_S1 : DFF_X1 port map( D => n3263, CK => CLK, Q => n_3227, QN 
                           => n29580);
   clk_r_REG9322_S1 : DFF_X1 port map( D => n2559, CK => CLK, Q => n_3228, QN 
                           => n29579);
   clk_r_REG8432_S1 : DFF_X1 port map( D => n3103, CK => CLK, Q => n_3229, QN 
                           => n29578);
   clk_r_REG8430_S1 : DFF_X1 port map( D => n3104, CK => CLK, Q => n_3230, QN 
                           => n29577);
   clk_r_REG9794_S1 : DFF_X1 port map( D => n2900, CK => CLK, Q => n_3231, QN 
                           => n29576);
   clk_r_REG9792_S1 : DFF_X1 port map( D => n2901, CK => CLK, Q => n_3232, QN 
                           => n29575);
   clk_r_REG8428_S1 : DFF_X1 port map( D => n3105, CK => CLK, Q => n_3233, QN 
                           => n29574);
   clk_r_REG8749_S1 : DFF_X1 port map( D => n2944, CK => CLK, Q => n_3234, QN 
                           => n29573);
   clk_r_REG8747_S1 : DFF_X1 port map( D => n2945, CK => CLK, Q => n_3235, QN 
                           => n29572);
   clk_r_REG8745_S1 : DFF_X1 port map( D => n2946, CK => CLK, Q => n_3236, QN 
                           => n29571);
   clk_r_REG9790_S1 : DFF_X1 port map( D => n2902, CK => CLK, Q => n_3237, QN 
                           => n29570);
   clk_r_REG9210_S1 : DFF_X1 port map( D => n2808, CK => CLK, Q => n_3238, QN 
                           => n29569);
   clk_r_REG9208_S1 : DFF_X1 port map( D => n2809, CK => CLK, Q => n_3239, QN 
                           => n29568);
   clk_r_REG9206_S1 : DFF_X1 port map( D => n2810, CK => CLK, Q => n_3240, QN 
                           => n29567);
   clk_r_REG9274_S1 : DFF_X1 port map( D => n2840, CK => CLK, Q => n_3241, QN 
                           => n29566);
   clk_r_REG9272_S1 : DFF_X1 port map( D => n2841, CK => CLK, Q => n_3242, QN 
                           => n29565);
   clk_r_REG9270_S1 : DFF_X1 port map( D => n2842, CK => CLK, Q => n_3243, QN 
                           => n29564);
   clk_r_REG8813_S1 : DFF_X1 port map( D => n2976, CK => CLK, Q => n_3244, QN 
                           => n29563);
   clk_r_REG8811_S1 : DFF_X1 port map( D => n2977, CK => CLK, Q => n_3245, QN 
                           => n29562);
   clk_r_REG8809_S1 : DFF_X1 port map( D => n2978, CK => CLK, Q => n_3246, QN 
                           => n29561);
   clk_r_REG8426_S1 : DFF_X1 port map( D => n3106, CK => CLK, Q => n_3247, QN 
                           => n29560);
   clk_r_REG8807_S1 : DFF_X1 port map( D => n2979, CK => CLK, Q => n_3248, QN 
                           => n29559);
   clk_r_REG8743_S1 : DFF_X1 port map( D => n2947, CK => CLK, Q => n_3249, QN 
                           => n29558);
   clk_r_REG9788_S1 : DFF_X1 port map( D => n2903, CK => CLK, Q => n_3250, QN 
                           => n29557);
   clk_r_REG9268_S1 : DFF_X1 port map( D => n2843, CK => CLK, Q => n_3251, QN 
                           => n29556);
   clk_r_REG9204_S1 : DFF_X1 port map( D => n2811, CK => CLK, Q => n_3252, QN 
                           => n29555);
   clk_r_REG9003_S1 : DFF_X1 port map( D => n2784, CK => CLK, Q => n_3253, QN 
                           => n29554);
   clk_r_REG8424_S1 : DFF_X1 port map( D => n3107, CK => CLK, Q => n_3254, QN 
                           => n29553);
   clk_r_REG8805_S1 : DFF_X1 port map( D => n2980, CK => CLK, Q => n_3255, QN 
                           => n29552);
   clk_r_REG8741_S1 : DFF_X1 port map( D => n2948, CK => CLK, Q => n_3256, QN 
                           => n29551);
   clk_r_REG9786_S1 : DFF_X1 port map( D => n2904, CK => CLK, Q => n_3257, QN 
                           => n29550);
   clk_r_REG9266_S1 : DFF_X1 port map( D => n2844, CK => CLK, Q => n_3258, QN 
                           => n29549);
   clk_r_REG9202_S1 : DFF_X1 port map( D => n2812, CK => CLK, Q => n_3259, QN 
                           => n29548);
   clk_r_REG7451_S1 : DFF_X1 port map( D => n3296, CK => CLK, Q => n_3260, QN 
                           => n29547);
   clk_r_REG7449_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n_3261, QN 
                           => n29546);
   clk_r_REG7447_S1 : DFF_X1 port map( D => n3298, CK => CLK, Q => n_3262, QN 
                           => n29545);
   clk_r_REG8422_S1 : DFF_X1 port map( D => n3108, CK => CLK, Q => n_3263, QN 
                           => n29544);
   clk_r_REG7445_S1 : DFF_X1 port map( D => n3299, CK => CLK, Q => n_3264, QN 
                           => n29543);
   clk_r_REG7443_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n_3265, QN 
                           => n29542);
   clk_r_REG7398_S1 : DFF_X1 port map( D => n3301, CK => CLK, Q => n_3266, QN 
                           => n29541);
   clk_r_REG7131_S1 : DFF_X1 port map( D => n2981, CK => CLK, Q => n_3267, QN 
                           => n29540);
   clk_r_REG7138_S1 : DFF_X1 port map( D => n2949, CK => CLK, Q => n_3268, QN 
                           => n29539);
   clk_r_REG9784_S1 : DFF_X1 port map( D => n2905, CK => CLK, Q => n_3269, QN 
                           => n29538);
   clk_r_REG9264_S1 : DFF_X1 port map( D => n2845, CK => CLK, Q => n_3270, QN 
                           => n29537);
   clk_r_REG9200_S1 : DFF_X1 port map( D => n2813, CK => CLK, Q => n_3271, QN 
                           => n29536);
   clk_r_REG8284_S1 : DFF_X1 port map( D => n3264, CK => CLK, Q => n_3272, QN 
                           => n29535);
   clk_r_REG8282_S1 : DFF_X1 port map( D => n3265, CK => CLK, Q => n_3273, QN 
                           => n29534);
   clk_r_REG8280_S1 : DFF_X1 port map( D => n3266, CK => CLK, Q => n_3274, QN 
                           => n29533);
   clk_r_REG8278_S1 : DFF_X1 port map( D => n3267, CK => CLK, Q => n_3275, QN 
                           => n29532);
   clk_r_REG8276_S1 : DFF_X1 port map( D => n3268, CK => CLK, Q => n_3276, QN 
                           => n29531);
   clk_r_REG9144_S1 : DFF_X1 port map( D => n3225, CK => CLK, Q => n_3277, QN 
                           => n29530);
   clk_r_REG8502_S1 : DFF_X1 port map( D => n3068, CK => CLK, Q => n_3278, QN 
                           => n29529);
   clk_r_REG8500_S1 : DFF_X1 port map( D => n3069, CK => CLK, Q => n_3279, QN 
                           => n29528);
   clk_r_REG8498_S1 : DFF_X1 port map( D => n3070, CK => CLK, Q => n_3280, QN 
                           => n29527);
   clk_r_REG8496_S1 : DFF_X1 port map( D => n3071, CK => CLK, Q => n_3281, QN 
                           => n29526);
   clk_r_REG8494_S1 : DFF_X1 port map( D => n3072, CK => CLK, Q => n_3282, QN 
                           => n29525);
   clk_r_REG8492_S1 : DFF_X1 port map( D => n3073, CK => CLK, Q => n_3283, QN 
                           => n29524);
   clk_r_REG7255_S1 : DFF_X1 port map( D => n3109, CK => CLK, Q => n_3284, QN 
                           => n29523);
   clk_r_REG7328_S1 : DFF_X1 port map( D => n3269, CK => CLK, Q => n_3285, QN 
                           => n29522);
   clk_r_REG7501_S1 : DFF_X1 port map( D => n3271, CK => CLK, Q => n_3286, QN 
                           => n29521);
   clk_r_REG8608_S1 : DFF_X1 port map( D => n3111, CK => CLK, Q => n_3287, QN 
                           => n29520);
   clk_r_REG8556_S1 : DFF_X1 port map( D => n3137, CK => CLK, Q => n_3288, QN 
                           => n29519);
   clk_r_REG8554_S1 : DFF_X1 port map( D => n3138, CK => CLK, Q => n_3289, QN 
                           => n29518);
   clk_r_REG8552_S1 : DFF_X1 port map( D => n3139, CK => CLK, Q => n_3290, QN 
                           => n29517);
   clk_r_REG8550_S1 : DFF_X1 port map( D => n3140, CK => CLK, Q => n_3291, QN 
                           => n29516);
   clk_r_REG7185_S1 : DFF_X1 port map( D => n3141, CK => CLK, Q => n_3292, QN 
                           => n29515);
   clk_r_REG9198_S1 : DFF_X1 port map( D => n2814, CK => CLK, Q => n_3293, QN 
                           => n29514);
   clk_r_REG8622_S1 : DFF_X1 port map( D => n3168, CK => CLK, Q => n_3294, QN 
                           => n29513);
   clk_r_REG8620_S1 : DFF_X1 port map( D => n3169, CK => CLK, Q => n_3295, QN 
                           => n29512);
   clk_r_REG8618_S1 : DFF_X1 port map( D => n3170, CK => CLK, Q => n_3296, QN 
                           => n29511);
   clk_r_REG8616_S1 : DFF_X1 port map( D => n3171, CK => CLK, Q => n_3297, QN 
                           => n29510);
   clk_r_REG8614_S1 : DFF_X1 port map( D => n3172, CK => CLK, Q => n_3298, QN 
                           => n29509);
   clk_r_REG7167_S1 : DFF_X1 port map( D => n3173, CK => CLK, Q => n_3299, QN 
                           => n29508);
   clk_r_REG9262_S1 : DFF_X1 port map( D => n2846, CK => CLK, Q => n_3300, QN 
                           => n29507);
   clk_r_REG9782_S1 : DFF_X1 port map( D => n2906, CK => CLK, Q => n_3301, QN 
                           => n29506);
   clk_r_REG8799_S1 : DFF_X1 port map( D => n2919, CK => CLK, Q => n_3302, QN 
                           => n29505);
   clk_r_REG8863_S1 : DFF_X1 port map( D => n2951, CK => CLK, Q => n_3303, QN 
                           => n29504);
   clk_r_REG8490_S1 : DFF_X1 port map( D => n3074, CK => CLK, Q => n_3304, QN 
                           => n29503);
   clk_r_REG8480_S1 : DFF_X1 port map( D => n3079, CK => CLK, Q => n_3305, QN 
                           => n29502);
   clk_r_REG8606_S1 : DFF_X1 port map( D => n3112, CK => CLK, Q => n_3306, QN 
                           => n29501);
   clk_r_REG8674_S1 : DFF_X1 port map( D => n3142, CK => CLK, Q => n_3307, QN 
                           => n29500);
   clk_r_REG9083_S1 : DFF_X1 port map( D => n3200, CK => CLK, Q => n_3308, QN 
                           => n29499);
   clk_r_REG9081_S1 : DFF_X1 port map( D => n3201, CK => CLK, Q => n_3309, QN 
                           => n29498);
   clk_r_REG9079_S1 : DFF_X1 port map( D => n3202, CK => CLK, Q => n_3310, QN 
                           => n29497);
   clk_r_REG9077_S1 : DFF_X1 port map( D => n3203, CK => CLK, Q => n_3311, QN 
                           => n29496);
   clk_r_REG9075_S1 : DFF_X1 port map( D => n3204, CK => CLK, Q => n_3312, QN 
                           => n29495);
   clk_r_REG9073_S1 : DFF_X1 port map( D => n3205, CK => CLK, Q => n_3313, QN 
                           => n29494);
   clk_r_REG9071_S1 : DFF_X1 port map( D => n3181, CK => CLK, Q => n_3314, QN 
                           => n29493);
   clk_r_REG8336_S1 : DFF_X1 port map( D => n3238, CK => CLK, Q => n_3315, QN 
                           => n29492);
   clk_r_REG7499_S1 : DFF_X1 port map( D => n3272, CK => CLK, Q => n_3316, QN 
                           => n29491);
   clk_r_REG9182_S1 : DFF_X1 port map( D => n3206, CK => CLK, Q => n_3317, QN 
                           => n29490);
   clk_r_REG9142_S1 : DFF_X1 port map( D => n3226, CK => CLK, Q => n_3318, QN 
                           => n29489);
   clk_r_REG9140_S1 : DFF_X1 port map( D => n3227, CK => CLK, Q => n_3319, QN 
                           => n29488);
   clk_r_REG9138_S1 : DFF_X1 port map( D => n3228, CK => CLK, Q => n_3320, QN 
                           => n29487);
   clk_r_REG9136_S1 : DFF_X1 port map( D => n3229, CK => CLK, Q => n_3321, QN 
                           => n29486);
   clk_r_REG9134_S1 : DFF_X1 port map( D => n3230, CK => CLK, Q => n_3322, QN 
                           => n29485);
   clk_r_REG8334_S1 : DFF_X1 port map( D => n3239, CK => CLK, Q => n_3323, QN 
                           => n29484);
   clk_r_REG9720_S1 : DFF_X1 port map( D => n2745, CK => CLK, Q => n_3324, QN 
                           => n29483);
   clk_r_REG9718_S1 : DFF_X1 port map( D => n2746, CK => CLK, Q => n_3325, QN 
                           => n29482);
   clk_r_REG9716_S1 : DFF_X1 port map( D => n2747, CK => CLK, Q => n_3326, QN 
                           => n29481);
   clk_r_REG9714_S1 : DFF_X1 port map( D => n2748, CK => CLK, Q => n_3327, QN 
                           => n29480);
   clk_r_REG7497_S1 : DFF_X1 port map( D => n3273, CK => CLK, Q => n_3328, QN 
                           => n29479);
   clk_r_REG8332_S1 : DFF_X1 port map( D => n3240, CK => CLK, Q => n_3329, QN 
                           => n29478);
   clk_r_REG9132_S1 : DFF_X1 port map( D => n3231, CK => CLK, Q => n_3330, QN 
                           => n29477);
   clk_r_REG9069_S1 : DFF_X1 port map( D => n3180, CK => CLK, Q => n_3331, QN 
                           => n29476);
   clk_r_REG8672_S1 : DFF_X1 port map( D => n3143, CK => CLK, Q => n_3332, QN 
                           => n29475);
   clk_r_REG8604_S1 : DFF_X1 port map( D => n3113, CK => CLK, Q => n_3333, QN 
                           => n29474);
   clk_r_REG8478_S1 : DFF_X1 port map( D => n3080, CK => CLK, Q => n_3334, QN 
                           => n29473);
   clk_r_REG9642_S1 : DFF_X1 port map( D => n2720, CK => CLK, Q => n_3335, QN 
                           => n29472);
   clk_r_REG8488_S1 : DFF_X1 port map( D => n3075, CK => CLK, Q => n_3336, QN 
                           => n29471);
   clk_r_REG8861_S1 : DFF_X1 port map( D => n2952, CK => CLK, Q => n_3337, QN 
                           => n29470);
   clk_r_REG9640_S1 : DFF_X1 port map( D => n2721, CK => CLK, Q => n_3338, QN 
                           => n29469);
   clk_r_REG9638_S1 : DFF_X1 port map( D => n2722, CK => CLK, Q => n_3339, QN 
                           => n29468);
   clk_r_REG9636_S1 : DFF_X1 port map( D => n2723, CK => CLK, Q => n_3340, QN 
                           => n29467);
   clk_r_REG9634_S1 : DFF_X1 port map( D => n2724, CK => CLK, Q => n_3341, QN 
                           => n29466);
   clk_r_REG6965_S1 : DFF_X1 port map( D => n2725, CK => CLK, Q => n_3342, QN 
                           => n29465);
   clk_r_REG9692_S1 : DFF_X1 port map( D => n2695, CK => CLK, Q => n_3343, QN 
                           => n29464);
   clk_r_REG9690_S1 : DFF_X1 port map( D => n2696, CK => CLK, Q => n_3344, QN 
                           => n29463);
   clk_r_REG9196_S1 : DFF_X1 port map( D => n2815, CK => CLK, Q => n_3345, QN 
                           => n29462);
   clk_r_REG9688_S1 : DFF_X1 port map( D => n2697, CK => CLK, Q => n_3346, QN 
                           => n29461);
   clk_r_REG8797_S1 : DFF_X1 port map( D => n2920, CK => CLK, Q => n_3347, QN 
                           => n29460);
   clk_r_REG9780_S1 : DFF_X1 port map( D => n2907, CK => CLK, Q => n_3348, QN 
                           => n29459);
   clk_r_REG9260_S1 : DFF_X1 port map( D => n2847, CK => CLK, Q => n_3349, QN 
                           => n29458);
   clk_r_REG9194_S1 : DFF_X1 port map( D => n2816, CK => CLK, Q => n_3350, QN 
                           => n29457);
   clk_r_REG9258_S1 : DFF_X1 port map( D => n2848, CK => CLK, Q => n_3351, QN 
                           => n29456);
   clk_r_REG9778_S1 : DFF_X1 port map( D => n2908, CK => CLK, Q => n_3352, QN 
                           => n29455);
   clk_r_REG8795_S1 : DFF_X1 port map( D => n2921, CK => CLK, Q => n_3353, QN 
                           => n29454);
   clk_r_REG9686_S1 : DFF_X1 port map( D => n2698, CK => CLK, Q => n_3354, QN 
                           => n29453);
   clk_r_REG8859_S1 : DFF_X1 port map( D => n2953, CK => CLK, Q => n_3355, QN 
                           => n29452);
   clk_r_REG8486_S1 : DFF_X1 port map( D => n3076, CK => CLK, Q => n_3356, QN 
                           => n29451);
   clk_r_REG9528_S1 : DFF_X1 port map( D => n2649, CK => CLK, Q => n_3357, QN 
                           => n29450);
   clk_r_REG9526_S1 : DFF_X1 port map( D => n2650, CK => CLK, Q => n_3358, QN 
                           => n29449);
   clk_r_REG8476_S1 : DFF_X1 port map( D => n3081, CK => CLK, Q => n_3359, QN 
                           => n29448);
   clk_r_REG8602_S1 : DFF_X1 port map( D => n3114, CK => CLK, Q => n_3360, QN 
                           => n29447);
   clk_r_REG8670_S1 : DFF_X1 port map( D => n3144, CK => CLK, Q => n_3361, QN 
                           => n29446);
   clk_r_REG9067_S1 : DFF_X1 port map( D => n3179, CK => CLK, Q => n_3362, QN 
                           => n29445);
   clk_r_REG9524_S1 : DFF_X1 port map( D => n2651, CK => CLK, Q => n_3363, QN 
                           => n29444);
   clk_r_REG9522_S1 : DFF_X1 port map( D => n2652, CK => CLK, Q => n_3364, QN 
                           => n29443);
   clk_r_REG9130_S1 : DFF_X1 port map( D => n3232, CK => CLK, Q => n_3365, QN 
                           => n29442);
   clk_r_REG9520_S1 : DFF_X1 port map( D => n2653, CK => CLK, Q => n_3366, QN 
                           => n29441);
   clk_r_REG8330_S1 : DFF_X1 port map( D => n3241, CK => CLK, Q => n_3367, QN 
                           => n29440);
   clk_r_REG9518_S1 : DFF_X1 port map( D => n2654, CK => CLK, Q => n_3368, QN 
                           => n29439);
   clk_r_REG7495_S1 : DFF_X1 port map( D => n3274, CK => CLK, Q => n_3369, QN 
                           => n29438);
   clk_r_REG9516_S1 : DFF_X1 port map( D => n2655, CK => CLK, Q => n_3370, QN 
                           => n29437);
   clk_r_REG9592_S1 : DFF_X1 port map( D => n2681, CK => CLK, Q => n_3371, QN 
                           => n29436);
   clk_r_REG9590_S1 : DFF_X1 port map( D => n2682, CK => CLK, Q => n_3372, QN 
                           => n29435);
   clk_r_REG9588_S1 : DFF_X1 port map( D => n2683, CK => CLK, Q => n_3373, QN 
                           => n29434);
   clk_r_REG9586_S1 : DFF_X1 port map( D => n2684, CK => CLK, Q => n_3374, QN 
                           => n29433);
   clk_r_REG9584_S1 : DFF_X1 port map( D => n2685, CK => CLK, Q => n_3375, QN 
                           => n29432);
   clk_r_REG9582_S1 : DFF_X1 port map( D => n2686, CK => CLK, Q => n_3376, QN 
                           => n29431);
   clk_r_REG9580_S1 : DFF_X1 port map( D => n2687, CK => CLK, Q => n_3377, QN 
                           => n29430);
   clk_r_REG9578_S1 : DFF_X1 port map( D => n2688, CK => CLK, Q => n_3378, QN 
                           => n29429);
   clk_r_REG9684_S1 : DFF_X1 port map( D => n2699, CK => CLK, Q => n_3379, QN 
                           => n29428);
   clk_r_REG9400_S1 : DFF_X1 port map( D => n2585, CK => CLK, Q => n_3380, QN 
                           => n29427);
   clk_r_REG9398_S1 : DFF_X1 port map( D => n2586, CK => CLK, Q => n_3381, QN 
                           => n29426);
   clk_r_REG9712_S1 : DFF_X1 port map( D => n2749, CK => CLK, Q => n_3382, QN 
                           => n29425);
   clk_r_REG9396_S1 : DFF_X1 port map( D => n2587, CK => CLK, Q => n_3383, QN 
                           => n29424);
   clk_r_REG9394_S1 : DFF_X1 port map( D => n2588, CK => CLK, Q => n_3384, QN 
                           => n29423);
   clk_r_REG9392_S1 : DFF_X1 port map( D => n2589, CK => CLK, Q => n_3385, QN 
                           => n29422);
   clk_r_REG9390_S1 : DFF_X1 port map( D => n2590, CK => CLK, Q => n_3386, QN 
                           => n29421);
   clk_r_REG9514_S1 : DFF_X1 port map( D => n2656, CK => CLK, Q => n_3387, QN 
                           => n29420);
   clk_r_REG9388_S1 : DFF_X1 port map( D => n2591, CK => CLK, Q => n_3388, QN 
                           => n29419);
   clk_r_REG9386_S1 : DFF_X1 port map( D => n2592, CK => CLK, Q => n_3389, QN 
                           => n29418);
   clk_r_REG8793_S1 : DFF_X1 port map( D => n2922, CK => CLK, Q => n_3390, QN 
                           => n29417);
   clk_r_REG8857_S1 : DFF_X1 port map( D => n2954, CK => CLK, Q => n_3391, QN 
                           => n29416);
   clk_r_REG7236_S1 : DFF_X1 port map( D => n3077, CK => CLK, Q => n_3392, QN 
                           => n29415);
   clk_r_REG9450_S1 : DFF_X1 port map( D => n2624, CK => CLK, Q => n_3393, QN 
                           => n29414);
   clk_r_REG9448_S1 : DFF_X1 port map( D => n2625, CK => CLK, Q => n_3394, QN 
                           => n29413);
   clk_r_REG9446_S1 : DFF_X1 port map( D => n2626, CK => CLK, Q => n_3395, QN 
                           => n29412);
   clk_r_REG9444_S1 : DFF_X1 port map( D => n2627, CK => CLK, Q => n_3396, QN 
                           => n29411);
   clk_r_REG9442_S1 : DFF_X1 port map( D => n2628, CK => CLK, Q => n_3397, QN 
                           => n29410);
   clk_r_REG6986_S1 : DFF_X1 port map( D => n2629, CK => CLK, Q => n_3398, QN 
                           => n29409);
   clk_r_REG8474_S1 : DFF_X1 port map( D => n3082, CK => CLK, Q => n_3399, QN 
                           => n29408);
   clk_r_REG9478_S1 : DFF_X1 port map( D => n2605, CK => CLK, Q => n_3400, QN 
                           => n29407);
   clk_r_REG9476_S1 : DFF_X1 port map( D => n2604, CK => CLK, Q => n_3401, QN 
                           => n29406);
   clk_r_REG8600_S1 : DFF_X1 port map( D => n3115, CK => CLK, Q => n_3402, QN 
                           => n29405);
   clk_r_REG8668_S1 : DFF_X1 port map( D => n3145, CK => CLK, Q => n_3403, QN 
                           => n29404);
   clk_r_REG7493_S1 : DFF_X1 port map( D => n3275, CK => CLK, Q => n_3404, QN 
                           => n29403);
   clk_r_REG8328_S1 : DFF_X1 port map( D => n3242, CK => CLK, Q => n_3405, QN 
                           => n29402);
   clk_r_REG9474_S1 : DFF_X1 port map( D => n2603, CK => CLK, Q => n_3406, QN 
                           => n29401);
   clk_r_REG9472_S1 : DFF_X1 port map( D => n2602, CK => CLK, Q => n_3407, QN 
                           => n29400);
   clk_r_REG9065_S1 : DFF_X1 port map( D => n3178, CK => CLK, Q => n_3408, QN 
                           => n29399);
   clk_r_REG8326_S1 : DFF_X1 port map( D => n3243, CK => CLK, Q => n_3409, QN 
                           => n29398);
   clk_r_REG7491_S1 : DFF_X1 port map( D => n3276, CK => CLK, Q => n_3410, QN 
                           => n29397);
   clk_r_REG9063_S1 : DFF_X1 port map( D => n3177, CK => CLK, Q => n_3411, QN 
                           => n29396);
   clk_r_REG8666_S1 : DFF_X1 port map( D => n3146, CK => CLK, Q => n_3412, QN 
                           => n29395);
   clk_r_REG8598_S1 : DFF_X1 port map( D => n3116, CK => CLK, Q => n_3413, QN 
                           => n29394);
   clk_r_REG9384_S1 : DFF_X1 port map( D => n2593, CK => CLK, Q => n_3414, QN 
                           => n29393);
   clk_r_REG9470_S1 : DFF_X1 port map( D => n2601, CK => CLK, Q => n_3415, QN 
                           => n29392);
   clk_r_REG9512_S1 : DFF_X1 port map( D => n2657, CK => CLK, Q => n_3416, QN 
                           => n29391);
   clk_r_REG9576_S1 : DFF_X1 port map( D => n2689, CK => CLK, Q => n_3417, QN 
                           => n29390);
   clk_r_REG9682_S1 : DFF_X1 port map( D => n2700, CK => CLK, Q => n_3418, QN 
                           => n29389);
   clk_r_REG8472_S1 : DFF_X1 port map( D => n3083, CK => CLK, Q => n_3419, QN 
                           => n29388);
   clk_r_REG8544_S1 : DFF_X1 port map( D => n3047, CK => CLK, Q => n_3420, QN 
                           => n29387);
   clk_r_REG8855_S1 : DFF_X1 port map( D => n2955, CK => CLK, Q => n_3421, QN 
                           => n29386);
   clk_r_REG8791_S1 : DFF_X1 port map( D => n2923, CK => CLK, Q => n_3422, QN 
                           => n29385);
   clk_r_REG9776_S1 : DFF_X1 port map( D => n2909, CK => CLK, Q => n_3423, QN 
                           => n29384);
   clk_r_REG9256_S1 : DFF_X1 port map( D => n2849, CK => CLK, Q => n_3424, QN 
                           => n29383);
   clk_r_REG9320_S1 : DFF_X1 port map( D => n2560, CK => CLK, Q => n_3425, QN 
                           => n29382);
   clk_r_REG9318_S1 : DFF_X1 port map( D => n2561, CK => CLK, Q => n_3426, QN 
                           => n29381);
   clk_r_REG9316_S1 : DFF_X1 port map( D => n2562, CK => CLK, Q => n_3427, QN 
                           => n29380);
   clk_r_REG9192_S1 : DFF_X1 port map( D => n2817, CK => CLK, Q => n_3428, QN 
                           => n29379);
   clk_r_REG9680_S1 : DFF_X1 port map( D => n2701, CK => CLK, Q => n_3429, QN 
                           => n29378);
   clk_r_REG9314_S1 : DFF_X1 port map( D => n2563, CK => CLK, Q => n_3430, QN 
                           => n29377);
   clk_r_REG9312_S1 : DFF_X1 port map( D => n2564, CK => CLK, Q => n_3431, QN 
                           => n29376);
   clk_r_REG7004_S1 : DFF_X1 port map( D => n2565, CK => CLK, Q => n_3432, QN 
                           => n29375);
   clk_r_REG9370_S1 : DFF_X1 port map( D => n2535, CK => CLK, Q => n_3433, QN 
                           => n29374);
   clk_r_REG9368_S1 : DFF_X1 port map( D => n2536, CK => CLK, Q => n_3434, QN 
                           => n29373);
   clk_r_REG9366_S1 : DFF_X1 port map( D => n2537, CK => CLK, Q => n_3435, QN 
                           => n29372);
   clk_r_REG9364_S1 : DFF_X1 port map( D => n2538, CK => CLK, Q => n_3436, QN 
                           => n29371);
   clk_r_REG9362_S1 : DFF_X1 port map( D => n2539, CK => CLK, Q => n_3437, QN 
                           => n29370);
   clk_r_REG9360_S1 : DFF_X1 port map( D => n2540, CK => CLK, Q => n_3438, QN 
                           => n29369);
   clk_r_REG9574_S1 : DFF_X1 port map( D => n2690, CK => CLK, Q => n_3439, QN 
                           => n29368);
   clk_r_REG9510_S1 : DFF_X1 port map( D => n2658, CK => CLK, Q => n_3440, QN 
                           => n29367);
   clk_r_REG9468_S1 : DFF_X1 port map( D => n2600, CK => CLK, Q => n_3441, QN 
                           => n29366);
   clk_r_REG9382_S1 : DFF_X1 port map( D => n2594, CK => CLK, Q => n_3442, QN 
                           => n29365);
   clk_r_REG9358_S1 : DFF_X1 port map( D => n2541, CK => CLK, Q => n_3443, QN 
                           => n29364);
   clk_r_REG8789_S1 : DFF_X1 port map( D => n2924, CK => CLK, Q => n_3444, QN 
                           => n29363);
   clk_r_REG8853_S1 : DFF_X1 port map( D => n2956, CK => CLK, Q => n_3445, QN 
                           => n29362);
   clk_r_REG8542_S1 : DFF_X1 port map( D => n3048, CK => CLK, Q => n_3446, QN 
                           => n29361);
   clk_r_REG8470_S1 : DFF_X1 port map( D => n3084, CK => CLK, Q => n_3447, QN 
                           => n29360);
   clk_r_REG8596_S1 : DFF_X1 port map( D => n3117, CK => CLK, Q => n_3448, QN 
                           => n29359);
   clk_r_REG8664_S1 : DFF_X1 port map( D => n3147, CK => CLK, Q => n_3449, QN 
                           => n29358);
   clk_r_REG9061_S1 : DFF_X1 port map( D => n3176, CK => CLK, Q => n_3450, QN 
                           => n29357);
   clk_r_REG7489_S1 : DFF_X1 port map( D => n3277, CK => CLK, Q => n_3451, QN 
                           => n29356);
   clk_r_REG8324_S1 : DFF_X1 port map( D => n3244, CK => CLK, Q => n_3452, QN 
                           => n29355);
   clk_r_REG9128_S1 : DFF_X1 port map( D => n3233, CK => CLK, Q => n_3453, QN 
                           => n29354);
   clk_r_REG9710_S1 : DFF_X1 port map( D => n2750, CK => CLK, Q => n_3454, QN 
                           => n29353);
   clk_r_REG9708_S1 : DFF_X1 port map( D => n2751, CK => CLK, Q => n_3455, QN 
                           => n29352);
   clk_r_REG9706_S1 : DFF_X1 port map( D => n2752, CK => CLK, Q => n_3456, QN 
                           => n29351);
   clk_r_REG8685_S1 : DFF_X1 port map( D => n2880, CK => CLK, Q => n_3457, QN 
                           => n29350);
   clk_r_REG8683_S1 : DFF_X1 port map( D => n2881, CK => CLK, Q => n_3458, QN 
                           => n29349);
   clk_r_REG8681_S1 : DFF_X1 port map( D => n2882, CK => CLK, Q => n_3459, QN 
                           => n29348);
   clk_r_REG8679_S1 : DFF_X1 port map( D => n2883, CK => CLK, Q => n_3460, QN 
                           => n29347);
   clk_r_REG8677_S1 : DFF_X1 port map( D => n2884, CK => CLK, Q => n_3461, QN 
                           => n29346);
   clk_r_REG7145_S1 : DFF_X1 port map( D => n2885, CK => CLK, Q => n_3462, QN 
                           => n29345);
   clk_r_REG9190_S1 : DFF_X1 port map( D => n2818, CK => CLK, Q => n_3463, QN 
                           => n29344);
   clk_r_REG9254_S1 : DFF_X1 port map( D => n2850, CK => CLK, Q => n_3464, QN 
                           => n29343);
   clk_r_REG9774_S1 : DFF_X1 port map( D => n2910, CK => CLK, Q => n_3465, QN 
                           => n29342);
   clk_r_REG8787_S1 : DFF_X1 port map( D => n2925, CK => CLK, Q => n_3466, QN 
                           => n29341);
   clk_r_REG8735_S1 : DFF_X1 port map( D => n2855, CK => CLK, Q => n_3467, QN 
                           => n29340);
   clk_r_REG8733_S1 : DFF_X1 port map( D => n2856, CK => CLK, Q => n_3468, QN 
                           => n29339);
   clk_r_REG8731_S1 : DFF_X1 port map( D => n2857, CK => CLK, Q => n_3469, QN 
                           => n29338);
   clk_r_REG8729_S1 : DFF_X1 port map( D => n2858, CK => CLK, Q => n_3470, QN 
                           => n29337);
   clk_r_REG8727_S1 : DFF_X1 port map( D => n2859, CK => CLK, Q => n_3471, QN 
                           => n29336);
   clk_r_REG8725_S1 : DFF_X1 port map( D => n2860, CK => CLK, Q => n_3472, QN 
                           => n29335);
   clk_r_REG8723_S1 : DFF_X1 port map( D => n2861, CK => CLK, Q => n_3473, QN 
                           => n29334);
   clk_r_REG8851_S1 : DFF_X1 port map( D => n2957, CK => CLK, Q => n_3474, QN 
                           => n29333);
   clk_r_REG8540_S1 : DFF_X1 port map( D => n3049, CK => CLK, Q => n_3475, QN 
                           => n29332);
   clk_r_REG8468_S1 : DFF_X1 port map( D => n3085, CK => CLK, Q => n_3476, QN 
                           => n29331);
   clk_r_REG9704_S1 : DFF_X1 port map( D => n2753, CK => CLK, Q => n_3477, QN 
                           => n29330);
   clk_r_REG8594_S1 : DFF_X1 port map( D => n3118, CK => CLK, Q => n_3478, QN 
                           => n29329);
   clk_r_REG8662_S1 : DFF_X1 port map( D => n3148, CK => CLK, Q => n_3479, QN 
                           => n29328);
   clk_r_REG9059_S1 : DFF_X1 port map( D => n3175, CK => CLK, Q => n_3480, QN 
                           => n29327);
   clk_r_REG9126_S1 : DFF_X1 port map( D => n3234, CK => CLK, Q => n_3481, QN 
                           => n29326);
   clk_r_REG8885_S1 : DFF_X1 port map( D => n3004, CK => CLK, Q => n_3482, QN 
                           => n29325);
   clk_r_REG7064_S1 : DFF_X1 port map( D => n3174, CK => CLK, Q => n_3483, QN 
                           => n29324);
   clk_r_REG8883_S1 : DFF_X1 port map( D => n3005, CK => CLK, Q => n_3484, QN 
                           => n29323);
   clk_r_REG8881_S1 : DFF_X1 port map( D => n3006, CK => CLK, Q => n_3485, QN 
                           => n29322);
   clk_r_REG8879_S1 : DFF_X1 port map( D => n3007, CK => CLK, Q => n_3486, QN 
                           => n29321);
   clk_r_REG8877_S1 : DFF_X1 port map( D => n3008, CK => CLK, Q => n_3487, QN 
                           => n29320);
   clk_r_REG8875_S1 : DFF_X1 port map( D => n3009, CK => CLK, Q => n_3488, QN 
                           => n29319);
   clk_r_REG8873_S1 : DFF_X1 port map( D => n3010, CK => CLK, Q => n_3489, QN 
                           => n29318);
   clk_r_REG8322_S1 : DFF_X1 port map( D => n3245, CK => CLK, Q => n_3490, QN 
                           => n29317);
   clk_r_REG7487_S1 : DFF_X1 port map( D => n3278, CK => CLK, Q => n_3491, QN 
                           => n29316);
   clk_r_REG8871_S1 : DFF_X1 port map( D => n3011, CK => CLK, Q => n_3492, QN 
                           => n29315);
   clk_r_REG8869_S1 : DFF_X1 port map( D => n3012, CK => CLK, Q => n_3493, QN 
                           => n29314);
   clk_r_REG7124_S1 : DFF_X1 port map( D => n3013, CK => CLK, Q => n_3494, QN 
                           => n29313);
   clk_r_REG8927_S1 : DFF_X1 port map( D => n2983, CK => CLK, Q => n_3495, QN 
                           => n29312);
   clk_r_REG8925_S1 : DFF_X1 port map( D => n2984, CK => CLK, Q => n_3496, QN 
                           => n29311);
   clk_r_REG8923_S1 : DFF_X1 port map( D => n2985, CK => CLK, Q => n_3497, QN 
                           => n29310);
   clk_r_REG9356_S1 : DFF_X1 port map( D => n2542, CK => CLK, Q => n_3498, QN 
                           => n29309);
   clk_r_REG9380_S1 : DFF_X1 port map( D => n2595, CK => CLK, Q => n_3499, QN 
                           => n29308);
   clk_r_REG9466_S1 : DFF_X1 port map( D => n2599, CK => CLK, Q => n_3500, QN 
                           => n29307);
   clk_r_REG9001_S1 : DFF_X1 port map( D => n2785, CK => CLK, Q => n_3501, QN 
                           => n29306);
   clk_r_REG8999_S1 : DFF_X1 port map( D => n2786, CK => CLK, Q => n_3502, QN 
                           => n29305);
   clk_r_REG8997_S1 : DFF_X1 port map( D => n2787, CK => CLK, Q => n_3503, QN 
                           => n29304);
   clk_r_REG8995_S1 : DFF_X1 port map( D => n2788, CK => CLK, Q => n_3504, QN 
                           => n29303);
   clk_r_REG7105_S1 : DFF_X1 port map( D => n2789, CK => CLK, Q => n_3505, QN 
                           => n29302);
   clk_r_REG9053_S1 : DFF_X1 port map( D => n2759, CK => CLK, Q => n_3506, QN 
                           => n29301);
   clk_r_REG9508_S1 : DFF_X1 port map( D => n2659, CK => CLK, Q => n_3507, QN 
                           => n29300);
   clk_r_REG9572_S1 : DFF_X1 port map( D => n2691, CK => CLK, Q => n_3508, QN 
                           => n29299);
   clk_r_REG9678_S1 : DFF_X1 port map( D => n2702, CK => CLK, Q => n_3509, QN 
                           => n29298);
   clk_r_REG9702_S1 : DFF_X1 port map( D => n2754, CK => CLK, Q => n_3510, QN 
                           => n29297);
   clk_r_REG9051_S1 : DFF_X1 port map( D => n2760, CK => CLK, Q => n_3511, QN 
                           => n29296);
   clk_r_REG8991_S1 : DFF_X1 port map( D => n3015, CK => CLK, Q => n_3512, QN 
                           => n29295);
   clk_r_REG8939_S1 : DFF_X1 port map( D => n3041, CK => CLK, Q => n_3513, QN 
                           => n29294);
   clk_r_REG8937_S1 : DFF_X1 port map( D => n3042, CK => CLK, Q => n_3514, QN 
                           => n29293);
   clk_r_REG8935_S1 : DFF_X1 port map( D => n3043, CK => CLK, Q => n_3515, QN 
                           => n29292);
   clk_r_REG8933_S1 : DFF_X1 port map( D => n3044, CK => CLK, Q => n_3516, QN 
                           => n29291);
   clk_r_REG7117_S1 : DFF_X1 port map( D => n3045, CK => CLK, Q => n_3517, QN 
                           => n29290);
   clk_r_REG8989_S1 : DFF_X1 port map( D => n3016, CK => CLK, Q => n_3518, QN 
                           => n29289);
   clk_r_REG9049_S1 : DFF_X1 port map( D => n2761, CK => CLK, Q => n_3519, QN 
                           => n29288);
   clk_r_REG9047_S1 : DFF_X1 port map( D => n2762, CK => CLK, Q => n_3520, QN 
                           => n29287);
   clk_r_REG9045_S1 : DFF_X1 port map( D => n2763, CK => CLK, Q => n_3521, QN 
                           => n29286);
   clk_r_REG8987_S1 : DFF_X1 port map( D => n3017, CK => CLK, Q => n_3522, QN 
                           => n29285);
   clk_r_REG9043_S1 : DFF_X1 port map( D => n2764, CK => CLK, Q => n_3523, QN 
                           => n29284);
   clk_r_REG9041_S1 : DFF_X1 port map( D => n2765, CK => CLK, Q => n_3524, QN 
                           => n29283);
   clk_r_REG8921_S1 : DFF_X1 port map( D => n2986, CK => CLK, Q => n_3525, QN 
                           => n29282);
   clk_r_REG9464_S1 : DFF_X1 port map( D => n2598, CK => CLK, Q => n_3526, QN 
                           => n29281);
   clk_r_REG8985_S1 : DFF_X1 port map( D => n3018, CK => CLK, Q => n_3527, QN 
                           => n29280);
   clk_r_REG8983_S1 : DFF_X1 port map( D => n3019, CK => CLK, Q => n_3528, QN 
                           => n29279);
   clk_r_REG9700_S1 : DFF_X1 port map( D => n2755, CK => CLK, Q => n_3529, QN 
                           => n29278);
   clk_r_REG8981_S1 : DFF_X1 port map( D => n3020, CK => CLK, Q => n_3530, QN 
                           => n29277);
   clk_r_REG9039_S1 : DFF_X1 port map( D => n2766, CK => CLK, Q => n_3531, QN 
                           => n29276);
   clk_r_REG9188_S1 : DFF_X1 port map( D => n2819, CK => CLK, Q => n_3532, QN 
                           => n29275);
   clk_r_REG9252_S1 : DFF_X1 port map( D => n2851, CK => CLK, Q => n_3533, QN 
                           => n29274);
   clk_r_REG8721_S1 : DFF_X1 port map( D => n2862, CK => CLK, Q => n_3534, QN 
                           => n29273);
   clk_r_REG9772_S1 : DFF_X1 port map( D => n2911, CK => CLK, Q => n_3535, QN 
                           => n29272);
   clk_r_REG8785_S1 : DFF_X1 port map( D => n2926, CK => CLK, Q => n_3536, QN 
                           => n29271);
   clk_r_REG8849_S1 : DFF_X1 port map( D => n2958, CK => CLK, Q => n_3537, QN 
                           => n29270);
   clk_r_REG8538_S1 : DFF_X1 port map( D => n3050, CK => CLK, Q => n_3538, QN 
                           => n29269);
   clk_r_REG8979_S1 : DFF_X1 port map( D => n3021, CK => CLK, Q => n_3539, QN 
                           => n29268);
   clk_r_REG8592_S1 : DFF_X1 port map( D => n3119, CK => CLK, Q => n_3540, QN 
                           => n29267);
   clk_r_REG8466_S1 : DFF_X1 port map( D => n3086, CK => CLK, Q => n_3541, QN 
                           => n29266);
   clk_r_REG8977_S1 : DFF_X1 port map( D => n3022, CK => CLK, Q => n_3542, QN 
                           => n29265);
   clk_r_REG8975_S1 : DFF_X1 port map( D => n3023, CK => CLK, Q => n_3543, QN 
                           => n29264);
   clk_r_REG8660_S1 : DFF_X1 port map( D => n3149, CK => CLK, Q => n_3544, QN 
                           => n29263);
   clk_r_REG9934_S1 : DFF_X1 port map( D => n3548, CK => CLK, Q => n_3545, QN 
                           => n29262);
   clk_r_REG9932_S1 : DFF_X1 port map( D => n3549, CK => CLK, Q => n_3546, QN 
                           => n29261);
   clk_r_REG9930_S1 : DFF_X1 port map( D => n3550, CK => CLK, Q => n_3547, QN 
                           => n29260);
   clk_r_REG9124_S1 : DFF_X1 port map( D => n3235, CK => CLK, Q => n_3548, QN 
                           => n29259);
   clk_r_REG9122_S1 : DFF_X1 port map( D => n3236, CK => CLK, Q => n_3549, QN 
                           => n29258);
   clk_r_REG7045_S1 : DFF_X1 port map( D => n3237, CK => CLK, Q => n_3550, QN 
                           => n29257);
   clk_r_REG9180_S1 : DFF_X1 port map( D => n3207, CK => CLK, Q => n_3551, QN 
                           => n29256);
   clk_r_REG9178_S1 : DFF_X1 port map( D => n3208, CK => CLK, Q => n_3552, QN 
                           => n29255);
   clk_r_REG9176_S1 : DFF_X1 port map( D => n3209, CK => CLK, Q => n_3553, QN 
                           => n29254);
   clk_r_REG9174_S1 : DFF_X1 port map( D => n3210, CK => CLK, Q => n_3554, QN 
                           => n29253);
   clk_r_REG9172_S1 : DFF_X1 port map( D => n3211, CK => CLK, Q => n_3555, QN 
                           => n29252);
   clk_r_REG9170_S1 : DFF_X1 port map( D => n3212, CK => CLK, Q => n_3556, QN 
                           => n29251);
   clk_r_REG9168_S1 : DFF_X1 port map( D => n3213, CK => CLK, Q => n_3557, QN 
                           => n29250);
   clk_r_REG9166_S1 : DFF_X1 port map( D => n3214, CK => CLK, Q => n_3558, QN 
                           => n29249);
   clk_r_REG9928_S1 : DFF_X1 port map( D => n3551, CK => CLK, Q => n_3559, QN 
                           => n29248);
   clk_r_REG7599_S1 : DFF_X1 port map( D => n3316, CK => CLK, Q => n_3560, QN 
                           => n29247);
   clk_r_REG7597_S1 : DFF_X1 port map( D => n3317, CK => CLK, Q => n_3561, QN 
                           => n29246);
   clk_r_REG7595_S1 : DFF_X1 port map( D => n3318, CK => CLK, Q => n_3562, QN 
                           => n29245);
   clk_r_REG7593_S1 : DFF_X1 port map( D => n3319, CK => CLK, Q => n_3563, QN 
                           => n29244);
   clk_r_REG9770_S1 : DFF_X1 port map( D => n2912, CK => CLK, Q => n_3564, QN 
                           => n29243);
   clk_r_REG9768_S1 : DFF_X1 port map( D => n2913, CK => CLK, Q => n_3565, QN 
                           => n29242);
   clk_r_REG9766_S1 : DFF_X1 port map( D => n2914, CK => CLK, Q => n_3566, QN 
                           => n29241);
   clk_r_REG9764_S1 : DFF_X1 port map( D => n2915, CK => CLK, Q => n_3567, QN 
                           => n29240);
   clk_r_REG7591_S1 : DFF_X1 port map( D => n3320, CK => CLK, Q => n_3568, QN 
                           => n29239);
   clk_r_REG9762_S1 : DFF_X1 port map( D => n2916, CK => CLK, Q => n_3569, QN 
                           => n29238);
   clk_r_REG7589_S1 : DFF_X1 port map( D => n3321, CK => CLK, Q => n_3570, QN 
                           => n29237);
   clk_r_REG7587_S1 : DFF_X1 port map( D => n3322, CK => CLK, Q => n_3571, QN 
                           => n29236);
   clk_r_REG6950_S1 : DFF_X1 port map( D => n2917, CK => CLK, Q => n_3572, QN 
                           => n29235);
   clk_r_REG9822_S1 : DFF_X1 port map( D => n2886, CK => CLK, Q => n_3573, QN 
                           => n29234);
   clk_r_REG7585_S1 : DFF_X1 port map( D => n3323, CK => CLK, Q => n_3574, QN 
                           => n29233);
   clk_r_REG9820_S1 : DFF_X1 port map( D => n2887, CK => CLK, Q => n_3575, QN 
                           => n29232);
   clk_r_REG9186_S1 : DFF_X1 port map( D => n2820, CK => CLK, Q => n_3576, QN 
                           => n29231);
   clk_r_REG7026_S1 : DFF_X1 port map( D => n2821, CK => CLK, Q => n_3577, QN 
                           => n29230);
   clk_r_REG9250_S1 : DFF_X1 port map( D => n2852, CK => CLK, Q => n_3578, QN 
                           => n29229);
   clk_r_REG9246_S1 : DFF_X1 port map( D => n2790, CK => CLK, Q => n_3579, QN 
                           => n29228);
   clk_r_REG7018_S1 : DFF_X1 port map( D => n2853, CK => CLK, Q => n_3580, QN 
                           => n29227);
   clk_r_REG9244_S1 : DFF_X1 port map( D => n2791, CK => CLK, Q => n_3581, QN 
                           => n29226);
   clk_r_REG9242_S1 : DFF_X1 port map( D => n2792, CK => CLK, Q => n_3582, QN 
                           => n29225);
   clk_r_REG9310_S1 : DFF_X1 port map( D => n2822, CK => CLK, Q => n_3583, QN 
                           => n29224);
   clk_r_REG9698_S1 : DFF_X1 port map( D => n2756, CK => CLK, Q => n_3584, QN 
                           => n29223);
   clk_r_REG9308_S1 : DFF_X1 port map( D => n2823, CK => CLK, Q => n_3585, QN 
                           => n29222);
   clk_r_REG9240_S1 : DFF_X1 port map( D => n2793, CK => CLK, Q => n_3586, QN 
                           => n29221);
   clk_r_REG9306_S1 : DFF_X1 port map( D => n2824, CK => CLK, Q => n_3587, QN 
                           => n29220);
   clk_r_REG9304_S1 : DFF_X1 port map( D => n2825, CK => CLK, Q => n_3588, QN 
                           => n29219);
   clk_r_REG9302_S1 : DFF_X1 port map( D => n2826, CK => CLK, Q => n_3589, QN 
                           => n29218);
   clk_r_REG9300_S1 : DFF_X1 port map( D => n2827, CK => CLK, Q => n_3590, QN 
                           => n29217);
   clk_r_REG9298_S1 : DFF_X1 port map( D => n2828, CK => CLK, Q => n_3591, QN 
                           => n29216);
   clk_r_REG9926_S1 : DFF_X1 port map( D => n3552, CK => CLK, Q => n_3592, QN 
                           => n29215);
   clk_r_REG9296_S1 : DFF_X1 port map( D => n2829, CK => CLK, Q => n_3593, QN 
                           => n29214);
   clk_r_REG6957_S1 : DFF_X1 port map( D => n2757, CK => CLK, Q => n_3594, QN 
                           => n29213);
   clk_r_REG9238_S1 : DFF_X1 port map( D => n2794, CK => CLK, Q => n_3595, QN 
                           => n29212);
   clk_r_REG9818_S1 : DFF_X1 port map( D => n2888, CK => CLK, Q => n_3596, QN 
                           => n29211);
   clk_r_REG9924_S1 : DFF_X1 port map( D => n3553, CK => CLK, Q => n_3597, QN 
                           => n29210);
   clk_r_REG9378_S1 : DFF_X1 port map( D => n2596, CK => CLK, Q => n_3598, QN 
                           => n29209);
   clk_r_REG9236_S1 : DFF_X1 port map( D => n2795, CK => CLK, Q => n_3599, QN 
                           => n29208);
   clk_r_REG9234_S1 : DFF_X1 port map( D => n2796, CK => CLK, Q => n_3600, QN 
                           => n29207);
   clk_r_REG6995_S1 : DFF_X1 port map( D => n2597, CK => CLK, Q => n_3601, QN 
                           => n29206);
   clk_r_REG9438_S1 : DFF_X1 port map( D => n2566, CK => CLK, Q => n_3602, QN 
                           => n29205);
   clk_r_REG9436_S1 : DFF_X1 port map( D => n2567, CK => CLK, Q => n_3603, QN 
                           => n29204);
   clk_r_REG9434_S1 : DFF_X1 port map( D => n2568, CK => CLK, Q => n_3604, QN 
                           => n29203);
   clk_r_REG9432_S1 : DFF_X1 port map( D => n2569, CK => CLK, Q => n_3605, QN 
                           => n29202);
   clk_r_REG9922_S1 : DFF_X1 port map( D => n3554, CK => CLK, Q => n_3606, QN 
                           => n29201);
   clk_r_REG9506_S1 : DFF_X1 port map( D => n2660, CK => CLK, Q => n_3607, QN 
                           => n29200);
   clk_r_REG9430_S1 : DFF_X1 port map( D => n2570, CK => CLK, Q => n_3608, QN 
                           => n29199);
   clk_r_REG6979_S1 : DFF_X1 port map( D => n2661, CK => CLK, Q => n_3609, QN 
                           => n29198);
   clk_r_REG9566_S1 : DFF_X1 port map( D => n2630, CK => CLK, Q => n_3610, QN 
                           => n29197);
   clk_r_REG9564_S1 : DFF_X1 port map( D => n2631, CK => CLK, Q => n_3611, QN 
                           => n29196);
   clk_r_REG9232_S1 : DFF_X1 port map( D => n2797, CK => CLK, Q => n_3612, QN 
                           => n29195);
   clk_r_REG9428_S1 : DFF_X1 port map( D => n2571, CK => CLK, Q => n_3613, QN 
                           => n29194);
   clk_r_REG9570_S1 : DFF_X1 port map( D => n2692, CK => CLK, Q => n_3614, QN 
                           => n29193);
   clk_r_REG9756_S1 : DFF_X1 port map( D => n2727, CK => CLK, Q => n_3615, QN 
                           => n29192);
   clk_r_REG9562_S1 : DFF_X1 port map( D => n2632, CK => CLK, Q => n_3616, QN 
                           => n29191);
   clk_r_REG9560_S1 : DFF_X1 port map( D => n2633, CK => CLK, Q => n_3617, QN 
                           => n29190);
   clk_r_REG9426_S1 : DFF_X1 port map( D => n2572, CK => CLK, Q => n_3618, QN 
                           => n29189);
   clk_r_REG6972_S1 : DFF_X1 port map( D => n2693, CK => CLK, Q => n_3619, QN 
                           => n29188);
   clk_r_REG9630_S1 : DFF_X1 port map( D => n2662, CK => CLK, Q => n_3620, QN 
                           => n29187);
   clk_r_REG9558_S1 : DFF_X1 port map( D => n2634, CK => CLK, Q => n_3621, QN 
                           => n29186);
   clk_r_REG9556_S1 : DFF_X1 port map( D => n2635, CK => CLK, Q => n_3622, QN 
                           => n29185);
   clk_r_REG9554_S1 : DFF_X1 port map( D => n2636, CK => CLK, Q => n_3623, QN 
                           => n29184);
   clk_r_REG9552_S1 : DFF_X1 port map( D => n2637, CK => CLK, Q => n_3624, QN 
                           => n29183);
   clk_r_REG9628_S1 : DFF_X1 port map( D => n2663, CK => CLK, Q => n_3625, QN 
                           => n29182);
   clk_r_REG9626_S1 : DFF_X1 port map( D => n2664, CK => CLK, Q => n_3626, QN 
                           => n29181);
   clk_r_REG9624_S1 : DFF_X1 port map( D => n2665, CK => CLK, Q => n_3627, QN 
                           => n29180);
   clk_r_REG9424_S1 : DFF_X1 port map( D => n2573, CK => CLK, Q => n_3628, QN 
                           => n29179);
   clk_r_REG9622_S1 : DFF_X1 port map( D => n2666, CK => CLK, Q => n_3629, QN 
                           => n29178);
   clk_r_REG9620_S1 : DFF_X1 port map( D => n2667, CK => CLK, Q => n_3630, QN 
                           => n29177);
   clk_r_REG9754_S1 : DFF_X1 port map( D => n2728, CK => CLK, Q => n_3631, QN 
                           => n29176);
   clk_r_REG9618_S1 : DFF_X1 port map( D => n2668, CK => CLK, Q => n_3632, QN 
                           => n29175);
   clk_r_REG9752_S1 : DFF_X1 port map( D => n2729, CK => CLK, Q => n_3633, QN 
                           => n29174);
   clk_r_REG9750_S1 : DFF_X1 port map( D => n2730, CK => CLK, Q => n_3634, QN 
                           => n29173);
   clk_r_REG9816_S1 : DFF_X1 port map( D => n2889, CK => CLK, Q => n_3635, QN 
                           => n29172);
   clk_r_REG9748_S1 : DFF_X1 port map( D => n2731, CK => CLK, Q => n_3636, QN 
                           => n29171);
   clk_r_REG9746_S1 : DFF_X1 port map( D => n2732, CK => CLK, Q => n_3637, QN 
                           => n29170);
   clk_r_REG9744_S1 : DFF_X1 port map( D => n2733, CK => CLK, Q => n_3638, QN 
                           => n29169);
   clk_r_REG9742_S1 : DFF_X1 port map( D => n2734, CK => CLK, Q => n_3639, QN 
                           => n29168);
   clk_r_REG9616_S1 : DFF_X1 port map( D => n2669, CK => CLK, Q => n_3640, QN 
                           => n29167);
   clk_r_REG8230_S1 : DFF_X1 port map( D => n3484, CK => CLK, Q => n_3641, QN 
                           => n29166);
   clk_r_REG8228_S1 : DFF_X1 port map( D => n3485, CK => CLK, Q => n_3642, QN 
                           => n29165);
   clk_r_REG9814_S1 : DFF_X1 port map( D => n2890, CK => CLK, Q => n_3643, QN 
                           => n29164);
   clk_r_REG8919_S1 : DFF_X1 port map( D => n2987, CK => CLK, Q => n_3644, QN 
                           => n29163);
   clk_r_REG8536_S1 : DFF_X1 port map( D => n3051, CK => CLK, Q => n_3645, QN 
                           => n29162);
   clk_r_REG9812_S1 : DFF_X1 port map( D => n2891, CK => CLK, Q => n_3646, QN 
                           => n29161);
   clk_r_REG8917_S1 : DFF_X1 port map( D => n2988, CK => CLK, Q => n_3647, QN 
                           => n29160);
   clk_r_REG8226_S1 : DFF_X1 port map( D => n3486, CK => CLK, Q => n_3648, QN 
                           => n29159);
   clk_r_REG9845_S1 : DFF_X1 port map( D => n3452, CK => CLK, Q => n_3649, QN 
                           => n29158);
   clk_r_REG9810_S1 : DFF_X1 port map( D => n2892, CK => CLK, Q => n_3650, QN 
                           => n29157);
   clk_r_REG7675_S1 : DFF_X1 port map( D => n3356, CK => CLK, Q => n_3651, QN 
                           => n29156);
   clk_r_REG7583_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n_3652, QN 
                           => n29155);
   clk_r_REG9843_S1 : DFF_X1 port map( D => n3453, CK => CLK, Q => n_3653, QN 
                           => n29154);
   clk_r_REG7889_S1 : DFF_X1 port map( D => n3420, CK => CLK, Q => n_3654, QN 
                           => n29153);
   clk_r_REG7581_S1 : DFF_X1 port map( D => n3325, CK => CLK, Q => n_3655, QN 
                           => n29152);
   clk_r_REG7971_S1 : DFF_X1 port map( D => n3388, CK => CLK, Q => n_3656, QN 
                           => n29151);
   clk_r_REG7579_S1 : DFF_X1 port map( D => n3326, CK => CLK, Q => n_3657, QN 
                           => n29150);
   clk_r_REG8370_S1 : DFF_X1 port map( D => n3516, CK => CLK, Q => n_3658, QN 
                           => n29149);
   clk_r_REG8534_S1 : DFF_X1 port map( D => n3052, CK => CLK, Q => n_3659, QN 
                           => n29148);
   clk_r_REG9841_S1 : DFF_X1 port map( D => n3454, CK => CLK, Q => n_3660, QN 
                           => n29147);
   clk_r_REG8532_S1 : DFF_X1 port map( D => n3053, CK => CLK, Q => n_3661, QN 
                           => n29146);
   clk_r_REG8915_S1 : DFF_X1 port map( D => n2989, CK => CLK, Q => n_3662, QN 
                           => n29145);
   clk_r_REG7887_S1 : DFF_X1 port map( D => n3421, CK => CLK, Q => n_3663, QN 
                           => n29144);
   clk_r_REG8368_S1 : DFF_X1 port map( D => n3517, CK => CLK, Q => n_3664, QN 
                           => n29143);
   clk_r_REG7885_S1 : DFF_X1 port map( D => n3422, CK => CLK, Q => n_3665, QN 
                           => n29142);
   clk_r_REG7673_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n_3666, QN 
                           => n29141);
   clk_r_REG7671_S1 : DFF_X1 port map( D => n3358, CK => CLK, Q => n_3667, QN 
                           => n29140);
   clk_r_REG8366_S1 : DFF_X1 port map( D => n3518, CK => CLK, Q => n_3668, QN 
                           => n29139);
   clk_r_REG7969_S1 : DFF_X1 port map( D => n3389, CK => CLK, Q => n_3669, QN 
                           => n29138);
   clk_r_REG7967_S1 : DFF_X1 port map( D => n3390, CK => CLK, Q => n_3670, QN 
                           => n29137);
   clk_r_REG9920_S1 : DFF_X1 port map( D => n3555, CK => CLK, Q => n_3671, QN 
                           => n29136);
   clk_r_REG9918_S1 : DFF_X1 port map( D => n3556, CK => CLK, Q => n_3672, QN 
                           => n29135);
   clk_r_REG6922_S1 : DFF_X1 port map( D => n3557, CK => CLK, Q => n_3673, QN 
                           => n29134);
   clk_r_REG9976_S1 : DFF_X1 port map( D => n3527, CK => CLK, Q => n_3674, QN 
                           => n29133);
   clk_r_REG9974_S1 : DFF_X1 port map( D => n3528, CK => CLK, Q => n_3675, QN 
                           => n29132);
   clk_r_REG9972_S1 : DFF_X1 port map( D => n3529, CK => CLK, Q => n_3676, QN 
                           => n29131);
   clk_r_REG9970_S1 : DFF_X1 port map( D => n3530, CK => CLK, Q => n_3677, QN 
                           => n29130);
   clk_r_REG9968_S1 : DFF_X1 port map( D => n3531, CK => CLK, Q => n_3678, QN 
                           => n29129);
   clk_r_REG9966_S1 : DFF_X1 port map( D => n3532, CK => CLK, Q => n_3679, QN 
                           => n29128);
   clk_r_REG9964_S1 : DFF_X1 port map( D => n3533, CK => CLK, Q => n_3680, QN 
                           => n29127);
   clk_r_REG9962_S1 : DFF_X1 port map( D => n3534, CK => CLK, Q => n_3681, QN 
                           => n29126);
   clk_r_REG9839_S1 : DFF_X1 port map( D => n3455, CK => CLK, Q => n_3682, QN 
                           => n29125);
   clk_r_REG7577_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n_3683, QN 
                           => n29124);
   clk_r_REG8224_S1 : DFF_X1 port map( D => n3487, CK => CLK, Q => n_3684, QN 
                           => n29123);
   clk_r_REG8530_S1 : DFF_X1 port map( D => n3054, CK => CLK, Q => n_3685, QN 
                           => n29122);
   clk_r_REG7965_S1 : DFF_X1 port map( D => n3391, CK => CLK, Q => n_3686, QN 
                           => n29121);
   clk_r_REG7669_S1 : DFF_X1 port map( D => n3359, CK => CLK, Q => n_3687, QN 
                           => n29120);
   clk_r_REG9808_S1 : DFF_X1 port map( D => n2893, CK => CLK, Q => n_3688, QN 
                           => n29119);
   clk_r_REG8913_S1 : DFF_X1 port map( D => n2990, CK => CLK, Q => n_3689, QN 
                           => n29118);
   clk_r_REG7883_S1 : DFF_X1 port map( D => n3423, CK => CLK, Q => n_3690, QN 
                           => n29117);
   clk_r_REG8364_S1 : DFF_X1 port map( D => n3519, CK => CLK, Q => n_3691, QN 
                           => n29116);
   clk_r_REG7667_S1 : DFF_X1 port map( D => n3360, CK => CLK, Q => n_3692, QN 
                           => n29115);
   clk_r_REG7575_S1 : DFF_X1 port map( D => n3328, CK => CLK, Q => n_3693, QN 
                           => n29114);
   clk_r_REG8222_S1 : DFF_X1 port map( D => n3488, CK => CLK, Q => n_3694, QN 
                           => n29113);
   clk_r_REG7881_S1 : DFF_X1 port map( D => n3424, CK => CLK, Q => n_3695, QN 
                           => n29112);
   clk_r_REG7573_S1 : DFF_X1 port map( D => n3329, CK => CLK, Q => n_3696, QN 
                           => n29111);
   clk_r_REG7963_S1 : DFF_X1 port map( D => n3392, CK => CLK, Q => n_3697, QN 
                           => n29110);
   clk_r_REG7961_S1 : DFF_X1 port map( D => n3393, CK => CLK, Q => n_3698, QN 
                           => n29109);
   clk_r_REG8362_S1 : DFF_X1 port map( D => n3520, CK => CLK, Q => n_3699, QN 
                           => n29108);
   clk_r_REG8220_S1 : DFF_X1 port map( D => n3489, CK => CLK, Q => n_3700, QN 
                           => n29107);
   clk_r_REG9837_S1 : DFF_X1 port map( D => n3456, CK => CLK, Q => n_3701, QN 
                           => n29106);
   clk_r_REG7665_S1 : DFF_X1 port map( D => n3361, CK => CLK, Q => n_3702, QN 
                           => n29105);
   clk_r_REG9835_S1 : DFF_X1 port map( D => n3457, CK => CLK, Q => n_3703, QN 
                           => n29104);
   clk_r_REG8360_S1 : DFF_X1 port map( D => n3521, CK => CLK, Q => n_3704, QN 
                           => n29103);
   clk_r_REG7879_S1 : DFF_X1 port map( D => n3425, CK => CLK, Q => n_3705, QN 
                           => n29102);
   clk_r_REG7877_S1 : DFF_X1 port map( D => n3426, CK => CLK, Q => n_3706, QN 
                           => n29101);
   clk_r_REG7875_S1 : DFF_X1 port map( D => n3427, CK => CLK, Q => n_3707, QN 
                           => n29100);
   clk_r_REG8358_S1 : DFF_X1 port map( D => n3522, CK => CLK, Q => n_3708, QN 
                           => n29099);
   clk_r_REG8356_S1 : DFF_X1 port map( D => n3523, CK => CLK, Q => n_3709, QN 
                           => n29098);
   clk_r_REG8354_S1 : DFF_X1 port map( D => n3524, CK => CLK, Q => n_3710, QN 
                           => n29097);
   clk_r_REG7873_S1 : DFF_X1 port map( D => n3428, CK => CLK, Q => n_3711, QN 
                           => n29096);
   clk_r_REG7309_S1 : DFF_X1 port map( D => n3525, CK => CLK, Q => n_3712, QN 
                           => n29095);
   clk_r_REG9833_S1 : DFF_X1 port map( D => n3458, CK => CLK, Q => n_3713, QN 
                           => n29094);
   clk_r_REG8218_S1 : DFF_X1 port map( D => n3490, CK => CLK, Q => n_3714, QN 
                           => n29093);
   clk_r_REG9831_S1 : DFF_X1 port map( D => n3459, CK => CLK, Q => n_3715, QN 
                           => n29092);
   clk_r_REG9829_S1 : DFF_X1 port map( D => n3460, CK => CLK, Q => n_3716, QN 
                           => n29091);
   clk_r_REG8216_S1 : DFF_X1 port map( D => n3491, CK => CLK, Q => n_3717, QN 
                           => n29090);
   clk_r_REG6935_S1 : DFF_X1 port map( D => n3461, CK => CLK, Q => n_3718, QN 
                           => n29089);
   clk_r_REG9887_S1 : DFF_X1 port map( D => n3431, CK => CLK, Q => n_3719, QN 
                           => n29088);
   clk_r_REG8412_S1 : DFF_X1 port map( D => n3495, CK => CLK, Q => n_3720, QN 
                           => n29087);
   clk_r_REG7571_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n_3721, QN 
                           => n29086);
   clk_r_REG7743_S1 : DFF_X1 port map( D => n3429, CK => CLK, Q => n_3722, QN 
                           => n29085);
   clk_r_REG8410_S1 : DFF_X1 port map( D => n3496, CK => CLK, Q => n_3723, QN 
                           => n29084);
   clk_r_REG8408_S1 : DFF_X1 port map( D => n3497, CK => CLK, Q => n_3724, QN 
                           => n29083);
   clk_r_REG9885_S1 : DFF_X1 port map( D => n3432, CK => CLK, Q => n_3725, QN 
                           => n29082);
   clk_r_REG9883_S1 : DFF_X1 port map( D => n3433, CK => CLK, Q => n_3726, QN 
                           => n29081);
   clk_r_REG7931_S1 : DFF_X1 port map( D => n3399, CK => CLK, Q => n_3727, QN 
                           => n29080);
   clk_r_REG7929_S1 : DFF_X1 port map( D => n3400, CK => CLK, Q => n_3728, QN 
                           => n29079);
   clk_r_REG7927_S1 : DFF_X1 port map( D => n3401, CK => CLK, Q => n_3729, QN 
                           => n29078);
   clk_r_REG7925_S1 : DFF_X1 port map( D => n3402, CK => CLK, Q => n_3730, QN 
                           => n29077);
   clk_r_REG9881_S1 : DFF_X1 port map( D => n3434, CK => CLK, Q => n_3731, QN 
                           => n29076);
   clk_r_REG8214_S1 : DFF_X1 port map( D => n3492, CK => CLK, Q => n_3732, QN 
                           => n29075);
   clk_r_REG8406_S1 : DFF_X1 port map( D => n3498, CK => CLK, Q => n_3733, QN 
                           => n29074);
   clk_r_REG7959_S1 : DFF_X1 port map( D => n3394, CK => CLK, Q => n_3734, QN 
                           => n29073);
   clk_r_REG8404_S1 : DFF_X1 port map( D => n3499, CK => CLK, Q => n_3735, QN 
                           => n29072);
   clk_r_REG7957_S1 : DFF_X1 port map( D => n3395, CK => CLK, Q => n_3736, QN 
                           => n29071);
   clk_r_REG7385_S1 : DFF_X1 port map( D => n3493, CK => CLK, Q => n_3737, QN 
                           => n29070);
   clk_r_REG7955_S1 : DFF_X1 port map( D => n3396, CK => CLK, Q => n_3738, QN 
                           => n29069);
   clk_r_REG7533_S1 : DFF_X1 port map( D => n3397, CK => CLK, Q => n_3739, QN 
                           => n29068);
   clk_r_REG9879_S1 : DFF_X1 port map( D => n3435, CK => CLK, Q => n_3740, QN 
                           => n29067);
   clk_r_REG7923_S1 : DFF_X1 port map( D => n3403, CK => CLK, Q => n_3741, QN 
                           => n29066);
   clk_r_REG8013_S1 : DFF_X1 port map( D => n3367, CK => CLK, Q => n_3742, QN 
                           => n29065);
   clk_r_REG8402_S1 : DFF_X1 port map( D => n3500, CK => CLK, Q => n_3743, QN 
                           => n29064);
   clk_r_REG8011_S1 : DFF_X1 port map( D => n3368, CK => CLK, Q => n_3744, QN 
                           => n29063);
   clk_r_REG8400_S1 : DFF_X1 port map( D => n3501, CK => CLK, Q => n_3745, QN 
                           => n29062);
   clk_r_REG8009_S1 : DFF_X1 port map( D => n3369, CK => CLK, Q => n_3746, QN 
                           => n29061);
   clk_r_REG8007_S1 : DFF_X1 port map( D => n3370, CK => CLK, Q => n_3747, QN 
                           => n29060);
   clk_r_REG9877_S1 : DFF_X1 port map( D => n3436, CK => CLK, Q => n_3748, QN 
                           => n29059);
   clk_r_REG8005_S1 : DFF_X1 port map( D => n3371, CK => CLK, Q => n_3749, QN 
                           => n29058);
   clk_r_REG8003_S1 : DFF_X1 port map( D => n3372, CK => CLK, Q => n_3750, QN 
                           => n29057);
   clk_r_REG7921_S1 : DFF_X1 port map( D => n3404, CK => CLK, Q => n_3751, QN 
                           => n29056);
   clk_r_REG9875_S1 : DFF_X1 port map( D => n3437, CK => CLK, Q => n_3752, QN 
                           => n29055);
   clk_r_REG7663_S1 : DFF_X1 port map( D => n3362, CK => CLK, Q => n_3753, QN 
                           => n29054);
   clk_r_REG7919_S1 : DFF_X1 port map( D => n3405, CK => CLK, Q => n_3754, QN 
                           => n29053);
   clk_r_REG8001_S1 : DFF_X1 port map( D => n3373, CK => CLK, Q => n_3755, QN 
                           => n29052);
   clk_r_REG7661_S1 : DFF_X1 port map( D => n3363, CK => CLK, Q => n_3756, QN 
                           => n29051);
   clk_r_REG7659_S1 : DFF_X1 port map( D => n3364, CK => CLK, Q => n_3757, QN 
                           => n29050);
   clk_r_REG7642_S1 : DFF_X1 port map( D => n3365, CK => CLK, Q => n_3758, QN 
                           => n29049);
   clk_r_REG7717_S1 : DFF_X1 port map( D => n3335, CK => CLK, Q => n_3759, QN 
                           => n29048);
   clk_r_REG7569_S1 : DFF_X1 port map( D => n3331, CK => CLK, Q => n_3760, QN 
                           => n29047);
   clk_r_REG7999_S1 : DFF_X1 port map( D => n3374, CK => CLK, Q => n_3761, QN 
                           => n29046);
   clk_r_REG8272_S1 : DFF_X1 port map( D => n3463, CK => CLK, Q => n_3762, QN 
                           => n29045);
   clk_r_REG7715_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n_3763, QN 
                           => n29044);
   clk_r_REG8270_S1 : DFF_X1 port map( D => n3464, CK => CLK, Q => n_3764, QN 
                           => n29043);
   clk_r_REG8268_S1 : DFF_X1 port map( D => n3465, CK => CLK, Q => n_3765, QN 
                           => n29042);
   clk_r_REG7713_S1 : DFF_X1 port map( D => n3337, CK => CLK, Q => n_3766, QN 
                           => n29041);
   clk_r_REG7711_S1 : DFF_X1 port map( D => n3338, CK => CLK, Q => n_3767, QN 
                           => n29040);
   clk_r_REG7709_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n_3768, QN 
                           => n29039);
   clk_r_REG7567_S1 : DFF_X1 port map( D => n3332, CK => CLK, Q => n_3769, QN 
                           => n29038);
   clk_r_REG8266_S1 : DFF_X1 port map( D => n3466, CK => CLK, Q => n_3770, QN 
                           => n29037);
   clk_r_REG8264_S1 : DFF_X1 port map( D => n3467, CK => CLK, Q => n_3771, QN 
                           => n29036);
   clk_r_REG7547_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n_3772, QN 
                           => n29035);
   clk_r_REG8262_S1 : DFF_X1 port map( D => n3468, CK => CLK, Q => n_3773, QN 
                           => n29034);
   clk_r_REG7627_S1 : DFF_X1 port map( D => n3302, CK => CLK, Q => n_3774, QN 
                           => n29033);
   clk_r_REG8398_S1 : DFF_X1 port map( D => n3502, CK => CLK, Q => n_3775, QN 
                           => n29032);
   clk_r_REG8260_S1 : DFF_X1 port map( D => n3469, CK => CLK, Q => n_3776, QN 
                           => n29031);
   clk_r_REG8258_S1 : DFF_X1 port map( D => n3470, CK => CLK, Q => n_3777, QN 
                           => n29030);
   clk_r_REG7707_S1 : DFF_X1 port map( D => n3340, CK => CLK, Q => n_3778, QN 
                           => n29029);
   clk_r_REG7625_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n_3779, QN 
                           => n29028);
   clk_r_REG9873_S1 : DFF_X1 port map( D => n3438, CK => CLK, Q => n_3780, QN 
                           => n29027);
   clk_r_REG7705_S1 : DFF_X1 port map( D => n3341, CK => CLK, Q => n_3781, QN 
                           => n29026);
   clk_r_REG7917_S1 : DFF_X1 port map( D => n3406, CK => CLK, Q => n_3782, QN 
                           => n29025);
   clk_r_REG7623_S1 : DFF_X1 port map( D => n3304, CK => CLK, Q => n_3783, QN 
                           => n29024);
   clk_r_REG7621_S1 : DFF_X1 port map( D => n3305, CK => CLK, Q => n_3784, QN 
                           => n29023);
   clk_r_REG7703_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n_3785, QN 
                           => n29022);
   clk_r_REG7619_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n_3786, QN 
                           => n29021);
   clk_r_REG7617_S1 : DFF_X1 port map( D => n3307, CK => CLK, Q => n_3787, QN 
                           => n29020);
   clk_r_REG7615_S1 : DFF_X1 port map( D => n3308, CK => CLK, Q => n_3788, QN 
                           => n29019);
   clk_r_REG7613_S1 : DFF_X1 port map( D => n3309, CK => CLK, Q => n_3789, QN 
                           => n29018);
   clk_r_REG10207_S7 : DFFR_X1 port map( D => n3576, CK => CLK, RN => RESET_BAR
                           , Q => n31216, QN => n_3790);
   clk_r_REG10136_S7 : DFFR_X1 port map( D => n3568, CK => CLK, RN => RESET_BAR
                           , Q => n31190, QN => n_3791);
   clk_r_REG10158_S7 : DFFS_X1 port map( D => n3564, CK => CLK, SN => RESET_BAR
                           , Q => n_3792, QN => n30052);
   clk_r_REG10137_S7 : DFFS_X1 port map( D => n3567, CK => CLK, SN => RESET_BAR
                           , Q => n_3793, QN => n30126);
   clk_r_REG10172_S7 : DFFS_X1 port map( D => n3562, CK => CLK, SN => RESET_BAR
                           , Q => n_3794, QN => n30128);
   clk_r_REG10151_S7 : DFFS_X1 port map( D => n3565, CK => CLK, SN => RESET_BAR
                           , Q => n_3795, QN => n30127);
   clk_r_REG10144_S7 : DFFR_X1 port map( D => n3566, CK => CLK, RN => RESET_BAR
                           , Q => n_3796, QN => n30051);
   clk_r_REG10215_S7 : DFFS_X1 port map( D => n3572, CK => CLK, SN => RESET_BAR
                           , Q => n_3797, QN => n30050);
   clk_r_REG10165_S7 : DFFS_X1 port map( D => n3561, CK => CLK, SN => RESET_BAR
                           , Q => n_3798, QN => n30125);
   clk_r_REG9982_S1 : DFFS_X2 port map( D => n18326, CK => CLK, SN => RESET_BAR
                           , Q => n30086, QN => n_3799);
   clk_r_REG9987_S1 : DFFS_X2 port map( D => n18331, CK => CLK, SN => RESET_BAR
                           , Q => n30091, QN => n_3800);
   clk_r_REG9988_S1 : DFFS_X2 port map( D => n18332, CK => CLK, SN => RESET_BAR
                           , Q => n30092, QN => n_3801);
   clk_r_REG9999_S1 : DFFS_X2 port map( D => n18335, CK => CLK, SN => RESET_BAR
                           , Q => n30095, QN => n_3802);
   clk_r_REG10004_S1 : DFFS_X2 port map( D => n18340, CK => CLK, SN => 
                           RESET_BAR, Q => n30100, QN => n_3803);
   clk_r_REG9990_S1 : DFFS_X2 port map( D => n18342, CK => CLK, SN => RESET_BAR
                           , Q => n30102, QN => n_3804);
   clk_r_REG9992_S1 : DFFS_X2 port map( D => n18344, CK => CLK, SN => RESET_BAR
                           , Q => n30104, QN => n_3805);
   clk_r_REG9994_S1 : DFFS_X2 port map( D => n18346, CK => CLK, SN => RESET_BAR
                           , Q => n30106, QN => n_3806);
   clk_r_REG9995_S1 : DFFS_X2 port map( D => n18347, CK => CLK, SN => RESET_BAR
                           , Q => n30107, QN => n_3807);
   clk_r_REG9996_S1 : DFFS_X2 port map( D => n18348, CK => CLK, SN => RESET_BAR
                           , Q => n30108, QN => n_3808);
   clk_r_REG10005_S1 : DFFS_X2 port map( D => n18349, CK => CLK, SN => 
                           RESET_BAR, Q => n30109, QN => n_3809);
   clk_r_REG10006_S1 : DFFS_X2 port map( D => n18351, CK => CLK, SN => 
                           RESET_BAR, Q => n30112, QN => n_3810);
   clk_r_REG10007_S1 : DFFS_X2 port map( D => n18353, CK => CLK, SN => 
                           RESET_BAR, Q => n30115, QN => n_3811);
   clk_r_REG10008_S1 : DFFS_X2 port map( D => n18354, CK => CLK, SN => 
                           RESET_BAR, Q => n30116, QN => n_3812);
   clk_r_REG10009_S1 : DFFS_X2 port map( D => n18355, CK => CLK, SN => 
                           RESET_BAR, Q => n30117, QN => n_3813);
   clk_r_REG10010_S1 : DFFS_X2 port map( D => n18357, CK => CLK, SN => 
                           RESET_BAR, Q => n30120, QN => n_3814);
   clk_r_REG10011_S1 : DFFS_X2 port map( D => n18359, CK => CLK, SN => 
                           RESET_BAR, Q => n30123, QN => n_3815);
   clk_r_REG10012_S1 : DFFS_X2 port map( D => n18360, CK => CLK, SN => 
                           RESET_BAR, Q => n30124, QN => n_3816);
   clk_r_REG9985_S1 : DFFS_X2 port map( D => n18329, CK => CLK, SN => RESET_BAR
                           , Q => n30089, QN => n_3817);
   clk_r_REG9986_S1 : DFFS_X2 port map( D => n18330, CK => CLK, SN => RESET_BAR
                           , Q => n30090, QN => n_3818);
   clk_r_REG9983_S1 : DFFS_X2 port map( D => n18327, CK => CLK, SN => RESET_BAR
                           , Q => n30087, QN => n_3819);
   clk_r_REG9984_S1 : DFFS_X2 port map( D => n18328, CK => CLK, SN => RESET_BAR
                           , Q => n30088, QN => n_3820);
   clk_r_REG9981_S1 : DFFS_X2 port map( D => n18325, CK => CLK, SN => RESET_BAR
                           , Q => n30085, QN => n_3821);
   clk_r_REG10001_S1 : DFFS_X2 port map( D => n18337, CK => CLK, SN => 
                           RESET_BAR, Q => n30097, QN => n_3822);
   clk_r_REG9989_S1 : DFFS_X2 port map( D => n18341, CK => CLK, SN => RESET_BAR
                           , Q => n30101, QN => n_3823);
   clk_r_REG9997_S1 : DFFS_X2 port map( D => n18333, CK => CLK, SN => RESET_BAR
                           , Q => n30093, QN => n_3824);
   clk_r_REG9998_S1 : DFFS_X2 port map( D => n18334, CK => CLK, SN => RESET_BAR
                           , Q => n30094, QN => n_3825);
   clk_r_REG10000_S1 : DFFS_X2 port map( D => n18336, CK => CLK, SN => 
                           RESET_BAR, Q => n30096, QN => n_3826);
   clk_r_REG10002_S1 : DFFS_X2 port map( D => n18338, CK => CLK, SN => 
                           RESET_BAR, Q => n30098, QN => n_3827);
   clk_r_REG10003_S1 : DFFS_X2 port map( D => n18339, CK => CLK, SN => 
                           RESET_BAR, Q => n30099, QN => n_3828);
   clk_r_REG9991_S1 : DFFS_X2 port map( D => n18343, CK => CLK, SN => RESET_BAR
                           , Q => n30103, QN => n_3829);
   clk_r_REG9993_S1 : DFFS_X2 port map( D => n18345, CK => CLK, SN => RESET_BAR
                           , Q => n30105, QN => n_3830);
   U3 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30094, ZN => n36813);
   U4 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30098, ZN => n36833);
   U5 : CLKBUF_X1 port map( A => n37627, Z => n37448);
   U6 : CLKBUF_X1 port map( A => n38342, Z => n38295);
   U7 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => ADD_RD1(2),
                           ZN => n19400);
   U8 : INV_X1 port map( A => n19400, ZN => n3566);
   U9 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), ZN => n35761);
   U10 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n35761, ZN => n19395);
   U11 : INV_X1 port map( A => n19395, ZN => n3561);
   U12 : INV_X1 port map( A => ADD_RD1(1), ZN => n35766);
   U13 : NOR2_X1 port map( A1 => n35766, A2 => n35761, ZN => n19398);
   U14 : INV_X1 port map( A => n19398, ZN => n3562);
   U15 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => ADD_RD2(2)
                           , ZN => n3570);
   U16 : INV_X1 port map( A => ADD_RD2(2), ZN => n35767);
   U17 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n35767, ZN => n35763);
   U18 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => n35763, ZN => n3571);
   U19 : INV_X1 port map( A => ADD_RD2(1), ZN => n35768);
   U20 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), ZN => n35762);
   U21 : NOR2_X1 port map( A1 => n35768, A2 => n35762, ZN => n3575);
   U22 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => n35762, ZN => n3577);
   U23 : NOR2_X1 port map( A1 => n35768, A2 => n35763, ZN => n3576);
   U24 : INV_X1 port map( A => ADD_RD1(2), ZN => n35764);
   U25 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => n35764, ZN
                           => n3568);
   U26 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n35766, ZN
                           => n19399);
   U27 : INV_X1 port map( A => n19399, ZN => n3564);
   U28 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => n35766, A3 => n35764, ZN => 
                           n3563);
   U29 : INV_X1 port map( A => ADD_RD1(3), ZN => n3560);
   U30 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n35764, ZN => n35765);
   U31 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n35765, ZN => n19396);
   U32 : INV_X1 port map( A => n19396, ZN => n3567);
   U33 : NOR2_X1 port map( A1 => n35766, A2 => n35765, ZN => n19397);
   U34 : INV_X1 port map( A => n19397, ZN => n3565);
   U35 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => n35767, ZN
                           => n3573);
   U36 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n35768, ZN
                           => n19402);
   U37 : INV_X1 port map( A => n19402, ZN => n3572);
   U38 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => n35768, A3 => n35767, ZN => 
                           n3574);
   U39 : INV_X1 port map( A => ADD_RD2(3), ZN => n3569);
   U40 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31248, ZN => n36748);
   U41 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30112, ZN => n36519);
   U42 : OAI22_X1 port map( A1 => n30112, A2 => n36748, B1 => n30267, B2 => 
                           n36519, ZN => n35769);
   U43 : INV_X1 port map( A => n35769, ZN => n3096);
   U44 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31235, ZN => n36425);
   U45 : CLKBUF_X1 port map( A => n36425, Z => n36321);
   U46 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30087, ZN => n36543);
   U47 : OAI22_X1 port map( A1 => n30087, A2 => n36321, B1 => n30430, B2 => 
                           n36543, ZN => n35770);
   U48 : INV_X1 port map( A => n35770, ZN => n3494);
   U49 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31240, ZN => n36454);
   U50 : OAI22_X1 port map( A1 => n30087, A2 => n36454, B1 => n30427, B2 => 
                           n36543, ZN => n35771);
   U51 : INV_X1 port map( A => n35771, ZN => n3352);
   U52 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31236, ZN => n36403);
   U53 : OAI22_X1 port map( A1 => n30087, A2 => n36403, B1 => n30431, B2 => 
                           n36543, ZN => n35772);
   U54 : INV_X1 port map( A => n35772, ZN => n3481);
   U55 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30088, ZN => n36535);
   U56 : OAI22_X1 port map( A1 => n30088, A2 => n36425, B1 => n30433, B2 => 
                           n36535, ZN => n35773);
   U57 : INV_X1 port map( A => n35773, ZN => n3514);
   U58 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31245, ZN => n36485);
   U59 : OAI22_X1 port map( A1 => n30112, A2 => n36485, B1 => n30315, B2 => 
                           n36519, ZN => n35774);
   U60 : INV_X1 port map( A => n35774, ZN => n3195);
   U61 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30090, ZN => n36511);
   U62 : OAI22_X1 port map( A1 => n30090, A2 => n36425, B1 => n30425, B2 => 
                           n36511, ZN => n35775);
   U63 : INV_X1 port map( A => n35775, ZN => n3512);
   U64 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31238, ZN => n36441);
   U65 : OAI22_X1 port map( A1 => n30088, A2 => n36441, B1 => n30437, B2 => 
                           n36535, ZN => n35776);
   U66 : INV_X1 port map( A => n35776, ZN => n3417);
   U67 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31239, ZN => n36469);
   U68 : CLKBUF_X1 port map( A => n36469, Z => n36303);
   U69 : OAI22_X1 port map( A1 => n30088, A2 => n36303, B1 => n30438, B2 => 
                           n36535, ZN => n35777);
   U70 : INV_X1 port map( A => n35777, ZN => n3366);
   U71 : CLKBUF_X1 port map( A => n36441, Z => n36315);
   U72 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30089, ZN => n36522);
   U73 : OAI22_X1 port map( A1 => n30089, A2 => n36315, B1 => n30439, B2 => 
                           n36522, ZN => n35778);
   U74 : INV_X1 port map( A => n35778, ZN => n3398);
   U75 : OAI22_X1 port map( A1 => n30087, A2 => n36469, B1 => n30440, B2 => 
                           n36543, ZN => n35779);
   U76 : INV_X1 port map( A => n35779, ZN => n3386);
   U77 : CLKBUF_X1 port map( A => n36403, Z => n36282);
   U78 : OAI22_X1 port map( A1 => n30089, A2 => n36282, B1 => n30441, B2 => 
                           n36522, ZN => n35780);
   U79 : INV_X1 port map( A => n35780, ZN => n3462);
   U80 : OAI22_X1 port map( A1 => n30090, A2 => n36441, B1 => n30442, B2 => 
                           n36511, ZN => n35781);
   U81 : INV_X1 port map( A => n35781, ZN => n3418);
   U82 : OAI22_X1 port map( A1 => n30087, A2 => n36441, B1 => n30443, B2 => 
                           n36543, ZN => n35782);
   U83 : INV_X1 port map( A => n35782, ZN => n3419);
   U84 : OAI22_X1 port map( A1 => n30090, A2 => n36454, B1 => n30444, B2 => 
                           n36511, ZN => n35783);
   U85 : INV_X1 port map( A => n35783, ZN => n3354);
   U86 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31237, ZN => n36327);
   U87 : CLKBUF_X1 port map( A => n36327, Z => n36489);
   U88 : OAI22_X1 port map( A1 => n30089, A2 => n36489, B1 => n30445, B2 => 
                           n36522, ZN => n35784);
   U89 : INV_X1 port map( A => n35784, ZN => n3430);
   U90 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31253, ZN => n36718);
   U91 : OAI22_X1 port map( A1 => n30112, A2 => n36718, B1 => n30338, B2 => 
                           n36519, ZN => n35785);
   U92 : INV_X1 port map( A => n35785, ZN => n2939);
   U93 : OAI22_X1 port map( A1 => n30089, A2 => n36454, B1 => n30446, B2 => 
                           n36522, ZN => n35786);
   U94 : INV_X1 port map( A => n35786, ZN => n3355);
   U95 : OAI22_X1 port map( A1 => n30090, A2 => n36403, B1 => n30447, B2 => 
                           n36511, ZN => n35787);
   U96 : INV_X1 port map( A => n35787, ZN => n3482);
   U97 : OAI22_X1 port map( A1 => n30090, A2 => n36327, B1 => n30448, B2 => 
                           n36511, ZN => n35788);
   U98 : INV_X1 port map( A => n35788, ZN => n3450);
   U99 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31234, ZN => n36493);
   U100 : OAI22_X1 port map( A1 => n30090, A2 => n36493, B1 => n30339, B2 => 
                           n36511, ZN => n35789);
   U101 : INV_X1 port map( A => n35789, ZN => n3535);
   U102 : OAI22_X1 port map( A1 => n30089, A2 => n36469, B1 => n30449, B2 => 
                           n36522, ZN => n35790);
   U103 : INV_X1 port map( A => n35790, ZN => n3387);
   U104 : OAI22_X1 port map( A1 => n30089, A2 => n36425, B1 => n30450, B2 => 
                           n36522, ZN => n35791);
   U105 : INV_X1 port map( A => n35791, ZN => n3515);
   U106 : OAI22_X1 port map( A1 => n30088, A2 => n36327, B1 => n30451, B2 => 
                           n36535, ZN => n35792);
   U107 : INV_X1 port map( A => n35792, ZN => n3451);
   U108 : OAI22_X1 port map( A1 => n30088, A2 => n36403, B1 => n30452, B2 => 
                           n36535, ZN => n35793);
   U109 : INV_X1 port map( A => n35793, ZN => n3483);
   U110 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31252, ZN => n36662);
   U111 : OAI22_X1 port map( A1 => n30112, A2 => n36662, B1 => n30332, B2 => 
                           n36519, ZN => n35794);
   U112 : INV_X1 port map( A => n35794, ZN => n2970);
   U113 : OAI22_X1 port map( A1 => n30089, A2 => n36493, B1 => n30342, B2 => 
                           n36522, ZN => n35795);
   U114 : INV_X1 port map( A => n35795, ZN => n3538);
   U115 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31244, ZN => n36643);
   U116 : CLKBUF_X1 port map( A => n36643, Z => n36184);
   U117 : OAI22_X1 port map( A1 => n30087, A2 => n36184, B1 => n30457, B2 => 
                           n36543, ZN => n35796);
   U118 : INV_X1 port map( A => n35796, ZN => n3219);
   U119 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31243, ZN => n36674);
   U120 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30108, ZN => n36538);
   U121 : OAI22_X1 port map( A1 => n30108, A2 => n36674, B1 => n30461, B2 => 
                           n36538, ZN => n35797);
   U122 : INV_X1 port map( A => n35797, ZN => n3260);
   U123 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30106, ZN => n36550);
   U124 : OAI22_X1 port map( A1 => n30106, A2 => n36184, B1 => n30462, B2 => 
                           n36550, ZN => n35798);
   U125 : INV_X1 port map( A => n35798, ZN => n3221);
   U126 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31247, ZN => n36712);
   U127 : OAI22_X1 port map( A1 => n30106, A2 => n36712, B1 => n30464, B2 => 
                           n36550, ZN => n35799);
   U128 : INV_X1 port map( A => n35799, ZN => n3134);
   U129 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31242, ZN => n36457);
   U130 : OAI22_X1 port map( A1 => n30106, A2 => n36457, B1 => n30467, B2 => 
                           n36550, ZN => n35800);
   U131 : INV_X1 port map( A => n35800, ZN => n3292);
   U132 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30107, ZN => n36525);
   U133 : OAI22_X1 port map( A1 => n30107, A2 => n36485, B1 => n30469, B2 => 
                           n36525, ZN => n35801);
   U134 : INV_X1 port map( A => n35801, ZN => n3196);
   U135 : OAI22_X1 port map( A1 => n30112, A2 => n36469, B1 => n30347, B2 => 
                           n36519, ZN => n35802);
   U136 : INV_X1 port map( A => n35802, ZN => n3377);
   U137 : OAI22_X1 port map( A1 => n30107, A2 => n36712, B1 => n30471, B2 => 
                           n36525, ZN => n35803);
   U138 : INV_X1 port map( A => n35803, ZN => n3135);
   U139 : OAI22_X1 port map( A1 => n30106, A2 => n36485, B1 => n30472, B2 => 
                           n36550, ZN => n35804);
   U140 : INV_X1 port map( A => n35804, ZN => n3197);
   U141 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31246, ZN => n36783);
   U142 : OAI22_X1 port map( A1 => n30106, A2 => n36783, B1 => n30473, B2 => 
                           n36550, ZN => n35805);
   U143 : INV_X1 port map( A => n35805, ZN => n3164);
   U144 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31255, ZN => n36715);
   U145 : OAI22_X1 port map( A1 => n30108, A2 => n36715, B1 => n30474, B2 => 
                           n36538, ZN => n35806);
   U146 : INV_X1 port map( A => n35806, ZN => n2876);
   U147 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31250, ZN => n36683);
   U148 : OAI22_X1 port map( A1 => n30108, A2 => n36683, B1 => n30475, B2 => 
                           n36538, ZN => n35807);
   U149 : INV_X1 port map( A => n35807, ZN => n3038);
   U150 : OAI22_X1 port map( A1 => n30106, A2 => n36748, B1 => n30477, B2 => 
                           n36550, ZN => n35808);
   U151 : INV_X1 port map( A => n35808, ZN => n3100);
   U152 : OAI22_X1 port map( A1 => n30112, A2 => n36712, B1 => n30279, B2 => 
                           n36519, ZN => n35809);
   U153 : INV_X1 port map( A => n35809, ZN => n3127);
   U154 : CLKBUF_X1 port map( A => n36712, Z => n36431);
   U155 : OAI22_X1 port map( A1 => n30108, A2 => n36431, B1 => n30481, B2 => 
                           n36538, ZN => n35810);
   U156 : INV_X1 port map( A => n35810, ZN => n3110);
   U157 : OAI22_X1 port map( A1 => n30108, A2 => n36718, B1 => n30482, B2 => 
                           n36538, ZN => n35811);
   U158 : INV_X1 port map( A => n35811, ZN => n2940);
   U159 : OAI22_X1 port map( A1 => n30106, A2 => n36662, B1 => n30483, B2 => 
                           n36550, ZN => n35812);
   U160 : INV_X1 port map( A => n35812, ZN => n2973);
   U161 : OAI22_X1 port map( A1 => n30106, A2 => n36718, B1 => n30484, B2 => 
                           n36550, ZN => n35813);
   U162 : INV_X1 port map( A => n35813, ZN => n2941);
   U163 : OAI22_X1 port map( A1 => n30112, A2 => n36454, B1 => n30353, B2 => 
                           n36519, ZN => n35814);
   U164 : INV_X1 port map( A => n35814, ZN => n3346);
   U165 : OAI22_X1 port map( A1 => n30090, A2 => n36469, B1 => n30420, B2 => 
                           n36511, ZN => n35815);
   U166 : INV_X1 port map( A => n35815, ZN => n3383);
   U167 : OAI22_X1 port map( A1 => n30107, A2 => n36718, B1 => n30487, B2 => 
                           n36525, ZN => n35816);
   U168 : INV_X1 port map( A => n35816, ZN => n2942);
   U169 : OAI22_X1 port map( A1 => n30108, A2 => n36485, B1 => n30489, B2 => 
                           n36538, ZN => n35817);
   U170 : INV_X1 port map( A => n35817, ZN => n3198);
   U171 : OAI22_X1 port map( A1 => n30087, A2 => n36327, B1 => n30417, B2 => 
                           n36543, ZN => n35818);
   U172 : INV_X1 port map( A => n35818, ZN => n3447);
   U173 : CLKBUF_X1 port map( A => n36683, Z => n36579);
   U174 : OAI22_X1 port map( A1 => n30107, A2 => n36579, B1 => n30492, B2 => 
                           n36525, ZN => n35819);
   U175 : INV_X1 port map( A => n35819, ZN => n3014);
   U176 : OAI22_X1 port map( A1 => n30088, A2 => n36454, B1 => n30428, B2 => 
                           n36535, ZN => n35820);
   U177 : INV_X1 port map( A => n35820, ZN => n3353);
   U178 : OAI22_X1 port map( A1 => n30112, A2 => n36493, B1 => n30410, B2 => 
                           n36519, ZN => n35821);
   U179 : INV_X1 port map( A => n35821, ZN => n3542);
   U180 : OAI22_X1 port map( A1 => n30089, A2 => n36457, B1 => n30187, B2 => 
                           n36522, ZN => n35822);
   U181 : INV_X1 port map( A => n35822, ZN => n3281);
   U182 : OAI22_X1 port map( A1 => n30088, A2 => n36715, B1 => n30191, B2 => 
                           n36535, ZN => n35823);
   U183 : INV_X1 port map( A => n35823, ZN => n2866);
   U184 : OAI22_X1 port map( A1 => n30088, A2 => n36718, B1 => n30192, B2 => 
                           n36535, ZN => n35824);
   U185 : INV_X1 port map( A => n35824, ZN => n2930);
   U186 : OAI22_X1 port map( A1 => n30088, A2 => n36662, B1 => n30193, B2 => 
                           n36535, ZN => n35825);
   U187 : INV_X1 port map( A => n35825, ZN => n2962);
   U188 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31251, ZN => n36398);
   U189 : OAI22_X1 port map( A1 => n30112, A2 => n36398, B1 => n30402, B2 => 
                           n36519, ZN => n35826);
   U190 : INV_X1 port map( A => n35826, ZN => n3000);
   U191 : OAI22_X1 port map( A1 => n30087, A2 => n36457, B1 => n30199, B2 => 
                           n36543, ZN => n35827);
   U192 : INV_X1 port map( A => n35827, ZN => n3282);
   U193 : OAI22_X1 port map( A1 => n30088, A2 => n36485, B1 => n30201, B2 => 
                           n36535, ZN => n35828);
   U194 : INV_X1 port map( A => n35828, ZN => n3185);
   U195 : OAI22_X1 port map( A1 => n30088, A2 => n36674, B1 => n30202, B2 => 
                           n36535, ZN => n35829);
   U196 : INV_X1 port map( A => n35829, ZN => n3249);
   U197 : OAI22_X1 port map( A1 => n30088, A2 => n36398, B1 => n30203, B2 => 
                           n36535, ZN => n35830);
   U198 : INV_X1 port map( A => n35830, ZN => n2996);
   U199 : CLKBUF_X1 port map( A => n36457, Z => n36420);
   U200 : OAI22_X1 port map( A1 => n30088, A2 => n36420, B1 => n30204, B2 => 
                           n36535, ZN => n35831);
   U201 : INV_X1 port map( A => n35831, ZN => n3283);
   U202 : OAI22_X1 port map( A1 => n30088, A2 => n36579, B1 => n30205, B2 => 
                           n36535, ZN => n35832);
   U203 : INV_X1 port map( A => n35832, ZN => n3028);
   U204 : CLKBUF_X1 port map( A => n36748, Z => n36433);
   U205 : OAI22_X1 port map( A1 => n30088, A2 => n36433, B1 => n30209, B2 => 
                           n36535, ZN => n35833);
   U206 : INV_X1 port map( A => n35833, ZN => n3091);
   U207 : OAI22_X1 port map( A1 => n30088, A2 => n36431, B1 => n30211, B2 => 
                           n36535, ZN => n35834);
   U208 : INV_X1 port map( A => n35834, ZN => n3123);
   U209 : OAI22_X1 port map( A1 => n30087, A2 => n36783, B1 => n30213, B2 => 
                           n36543, ZN => n35835);
   U210 : INV_X1 port map( A => n35835, ZN => n3153);
   U211 : CLKBUF_X1 port map( A => n36662, Z => n36692);
   U212 : OAI22_X1 port map( A1 => n30087, A2 => n36692, B1 => n30216, B2 => 
                           n36543, ZN => n35836);
   U213 : INV_X1 port map( A => n35836, ZN => n2964);
   U214 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31249, ZN => n36449);
   U215 : OAI22_X1 port map( A1 => n30087, A2 => n36449, B1 => n30218, B2 => 
                           n36543, ZN => n35837);
   U216 : INV_X1 port map( A => n35837, ZN => n3060);
   U217 : CLKBUF_X1 port map( A => n36718, Z => n36701);
   U218 : OAI22_X1 port map( A1 => n30087, A2 => n36701, B1 => n30219, B2 => 
                           n36543, ZN => n35838);
   U219 : INV_X1 port map( A => n35838, ZN => n2932);
   U220 : OAI22_X1 port map( A1 => n30112, A2 => n36425, B1 => n30382, B2 => 
                           n36519, ZN => n35839);
   U221 : INV_X1 port map( A => n35839, ZN => n3503);
   U222 : CLKBUF_X1 port map( A => n36783, Z => n36429);
   U223 : OAI22_X1 port map( A1 => n30088, A2 => n36429, B1 => n30225, B2 => 
                           n36535, ZN => n35840);
   U224 : INV_X1 port map( A => n35840, ZN => n3155);
   U225 : OAI22_X1 port map( A1 => n30112, A2 => n36489, B1 => n30377, B2 => 
                           n36519, ZN => n35841);
   U226 : INV_X1 port map( A => n35841, ZN => n3443);
   U227 : CLKBUF_X1 port map( A => n36715, Z => n36477);
   U228 : OAI22_X1 port map( A1 => n30087, A2 => n36477, B1 => n30226, B2 => 
                           n36543, ZN => n35842);
   U229 : INV_X1 port map( A => n35842, ZN => n2868);
   U230 : CLKBUF_X1 port map( A => n36485, Z => n36427);
   U231 : OAI22_X1 port map( A1 => n30087, A2 => n36427, B1 => n30229, B2 => 
                           n36543, ZN => n35843);
   U232 : INV_X1 port map( A => n35843, ZN => n3187);
   U233 : OAI22_X1 port map( A1 => n30087, A2 => n36748, B1 => n30230, B2 => 
                           n36543, ZN => n35844);
   U234 : INV_X1 port map( A => n35844, ZN => n3092);
   U235 : OAI22_X1 port map( A1 => n30087, A2 => n36431, B1 => n30231, B2 => 
                           n36543, ZN => n35845);
   U236 : INV_X1 port map( A => n35845, ZN => n3125);
   U237 : OAI22_X1 port map( A1 => n30112, A2 => n36403, B1 => n30371, B2 => 
                           n36519, ZN => n35846);
   U238 : INV_X1 port map( A => n35846, ZN => n3471);
   U239 : OAI22_X1 port map( A1 => n30112, A2 => n36683, B1 => n30314, B2 => 
                           n36519, ZN => n35847);
   U240 : INV_X1 port map( A => n35847, ZN => n3035);
   U241 : OAI22_X1 port map( A1 => n30112, A2 => n36441, B1 => n30369, B2 => 
                           n36519, ZN => n35848);
   U242 : INV_X1 port map( A => n35848, ZN => n3407);
   U243 : OAI22_X1 port map( A1 => n30112, A2 => n36457, B1 => n30254, B2 => 
                           n36519, ZN => n35849);
   U244 : INV_X1 port map( A => n35849, ZN => n3291);
   U245 : OAI22_X1 port map( A1 => n30112, A2 => n36449, B1 => n30357, B2 => 
                           n36519, ZN => n35850);
   U246 : INV_X1 port map( A => n35850, ZN => n3064);
   U247 : OAI22_X1 port map( A1 => n30090, A2 => n36457, B1 => n30157, B2 => 
                           n36511, ZN => n35851);
   U248 : INV_X1 port map( A => n35851, ZN => n3279);
   U249 : OAI22_X1 port map( A1 => n30090, A2 => n36674, B1 => n30158, B2 => 
                           n36511, ZN => n35852);
   U250 : INV_X1 port map( A => n35852, ZN => n3246);
   U251 : OAI22_X1 port map( A1 => n30090, A2 => n36485, B1 => n30159, B2 => 
                           n36511, ZN => n35853);
   U252 : INV_X1 port map( A => n35853, ZN => n3182);
   U253 : OAI22_X1 port map( A1 => n30090, A2 => n36783, B1 => n30160, B2 => 
                           n36511, ZN => n35854);
   U254 : INV_X1 port map( A => n35854, ZN => n3150);
   U255 : OAI22_X1 port map( A1 => n30090, A2 => n36712, B1 => n30161, B2 => 
                           n36511, ZN => n35855);
   U256 : INV_X1 port map( A => n35855, ZN => n3120);
   U257 : OAI22_X1 port map( A1 => n30090, A2 => n36748, B1 => n30162, B2 => 
                           n36511, ZN => n35856);
   U258 : INV_X1 port map( A => n35856, ZN => n3088);
   U259 : OAI22_X1 port map( A1 => n30087, A2 => n36398, B1 => n30164, B2 => 
                           n36543, ZN => n35857);
   U260 : INV_X1 port map( A => n35857, ZN => n2992);
   U261 : OAI22_X1 port map( A1 => n30090, A2 => n36449, B1 => n30165, B2 => 
                           n36511, ZN => n35858);
   U262 : INV_X1 port map( A => n35858, ZN => n3056);
   U263 : OAI22_X1 port map( A1 => n30090, A2 => n36683, B1 => n30166, B2 => 
                           n36511, ZN => n35859);
   U264 : INV_X1 port map( A => n35859, ZN => n3025);
   U265 : OAI22_X1 port map( A1 => n30090, A2 => n36398, B1 => n30167, B2 => 
                           n36511, ZN => n35860);
   U266 : INV_X1 port map( A => n35860, ZN => n2993);
   U267 : OAI22_X1 port map( A1 => n30090, A2 => n36662, B1 => n30168, B2 => 
                           n36511, ZN => n35861);
   U268 : INV_X1 port map( A => n35861, ZN => n2960);
   U269 : OAI22_X1 port map( A1 => n30090, A2 => n36718, B1 => n30169, B2 => 
                           n36511, ZN => n35862);
   U270 : INV_X1 port map( A => n35862, ZN => n2928);
   U271 : OAI22_X1 port map( A1 => n30089, A2 => n36449, B1 => n30170, B2 => 
                           n36522, ZN => n35863);
   U272 : INV_X1 port map( A => n35863, ZN => n3057);
   U273 : OAI22_X1 port map( A1 => n30089, A2 => n36398, B1 => n30171, B2 => 
                           n36522, ZN => n35864);
   U274 : INV_X1 port map( A => n35864, ZN => n2994);
   U275 : OAI22_X1 port map( A1 => n30089, A2 => n36748, B1 => n30172, B2 => 
                           n36522, ZN => n35865);
   U276 : INV_X1 port map( A => n35865, ZN => n3089);
   U277 : OAI22_X1 port map( A1 => n30089, A2 => n36712, B1 => n30174, B2 => 
                           n36522, ZN => n35866);
   U278 : INV_X1 port map( A => n35866, ZN => n3121);
   U279 : OAI22_X1 port map( A1 => n30089, A2 => n36485, B1 => n30176, B2 => 
                           n36522, ZN => n35867);
   U280 : INV_X1 port map( A => n35867, ZN => n3183);
   U281 : OAI22_X1 port map( A1 => n30089, A2 => n36662, B1 => n30177, B2 => 
                           n36522, ZN => n35868);
   U282 : INV_X1 port map( A => n35868, ZN => n2961);
   U283 : OAI22_X1 port map( A1 => n30089, A2 => n36674, B1 => n30178, B2 => 
                           n36522, ZN => n35869);
   U284 : INV_X1 port map( A => n35869, ZN => n3247);
   U285 : OAI22_X1 port map( A1 => n30089, A2 => n36715, B1 => n30184, B2 => 
                           n36522, ZN => n35870);
   U286 : INV_X1 port map( A => n35870, ZN => n2865);
   U287 : OAI22_X1 port map( A1 => n30087, A2 => n36493, B1 => n30341, B2 => 
                           n36543, ZN => n35871);
   U288 : INV_X1 port map( A => n35871, ZN => n3537);
   U289 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30103, ZN => n36508);
   U290 : OAI22_X1 port map( A1 => n30103, A2 => n36449, B1 => n30757, B2 => 
                           n36508, ZN => n35872);
   U291 : INV_X1 port map( A => n35872, ZN => n3077);
   U292 : OAI22_X1 port map( A1 => n30103, A2 => n36433, B1 => n30764, B2 => 
                           n36508, ZN => n35873);
   U293 : INV_X1 port map( A => n35873, ZN => n3082);
   U294 : OAI22_X1 port map( A1 => n30103, A2 => n36431, B1 => n30767, B2 => 
                           n36508, ZN => n35874);
   U295 : INV_X1 port map( A => n35874, ZN => n3115);
   U296 : OAI22_X1 port map( A1 => n30103, A2 => n36429, B1 => n30768, B2 => 
                           n36508, ZN => n35875);
   U297 : INV_X1 port map( A => n35875, ZN => n3145);
   U298 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30101, ZN => n36514);
   U299 : OAI22_X1 port map( A1 => n30101, A2 => n36420, B1 => n30769, B2 => 
                           n36514, ZN => n35876);
   U300 : INV_X1 port map( A => n35876, ZN => n3275);
   U301 : CLKBUF_X1 port map( A => n36674, Z => n36422);
   U302 : OAI22_X1 port map( A1 => n30101, A2 => n36422, B1 => n30770, B2 => 
                           n36514, ZN => n35877);
   U303 : INV_X1 port map( A => n35877, ZN => n3242);
   U304 : OAI22_X1 port map( A1 => n30103, A2 => n36427, B1 => n30773, B2 => 
                           n36508, ZN => n35878);
   U305 : INV_X1 port map( A => n35878, ZN => n3178);
   U306 : OAI22_X1 port map( A1 => n30103, A2 => n36422, B1 => n30774, B2 => 
                           n36508, ZN => n35879);
   U307 : INV_X1 port map( A => n35879, ZN => n3243);
   U308 : OAI22_X1 port map( A1 => n30103, A2 => n36420, B1 => n30775, B2 => 
                           n36508, ZN => n35880);
   U309 : INV_X1 port map( A => n35880, ZN => n3276);
   U310 : OAI22_X1 port map( A1 => n30101, A2 => n36427, B1 => n30776, B2 => 
                           n36514, ZN => n35881);
   U311 : INV_X1 port map( A => n35881, ZN => n3177);
   U312 : OAI22_X1 port map( A1 => n30101, A2 => n36429, B1 => n30777, B2 => 
                           n36514, ZN => n35882);
   U313 : INV_X1 port map( A => n35882, ZN => n3146);
   U314 : OAI22_X1 port map( A1 => n30101, A2 => n36431, B1 => n30778, B2 => 
                           n36514, ZN => n35883);
   U315 : INV_X1 port map( A => n35883, ZN => n3116);
   U316 : OAI22_X1 port map( A1 => n30101, A2 => n36433, B1 => n30784, B2 => 
                           n36514, ZN => n35884);
   U317 : INV_X1 port map( A => n35884, ZN => n3083);
   U318 : OAI22_X1 port map( A1 => n30101, A2 => n36692, B1 => n30786, B2 => 
                           n36514, ZN => n35885);
   U319 : INV_X1 port map( A => n35885, ZN => n2955);
   U320 : OAI22_X1 port map( A1 => n30101, A2 => n36701, B1 => n30787, B2 => 
                           n36514, ZN => n35886);
   U321 : INV_X1 port map( A => n35886, ZN => n2923);
   U322 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31254, ZN => n36472);
   U323 : OAI22_X1 port map( A1 => n30101, A2 => n36472, B1 => n30788, B2 => 
                           n36514, ZN => n35887);
   U324 : INV_X1 port map( A => n35887, ZN => n2909);
   U325 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31256, ZN => n36487);
   U326 : OAI22_X1 port map( A1 => n30101, A2 => n36487, B1 => n30789, B2 => 
                           n36514, ZN => n35888);
   U327 : INV_X1 port map( A => n35888, ZN => n2849);
   U328 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31257, ZN => n36730);
   U329 : OAI22_X1 port map( A1 => n30101, A2 => n36730, B1 => n30793, B2 => 
                           n36514, ZN => n35889);
   U330 : INV_X1 port map( A => n35889, ZN => n2817);
   U331 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30093, ZN => n36606);
   U332 : OAI22_X1 port map( A1 => n30093, A2 => n36715, B1 => n30825, B2 => 
                           n36606, ZN => n35890);
   U333 : INV_X1 port map( A => n35890, ZN => n2883);
   U334 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30099, ZN => n36572);
   U335 : OAI22_X1 port map( A1 => n30099, A2 => n36730, B1 => n30828, B2 => 
                           n36572, ZN => n35891);
   U336 : INV_X1 port map( A => n35891, ZN => n2818);
   U337 : OAI22_X1 port map( A1 => n30099, A2 => n36487, B1 => n30829, B2 => 
                           n36572, ZN => n35892);
   U338 : INV_X1 port map( A => n35892, ZN => n2850);
   U339 : OAI22_X1 port map( A1 => n30099, A2 => n36472, B1 => n30830, B2 => 
                           n36572, ZN => n35893);
   U340 : INV_X1 port map( A => n35893, ZN => n2910);
   U341 : OAI22_X1 port map( A1 => n30099, A2 => n36701, B1 => n30831, B2 => 
                           n36572, ZN => n35894);
   U342 : INV_X1 port map( A => n35894, ZN => n2925);
   U343 : OAI22_X1 port map( A1 => n30103, A2 => n36477, B1 => n30833, B2 => 
                           n36508, ZN => n35895);
   U344 : INV_X1 port map( A => n35895, ZN => n2856);
   U345 : OAI22_X1 port map( A1 => n30101, A2 => n36477, B1 => n30835, B2 => 
                           n36514, ZN => n35896);
   U346 : INV_X1 port map( A => n35896, ZN => n2858);
   U347 : OAI22_X1 port map( A1 => n30099, A2 => n36477, B1 => n30837, B2 => 
                           n36572, ZN => n35897);
   U348 : INV_X1 port map( A => n35897, ZN => n2860);
   U349 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30097, ZN => n36609);
   U350 : OAI22_X1 port map( A1 => n30097, A2 => n36477, B1 => n30838, B2 => 
                           n36609, ZN => n35898);
   U351 : INV_X1 port map( A => n35898, ZN => n2861);
   U352 : OAI22_X1 port map( A1 => n30099, A2 => n36692, B1 => n30839, B2 => 
                           n36572, ZN => n35899);
   U353 : INV_X1 port map( A => n35899, ZN => n2957);
   U354 : CLKBUF_X1 port map( A => n36449, Z => n36677);
   U355 : OAI22_X1 port map( A1 => n30099, A2 => n36677, B1 => n30840, B2 => 
                           n36572, ZN => n35900);
   U356 : INV_X1 port map( A => n35900, ZN => n3049);
   U357 : OAI22_X1 port map( A1 => n30099, A2 => n36433, B1 => n30841, B2 => 
                           n36572, ZN => n35901);
   U358 : INV_X1 port map( A => n35901, ZN => n3085);
   U359 : OAI22_X1 port map( A1 => n30099, A2 => n36712, B1 => n30843, B2 => 
                           n36572, ZN => n35902);
   U360 : INV_X1 port map( A => n35902, ZN => n3118);
   U361 : OAI22_X1 port map( A1 => n30099, A2 => n36429, B1 => n30844, B2 => 
                           n36572, ZN => n35903);
   U362 : INV_X1 port map( A => n35903, ZN => n3148);
   U363 : OAI22_X1 port map( A1 => n30099, A2 => n36427, B1 => n30845, B2 => 
                           n36572, ZN => n35904);
   U364 : INV_X1 port map( A => n35904, ZN => n3175);
   U365 : OAI22_X1 port map( A1 => n30097, A2 => n36398, B1 => n30847, B2 => 
                           n36609, ZN => n35905);
   U366 : INV_X1 port map( A => n35905, ZN => n3004);
   U367 : OAI22_X1 port map( A1 => n30107, A2 => n36441, B1 => n31019, B2 => 
                           n36525, ZN => n35906);
   U368 : INV_X1 port map( A => n35906, ZN => n3420);
   U369 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31241, ZN => n36515);
   U370 : OAI22_X1 port map( A1 => n30107, A2 => n36515, B1 => n31020, B2 => 
                           n36525, ZN => n35907);
   U371 : INV_X1 port map( A => n35907, ZN => n3325);
   U372 : OAI22_X1 port map( A1 => n30108, A2 => n36327, B1 => n31018, B2 => 
                           n36538, ZN => n35908);
   U373 : INV_X1 port map( A => n35908, ZN => n3453);
   U374 : OAI22_X1 port map( A1 => n30108, A2 => n36515, B1 => n31017, B2 => 
                           n36538, ZN => n35909);
   U375 : INV_X1 port map( A => n35909, ZN => n3324);
   U376 : OAI22_X1 port map( A1 => n30107, A2 => n36469, B1 => n31021, B2 => 
                           n36525, ZN => n35910);
   U377 : INV_X1 port map( A => n35910, ZN => n3388);
   U378 : OAI22_X1 port map( A1 => n30106, A2 => n36515, B1 => n31022, B2 => 
                           n36550, ZN => n35911);
   U379 : INV_X1 port map( A => n35911, ZN => n3326);
   U380 : OAI22_X1 port map( A1 => n30108, A2 => n36425, B1 => n31023, B2 => 
                           n36538, ZN => n35912);
   U381 : INV_X1 port map( A => n35912, ZN => n3516);
   U382 : OAI22_X1 port map( A1 => n30108, A2 => n36677, B1 => n31024, B2 => 
                           n36538, ZN => n35913);
   U383 : INV_X1 port map( A => n35913, ZN => n3052);
   U384 : OAI22_X1 port map( A1 => n30106, A2 => n36327, B1 => n31025, B2 => 
                           n36550, ZN => n35914);
   U385 : INV_X1 port map( A => n35914, ZN => n3454);
   U386 : OAI22_X1 port map( A1 => n30106, A2 => n36677, B1 => n31026, B2 => 
                           n36550, ZN => n35915);
   U387 : INV_X1 port map( A => n35915, ZN => n3053);
   U388 : CLKBUF_X1 port map( A => n36398, Z => n36618);
   U389 : OAI22_X1 port map( A1 => n30108, A2 => n36618, B1 => n31027, B2 => 
                           n36538, ZN => n35916);
   U390 : INV_X1 port map( A => n35916, ZN => n2989);
   U391 : OAI22_X1 port map( A1 => n30106, A2 => n36441, B1 => n31028, B2 => 
                           n36550, ZN => n35917);
   U392 : INV_X1 port map( A => n35917, ZN => n3421);
   U393 : OAI22_X1 port map( A1 => n30107, A2 => n36425, B1 => n31029, B2 => 
                           n36525, ZN => n35918);
   U394 : INV_X1 port map( A => n35918, ZN => n3517);
   U395 : OAI22_X1 port map( A1 => n30108, A2 => n36441, B1 => n31030, B2 => 
                           n36538, ZN => n35919);
   U396 : INV_X1 port map( A => n35919, ZN => n3422);
   U397 : OAI22_X1 port map( A1 => n30107, A2 => n36454, B1 => n31031, B2 => 
                           n36525, ZN => n35920);
   U398 : INV_X1 port map( A => n35920, ZN => n3357);
   U399 : OAI22_X1 port map( A1 => n30106, A2 => n36454, B1 => n31032, B2 => 
                           n36550, ZN => n35921);
   U400 : INV_X1 port map( A => n35921, ZN => n3358);
   U401 : OAI22_X1 port map( A1 => n30106, A2 => n36425, B1 => n31033, B2 => 
                           n36550, ZN => n35922);
   U402 : INV_X1 port map( A => n35922, ZN => n3518);
   U403 : OAI22_X1 port map( A1 => n30108, A2 => n36469, B1 => n31034, B2 => 
                           n36538, ZN => n35923);
   U404 : INV_X1 port map( A => n35923, ZN => n3389);
   U405 : OAI22_X1 port map( A1 => n30108, A2 => n36454, B1 => n31016, B2 => 
                           n36538, ZN => n35924);
   U406 : INV_X1 port map( A => n35924, ZN => n3356);
   U407 : OAI22_X1 port map( A1 => n30107, A2 => n36327, B1 => n31014, B2 => 
                           n36525, ZN => n35925);
   U408 : INV_X1 port map( A => n35925, ZN => n3452);
   U409 : OAI22_X1 port map( A1 => n30106, A2 => n36469, B1 => n31035, B2 => 
                           n36550, ZN => n35926);
   U410 : INV_X1 port map( A => n35926, ZN => n3390);
   U411 : OAI22_X1 port map( A1 => n30097, A2 => n36493, B1 => n31036, B2 => 
                           n36609, ZN => n35927);
   U412 : INV_X1 port map( A => n35927, ZN => n3555);
   U413 : OAI22_X1 port map( A1 => n30108, A2 => n36403, B1 => n31013, B2 => 
                           n36538, ZN => n35928);
   U414 : INV_X1 port map( A => n35928, ZN => n3486);
   U415 : OAI22_X1 port map( A1 => n30093, A2 => n36493, B1 => n31037, B2 => 
                           n36606, ZN => n35929);
   U416 : INV_X1 port map( A => n35929, ZN => n3556);
   U417 : OAI22_X1 port map( A1 => n30103, A2 => n36493, B1 => n31038, B2 => 
                           n36508, ZN => n35930);
   U418 : INV_X1 port map( A => n35930, ZN => n3557);
   U419 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30096, ZN => n36505);
   U420 : OAI22_X1 port map( A1 => n30096, A2 => n36398, B1 => n30849, B2 => 
                           n36505, ZN => n35931);
   U421 : INV_X1 port map( A => n35931, ZN => n3005);
   U422 : OAI22_X1 port map( A1 => n30093, A2 => n36398, B1 => n30852, B2 => 
                           n36606, ZN => n35932);
   U423 : INV_X1 port map( A => n35932, ZN => n3008);
   U424 : OAI22_X1 port map( A1 => n30099, A2 => n36422, B1 => n30855, B2 => 
                           n36572, ZN => n35933);
   U425 : INV_X1 port map( A => n35933, ZN => n3245);
   U426 : OAI22_X1 port map( A1 => n30099, A2 => n36457, B1 => n30856, B2 => 
                           n36572, ZN => n35934);
   U427 : INV_X1 port map( A => n35934, ZN => n3278);
   U428 : OAI22_X1 port map( A1 => n30103, A2 => n36398, B1 => n30858, B2 => 
                           n36508, ZN => n35935);
   U429 : INV_X1 port map( A => n35935, ZN => n3012);
   U430 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n30105, ZN => n36586);
   U431 : OAI22_X1 port map( A1 => n30105, A2 => n36327, B1 => n31047, B2 => 
                           n36586, ZN => n35936);
   U432 : INV_X1 port map( A => n35936, ZN => n3455);
   U433 : OAI22_X1 port map( A1 => n30105, A2 => n36515, B1 => n31048, B2 => 
                           n36586, ZN => n35937);
   U434 : INV_X1 port map( A => n35937, ZN => n3327);
   U435 : OAI22_X1 port map( A1 => n30105, A2 => n36403, B1 => n31049, B2 => 
                           n36586, ZN => n35938);
   U436 : INV_X1 port map( A => n35938, ZN => n3487);
   U437 : OAI22_X1 port map( A1 => n30105, A2 => n36449, B1 => n31050, B2 => 
                           n36586, ZN => n35939);
   U438 : INV_X1 port map( A => n35939, ZN => n3054);
   U439 : OAI22_X1 port map( A1 => n30105, A2 => n36469, B1 => n31051, B2 => 
                           n36586, ZN => n35940);
   U440 : INV_X1 port map( A => n35940, ZN => n3391);
   U441 : OAI22_X1 port map( A1 => n30105, A2 => n36454, B1 => n31052, B2 => 
                           n36586, ZN => n35941);
   U442 : INV_X1 port map( A => n35941, ZN => n3359);
   U443 : CLKBUF_X1 port map( A => n36472, Z => n36584);
   U444 : OAI22_X1 port map( A1 => n30105, A2 => n36584, B1 => n31053, B2 => 
                           n36586, ZN => n35942);
   U445 : INV_X1 port map( A => n35942, ZN => n2893);
   U446 : OAI22_X1 port map( A1 => n30105, A2 => n36398, B1 => n31054, B2 => 
                           n36586, ZN => n35943);
   U447 : INV_X1 port map( A => n35943, ZN => n2990);
   U448 : OAI22_X1 port map( A1 => n30105, A2 => n36441, B1 => n31055, B2 => 
                           n36586, ZN => n35944);
   U449 : INV_X1 port map( A => n35944, ZN => n3423);
   U450 : OAI22_X1 port map( A1 => n30105, A2 => n36425, B1 => n31056, B2 => 
                           n36586, ZN => n35945);
   U451 : INV_X1 port map( A => n35945, ZN => n3519);
   U452 : OAI22_X1 port map( A1 => n30103, A2 => n36403, B1 => n31059, B2 => 
                           n36508, ZN => n35946);
   U453 : INV_X1 port map( A => n35946, ZN => n3488);
   U454 : OAI22_X1 port map( A1 => n30106, A2 => n36618, B1 => n31012, B2 => 
                           n36550, ZN => n35947);
   U455 : INV_X1 port map( A => n35947, ZN => n2988);
   U456 : OAI22_X1 port map( A1 => n30103, A2 => n36515, B1 => n31061, B2 => 
                           n36508, ZN => n35948);
   U457 : INV_X1 port map( A => n35948, ZN => n3329);
   U458 : OAI22_X1 port map( A1 => n30103, A2 => n36469, B1 => n31063, B2 => 
                           n36508, ZN => n35949);
   U459 : INV_X1 port map( A => n35949, ZN => n3393);
   U460 : OAI22_X1 port map( A1 => n30106, A2 => n36584, B1 => n31011, B2 => 
                           n36550, ZN => n35950);
   U461 : INV_X1 port map( A => n35950, ZN => n2891);
   U462 : OAI22_X1 port map( A1 => n30103, A2 => n36327, B1 => n31066, B2 => 
                           n36508, ZN => n35951);
   U463 : INV_X1 port map( A => n35951, ZN => n3456);
   U464 : OAI22_X1 port map( A1 => n30103, A2 => n36454, B1 => n31067, B2 => 
                           n36508, ZN => n35952);
   U465 : INV_X1 port map( A => n35952, ZN => n3361);
   U466 : OAI22_X1 port map( A1 => n30103, A2 => n36425, B1 => n31069, B2 => 
                           n36508, ZN => n35953);
   U467 : INV_X1 port map( A => n35953, ZN => n3521);
   U468 : OAI22_X1 port map( A1 => n30103, A2 => n36441, B1 => n31070, B2 => 
                           n36508, ZN => n35954);
   U469 : INV_X1 port map( A => n35954, ZN => n3425);
   U470 : OAI22_X1 port map( A1 => n30107, A2 => n36677, B1 => n31010, B2 => 
                           n36525, ZN => n35955);
   U471 : INV_X1 port map( A => n35955, ZN => n3051);
   U472 : OAI22_X1 port map( A1 => n30107, A2 => n36618, B1 => n31009, B2 => 
                           n36525, ZN => n35956);
   U473 : INV_X1 port map( A => n35956, ZN => n2987);
   U474 : OAI22_X1 port map( A1 => n30107, A2 => n36403, B1 => n31007, B2 => 
                           n36525, ZN => n35957);
   U475 : INV_X1 port map( A => n35957, ZN => n3485);
   U476 : OAI22_X1 port map( A1 => n30106, A2 => n36403, B1 => n31006, B2 => 
                           n36550, ZN => n35958);
   U477 : INV_X1 port map( A => n35958, ZN => n3484);
   U478 : OAI22_X1 port map( A1 => n30103, A2 => n36683, B1 => n30878, B2 => 
                           n36508, ZN => n35959);
   U479 : INV_X1 port map( A => n35959, ZN => n3041);
   U480 : OAI22_X1 port map( A1 => n30107, A2 => n36662, B1 => n30493, B2 => 
                           n36525, ZN => n35960);
   U481 : INV_X1 port map( A => n35960, ZN => n2974);
   U482 : OAI22_X1 port map( A1 => n30101, A2 => n36683, B1 => n30880, B2 => 
                           n36514, ZN => n35961);
   U483 : INV_X1 port map( A => n35961, ZN => n3043);
   U484 : OAI22_X1 port map( A1 => n30108, A2 => n36457, B1 => n30494, B2 => 
                           n36538, ZN => n35962);
   U485 : INV_X1 port map( A => n35962, ZN => n3293);
   U486 : OAI22_X1 port map( A1 => n30107, A2 => n36674, B1 => n30495, B2 => 
                           n36525, ZN => n35963);
   U487 : INV_X1 port map( A => n35963, ZN => n3262);
   U488 : OAI22_X1 port map( A1 => n30108, A2 => n36748, B1 => n30498, B2 => 
                           n36538, ZN => n35964);
   U489 : INV_X1 port map( A => n35964, ZN => n3101);
   U490 : OAI22_X1 port map( A1 => n30107, A2 => n36457, B1 => n30499, B2 => 
                           n36525, ZN => n35965);
   U491 : INV_X1 port map( A => n35965, ZN => n3294);
   U492 : OAI22_X1 port map( A1 => n30107, A2 => n36748, B1 => n30500, B2 => 
                           n36525, ZN => n35966);
   U493 : INV_X1 port map( A => n35966, ZN => n3102);
   U494 : OAI22_X1 port map( A1 => n30108, A2 => n36783, B1 => n30502, B2 => 
                           n36538, ZN => n35967);
   U495 : INV_X1 port map( A => n35967, ZN => n3165);
   U496 : OAI22_X1 port map( A1 => n30107, A2 => n36783, B1 => n30503, B2 => 
                           n36525, ZN => n35968);
   U497 : INV_X1 port map( A => n35968, ZN => n3166);
   U498 : OAI22_X1 port map( A1 => n30088, A2 => n36515, B1 => n30504, B2 => 
                           n36535, ZN => n35969);
   U499 : INV_X1 port map( A => n35969, ZN => n3310);
   U500 : OAI22_X1 port map( A1 => n30090, A2 => n36515, B1 => n30505, B2 => 
                           n36511, ZN => n35970);
   U501 : INV_X1 port map( A => n35970, ZN => n3311);
   U502 : OAI22_X1 port map( A1 => n30093, A2 => n36579, B1 => n30892, B2 => 
                           n36606, ZN => n35971);
   U503 : INV_X1 port map( A => n35971, ZN => n3018);
   U504 : OAI22_X1 port map( A1 => n30087, A2 => n36515, B1 => n30508, B2 => 
                           n36543, ZN => n35972);
   U505 : INV_X1 port map( A => n35972, ZN => n3314);
   U506 : CLKBUF_X1 port map( A => n36515, Z => n36296);
   U507 : OAI22_X1 port map( A1 => n30089, A2 => n36296, B1 => n30509, B2 => 
                           n36522, ZN => n35973);
   U508 : INV_X1 port map( A => n35973, ZN => n3315);
   U509 : OAI22_X1 port map( A1 => n30089, A2 => n36730, B1 => n30512, B2 => 
                           n36522, ZN => n35974);
   U510 : INV_X1 port map( A => n35974, ZN => n2798);
   U511 : OAI22_X1 port map( A1 => n30089, A2 => n36487, B1 => n30514, B2 => 
                           n36522, ZN => n35975);
   U512 : INV_X1 port map( A => n35975, ZN => n2830);
   U513 : OAI22_X1 port map( A1 => n30108, A2 => n36730, B1 => n30515, B2 => 
                           n36538, ZN => n35976);
   U514 : INV_X1 port map( A => n35976, ZN => n2799);
   U515 : OAI22_X1 port map( A1 => n30108, A2 => n36487, B1 => n30516, B2 => 
                           n36538, ZN => n35977);
   U516 : INV_X1 port map( A => n35977, ZN => n2831);
   U517 : OAI22_X1 port map( A1 => n30107, A2 => n36730, B1 => n30521, B2 => 
                           n36525, ZN => n35978);
   U518 : INV_X1 port map( A => n35978, ZN => n2800);
   U519 : OAI22_X1 port map( A1 => n30107, A2 => n36487, B1 => n30522, B2 => 
                           n36525, ZN => n35979);
   U520 : INV_X1 port map( A => n35979, ZN => n2832);
   U521 : OAI22_X1 port map( A1 => n30106, A2 => n36730, B1 => n30528, B2 => 
                           n36550, ZN => n35980);
   U522 : INV_X1 port map( A => n35980, ZN => n2802);
   U523 : OAI22_X1 port map( A1 => n30106, A2 => n36487, B1 => n30529, B2 => 
                           n36550, ZN => n35981);
   U524 : INV_X1 port map( A => n35981, ZN => n2833);
   U525 : OAI22_X1 port map( A1 => n30088, A2 => n36487, B1 => n30530, B2 => 
                           n36535, ZN => n35982);
   U526 : INV_X1 port map( A => n35982, ZN => n2834);
   U527 : OAI22_X1 port map( A1 => n30088, A2 => n36472, B1 => n30531, B2 => 
                           n36535, ZN => n35983);
   U528 : INV_X1 port map( A => n35983, ZN => n2894);
   U529 : CLKBUF_X1 port map( A => n36487, Z => n36788);
   U530 : OAI22_X1 port map( A1 => n30090, A2 => n36788, B1 => n30542, B2 => 
                           n36511, ZN => n35984);
   U531 : INV_X1 port map( A => n35984, ZN => n2835);
   U532 : OAI22_X1 port map( A1 => n30087, A2 => n36487, B1 => n30543, B2 => 
                           n36543, ZN => n35985);
   U533 : INV_X1 port map( A => n35985, ZN => n2836);
   U534 : OAI22_X1 port map( A1 => n30096, A2 => n36683, B1 => n30907, B2 => 
                           n36505, ZN => n35986);
   U535 : INV_X1 port map( A => n35986, ZN => n3022);
   U536 : OAI22_X1 port map( A1 => n30097, A2 => n36683, B1 => n30908, B2 => 
                           n36609, ZN => n35987);
   U537 : INV_X1 port map( A => n35987, ZN => n3023);
   U538 : OAI22_X1 port map( A1 => n30090, A2 => n36472, B1 => n30544, B2 => 
                           n36511, ZN => n35988);
   U539 : INV_X1 port map( A => n35988, ZN => n2895);
   U540 : OAI22_X1 port map( A1 => n30107, A2 => n36493, B1 => n30910, B2 => 
                           n36525, ZN => n35989);
   U541 : INV_X1 port map( A => n35989, ZN => n3548);
   U542 : OAI22_X1 port map( A1 => n30106, A2 => n36493, B1 => n30911, B2 => 
                           n36550, ZN => n35990);
   U543 : INV_X1 port map( A => n35990, ZN => n3549);
   U544 : OAI22_X1 port map( A1 => n30108, A2 => n36493, B1 => n30912, B2 => 
                           n36538, ZN => n35991);
   U545 : INV_X1 port map( A => n35991, ZN => n3550);
   U546 : OAI22_X1 port map( A1 => n30089, A2 => n36472, B1 => n30556, B2 => 
                           n36522, ZN => n35992);
   U547 : INV_X1 port map( A => n35992, ZN => n2896);
   U548 : OAI22_X1 port map( A1 => n30101, A2 => n36184, B1 => n30917, B2 => 
                           n36514, ZN => n35993);
   U549 : INV_X1 port map( A => n35993, ZN => n3208);
   U550 : OAI22_X1 port map( A1 => n30112, A2 => n36184, B1 => n30918, B2 => 
                           n36519, ZN => n35994);
   U551 : INV_X1 port map( A => n35994, ZN => n3209);
   U552 : OAI22_X1 port map( A1 => n30087, A2 => n36730, B1 => n30565, B2 => 
                           n36543, ZN => n35995);
   U553 : INV_X1 port map( A => n35995, ZN => n2806);
   U554 : OAI22_X1 port map( A1 => n30096, A2 => n36184, B1 => n30921, B2 => 
                           n36505, ZN => n35996);
   U555 : INV_X1 port map( A => n35996, ZN => n3212);
   U556 : OAI22_X1 port map( A1 => n30105, A2 => n36783, B1 => n30579, B2 => 
                           n36586, ZN => n35997);
   U557 : INV_X1 port map( A => n35997, ZN => n3167);
   U558 : OAI22_X1 port map( A1 => n30105, A2 => n36493, B1 => n30924, B2 => 
                           n36586, ZN => n35998);
   U559 : INV_X1 port map( A => n35998, ZN => n3551);
   U560 : OAI22_X1 port map( A1 => n30105, A2 => n36485, B1 => n30580, B2 => 
                           n36586, ZN => n35999);
   U561 : INV_X1 port map( A => n35999, ZN => n3199);
   U562 : OAI22_X1 port map( A1 => n30112, A2 => n36296, B1 => n30926, B2 => 
                           n36519, ZN => n36000);
   U563 : INV_X1 port map( A => n36000, ZN => n3317);
   U564 : OAI22_X1 port map( A1 => n30105, A2 => n36487, B1 => n30583, B2 => 
                           n36586, ZN => n36001);
   U565 : INV_X1 port map( A => n36001, ZN => n2839);
   U566 : OAI22_X1 port map( A1 => n30105, A2 => n36683, B1 => n30586, B2 => 
                           n36586, ZN => n36002);
   U567 : INV_X1 port map( A => n36002, ZN => n3040);
   U568 : OAI22_X1 port map( A1 => n30105, A2 => n36712, B1 => n30587, B2 => 
                           n36586, ZN => n36003);
   U569 : INV_X1 port map( A => n36003, ZN => n3136);
   U570 : OAI22_X1 port map( A1 => n30112, A2 => n36472, B1 => n30930, B2 => 
                           n36519, ZN => n36004);
   U571 : INV_X1 port map( A => n36004, ZN => n2913);
   U572 : OAI22_X1 port map( A1 => n30105, A2 => n36662, B1 => n30588, B2 => 
                           n36586, ZN => n36005);
   U573 : INV_X1 port map( A => n36005, ZN => n2975);
   U574 : OAI22_X1 port map( A1 => n30105, A2 => n36457, B1 => n30590, B2 => 
                           n36586, ZN => n36006);
   U575 : INV_X1 port map( A => n36006, ZN => n3295);
   U576 : OAI22_X1 port map( A1 => n30105, A2 => n36730, B1 => n30591, B2 => 
                           n36586, ZN => n36007);
   U577 : INV_X1 port map( A => n36007, ZN => n2807);
   U578 : OAI22_X1 port map( A1 => n30105, A2 => n36674, B1 => n30592, B2 => 
                           n36586, ZN => n36008);
   U579 : INV_X1 port map( A => n36008, ZN => n3263);
   U580 : OAI22_X1 port map( A1 => n30105, A2 => n36748, B1 => n30594, B2 => 
                           n36586, ZN => n36009);
   U581 : INV_X1 port map( A => n36009, ZN => n3103);
   U582 : OAI22_X1 port map( A1 => n30096, A2 => n36748, B1 => n30595, B2 => 
                           n36505, ZN => n36010);
   U583 : INV_X1 port map( A => n36010, ZN => n3104);
   U584 : OAI22_X1 port map( A1 => n30096, A2 => n36584, B1 => n30597, B2 => 
                           n36505, ZN => n36011);
   U585 : INV_X1 port map( A => n36011, ZN => n2901);
   U586 : OAI22_X1 port map( A1 => n30097, A2 => n36748, B1 => n30598, B2 => 
                           n36609, ZN => n36012);
   U587 : INV_X1 port map( A => n36012, ZN => n3105);
   U588 : OAI22_X1 port map( A1 => n30097, A2 => n36472, B1 => n30602, B2 => 
                           n36609, ZN => n36013);
   U589 : INV_X1 port map( A => n36013, ZN => n2902);
   U590 : OAI22_X1 port map( A1 => n30096, A2 => n36730, B1 => n30604, B2 => 
                           n36505, ZN => n36014);
   U591 : INV_X1 port map( A => n36014, ZN => n2809);
   U592 : OAI22_X1 port map( A1 => n30097, A2 => n36730, B1 => n30605, B2 => 
                           n36609, ZN => n36015);
   U593 : INV_X1 port map( A => n36015, ZN => n2810);
   U594 : OAI22_X1 port map( A1 => n30103, A2 => n36730, B1 => n30942, B2 => 
                           n36508, ZN => n36016);
   U595 : INV_X1 port map( A => n36016, ZN => n2821);
   U596 : OAI22_X1 port map( A1 => n30096, A2 => n36487, B1 => n30606, B2 => 
                           n36505, ZN => n36017);
   U597 : INV_X1 port map( A => n36017, ZN => n2840);
   U598 : CLKBUF_X1 port map( A => n36730, Z => n36751);
   U599 : OAI22_X1 port map( A1 => n30112, A2 => n36751, B1 => n30944, B2 => 
                           n36519, ZN => n36018);
   U600 : INV_X1 port map( A => n36018, ZN => n2790);
   U601 : OAI22_X1 port map( A1 => n30112, A2 => n36487, B1 => n30945, B2 => 
                           n36519, ZN => n36019);
   U602 : INV_X1 port map( A => n36019, ZN => n2853);
   U603 : OAI22_X1 port map( A1 => n30097, A2 => n36487, B1 => n30607, B2 => 
                           n36609, ZN => n36020);
   U604 : INV_X1 port map( A => n36020, ZN => n2841);
   U605 : OAI22_X1 port map( A1 => n30096, A2 => n36662, B1 => n30609, B2 => 
                           n36505, ZN => n36021);
   U606 : INV_X1 port map( A => n36021, ZN => n2976);
   U607 : OAI22_X1 port map( A1 => n30096, A2 => n36457, B1 => n30625, B2 => 
                           n36505, ZN => n36022);
   U608 : INV_X1 port map( A => n36022, ZN => n3296);
   U609 : OAI22_X1 port map( A1 => n30089, A2 => n36683, B1 => n31172, B2 => 
                           n36522, ZN => n36023);
   U610 : INV_X1 port map( A => n36023, ZN => n3024);
   U611 : OAI22_X1 port map( A1 => n30097, A2 => n36457, B1 => n30626, B2 => 
                           n36609, ZN => n36024);
   U612 : INV_X1 port map( A => n36024, ZN => n3297);
   U613 : OAI22_X1 port map( A1 => n30093, A2 => n36748, B1 => n30628, B2 => 
                           n36606, ZN => n36025);
   U614 : INV_X1 port map( A => n36025, ZN => n3108);
   U615 : OAI22_X1 port map( A1 => n30093, A2 => n36457, B1 => n30631, B2 => 
                           n36606, ZN => n36026);
   U616 : INV_X1 port map( A => n36026, ZN => n3301);
   U617 : OAI22_X1 port map( A1 => n30093, A2 => n36662, B1 => n30632, B2 => 
                           n36606, ZN => n36027);
   U618 : INV_X1 port map( A => n36027, ZN => n2981);
   U619 : OAI22_X1 port map( A1 => n30093, A2 => n36472, B1 => n30634, B2 => 
                           n36606, ZN => n36028);
   U620 : INV_X1 port map( A => n36028, ZN => n2905);
   U621 : OAI22_X1 port map( A1 => n30093, A2 => n36487, B1 => n30635, B2 => 
                           n36606, ZN => n36029);
   U622 : INV_X1 port map( A => n36029, ZN => n2845);
   U623 : OAI22_X1 port map( A1 => n30093, A2 => n36674, B1 => n30640, B2 => 
                           n36606, ZN => n36030);
   U624 : INV_X1 port map( A => n36030, ZN => n3267);
   U625 : OAI22_X1 port map( A1 => n30097, A2 => n36449, B1 => n30643, B2 => 
                           n36609, ZN => n36031);
   U626 : INV_X1 port map( A => n36031, ZN => n3068);
   U627 : OAI22_X1 port map( A1 => n30103, A2 => n36788, B1 => n30958, B2 => 
                           n36508, ZN => n36032);
   U628 : INV_X1 port map( A => n36032, ZN => n2829);
   U629 : OAI22_X1 port map( A1 => n30096, A2 => n36296, B1 => n31154, B2 => 
                           n36505, ZN => n36033);
   U630 : INV_X1 port map( A => n36033, ZN => n3309);
   U631 : CLKBUF_X1 port map( A => n36454, Z => n36280);
   U632 : OAI22_X1 port map( A1 => n30093, A2 => n36280, B1 => n31146, B2 => 
                           n36606, ZN => n36034);
   U633 : INV_X1 port map( A => n36034, ZN => n3341);
   U634 : OAI22_X1 port map( A1 => n30096, A2 => n36449, B1 => n30644, B2 => 
                           n36505, ZN => n36035);
   U635 : INV_X1 port map( A => n36035, ZN => n3069);
   U636 : OAI22_X1 port map( A1 => n30099, A2 => n36493, B1 => n30957, B2 => 
                           n36572, ZN => n36036);
   U637 : INV_X1 port map( A => n36036, ZN => n3552);
   U638 : OAI22_X1 port map( A1 => n30097, A2 => n36441, B1 => n31072, B2 => 
                           n36609, ZN => n36037);
   U639 : INV_X1 port map( A => n36037, ZN => n3427);
   U640 : OAI22_X1 port map( A1 => n30099, A2 => n36425, B1 => n31074, B2 => 
                           n36572, ZN => n36038);
   U641 : INV_X1 port map( A => n36038, ZN => n3523);
   U642 : OAI22_X1 port map( A1 => n30097, A2 => n36296, B1 => n31144, B2 => 
                           n36609, ZN => n36039);
   U643 : INV_X1 port map( A => n36039, ZN => n3303);
   U644 : OAI22_X1 port map( A1 => n30093, A2 => n36282, B1 => n31141, B2 => 
                           n36606, ZN => n36040);
   U645 : INV_X1 port map( A => n36040, ZN => n3469);
   U646 : OAI22_X1 port map( A1 => n30097, A2 => n36425, B1 => n31075, B2 => 
                           n36609, ZN => n36041);
   U647 : INV_X1 port map( A => n36041, ZN => n3524);
   U648 : OAI22_X1 port map( A1 => n30096, A2 => n36441, B1 => n31076, B2 => 
                           n36505, ZN => n36042);
   U649 : INV_X1 port map( A => n36042, ZN => n3428);
   U650 : OAI22_X1 port map( A1 => n30096, A2 => n36425, B1 => n31077, B2 => 
                           n36505, ZN => n36043);
   U651 : INV_X1 port map( A => n36043, ZN => n3525);
   U652 : OAI22_X1 port map( A1 => n30097, A2 => n36184, B1 => n30682, B2 => 
                           n36609, ZN => n36044);
   U653 : INV_X1 port map( A => n36044, ZN => n3206);
   U654 : OAI22_X1 port map( A1 => n30093, A2 => n36449, B1 => n30645, B2 => 
                           n36606, ZN => n36045);
   U655 : INV_X1 port map( A => n36045, ZN => n3070);
   U656 : OAI22_X1 port map( A1 => n30099, A2 => n36469, B1 => n31104, B2 => 
                           n36572, ZN => n36046);
   U657 : INV_X1 port map( A => n36046, ZN => n3397);
   U658 : OAI22_X1 port map( A1 => n30093, A2 => n36485, B1 => n30677, B2 => 
                           n36606, ZN => n36047);
   U659 : INV_X1 port map( A => n36047, ZN => n3204);
   U660 : OAI22_X1 port map( A1 => n30099, A2 => n36327, B1 => n31078, B2 => 
                           n36572, ZN => n36048);
   U661 : INV_X1 port map( A => n36048, ZN => n3458);
   U662 : OAI22_X1 port map( A1 => n30097, A2 => n36327, B1 => n31080, B2 => 
                           n36609, ZN => n36049);
   U663 : INV_X1 port map( A => n36049, ZN => n3459);
   U664 : OAI22_X1 port map( A1 => n30096, A2 => n36327, B1 => n31081, B2 => 
                           n36505, ZN => n36050);
   U665 : INV_X1 port map( A => n36050, ZN => n3460);
   U666 : OAI22_X1 port map( A1 => n30093, A2 => n36303, B1 => n31115, B2 => 
                           n36606, ZN => n36051);
   U667 : INV_X1 port map( A => n36051, ZN => n3372);
   U668 : OAI22_X1 port map( A1 => n30103, A2 => n36584, B1 => n30961, B2 => 
                           n36508, ZN => n36052);
   U669 : INV_X1 port map( A => n36052, ZN => n2888);
   U670 : OAI22_X1 port map( A1 => n30099, A2 => n36403, B1 => n31082, B2 => 
                           n36572, ZN => n36053);
   U671 : INV_X1 port map( A => n36053, ZN => n3491);
   U672 : OAI22_X1 port map( A1 => n30101, A2 => n36441, B1 => n31087, B2 => 
                           n36514, ZN => n36054);
   U673 : INV_X1 port map( A => n36054, ZN => n3429);
   U674 : OAI22_X1 port map( A1 => n30096, A2 => n36493, B1 => n30971, B2 => 
                           n36505, ZN => n36055);
   U675 : INV_X1 port map( A => n36055, ZN => n3554);
   U676 : OAI22_X1 port map( A1 => n30101, A2 => n36489, B1 => n31096, B2 => 
                           n36514, ZN => n36056);
   U677 : INV_X1 port map( A => n36056, ZN => n3434);
   U678 : OAI22_X1 port map( A1 => n30101, A2 => n36403, B1 => n31097, B2 => 
                           n36514, ZN => n36057);
   U679 : INV_X1 port map( A => n36057, ZN => n3492);
   U680 : OAI22_X1 port map( A1 => n30096, A2 => n36485, B1 => n30674, B2 => 
                           n36505, ZN => n36058);
   U681 : INV_X1 port map( A => n36058, ZN => n3201);
   U682 : OAI22_X1 port map( A1 => n30101, A2 => n36493, B1 => n30962, B2 => 
                           n36514, ZN => n36059);
   U683 : INV_X1 port map( A => n36059, ZN => n3553);
   U684 : OAI22_X1 port map( A1 => n30093, A2 => n36425, B1 => n31140, B2 => 
                           n36606, ZN => n36060);
   U685 : INV_X1 port map( A => n36060, ZN => n3502);
   U686 : OAI22_X1 port map( A1 => n30097, A2 => n36485, B1 => n30673, B2 => 
                           n36609, ZN => n36061);
   U687 : INV_X1 port map( A => n36061, ZN => n3200);
   U688 : OAI22_X1 port map( A1 => n30101, A2 => n36321, B1 => n31098, B2 => 
                           n36514, ZN => n36062);
   U689 : INV_X1 port map( A => n36062, ZN => n3498);
   U690 : OAI22_X1 port map( A1 => n30096, A2 => n36469, B1 => n31101, B2 => 
                           n36505, ZN => n36063);
   U691 : INV_X1 port map( A => n36063, ZN => n3395);
   U692 : OAI22_X1 port map( A1 => n30093, A2 => n36783, B1 => n30662, B2 => 
                           n36606, ZN => n36064);
   U693 : INV_X1 port map( A => n36064, ZN => n3171);
   U694 : OAI22_X1 port map( A1 => n30093, A2 => n36296, B1 => n31139, B2 => 
                           n36606, ZN => n36065);
   U695 : INV_X1 port map( A => n36065, ZN => n3302);
   U696 : OAI22_X1 port map( A1 => n30096, A2 => n36783, B1 => n30660, B2 => 
                           n36505, ZN => n36066);
   U697 : INV_X1 port map( A => n36066, ZN => n3169);
   U698 : OAI22_X1 port map( A1 => n30097, A2 => n36469, B1 => n31103, B2 => 
                           n36609, ZN => n36067);
   U699 : INV_X1 port map( A => n36067, ZN => n3396);
   U700 : OAI22_X1 port map( A1 => n30093, A2 => n36712, B1 => n30655, B2 => 
                           n36606, ZN => n36068);
   U701 : INV_X1 port map( A => n36068, ZN => n3139);
   U702 : OAI22_X1 port map( A1 => n30096, A2 => n36454, B1 => n31123, B2 => 
                           n36505, ZN => n36069);
   U703 : INV_X1 port map( A => n36069, ZN => n3365);
   U704 : OAI22_X1 port map( A1 => n30101, A2 => n36303, B1 => n31109, B2 => 
                           n36514, ZN => n36070);
   U705 : INV_X1 port map( A => n36070, ZN => n3368);
   U706 : OAI22_X1 port map( A1 => n30097, A2 => n36783, B1 => n30659, B2 => 
                           n36609, ZN => n36071);
   U707 : INV_X1 port map( A => n36071, ZN => n3168);
   U708 : OAI22_X1 port map( A1 => n30097, A2 => n36280, B1 => n31124, B2 => 
                           n36609, ZN => n36072);
   U709 : INV_X1 port map( A => n36072, ZN => n3335);
   U710 : OAI22_X1 port map( A1 => n30099, A2 => n36515, B1 => n31134, B2 => 
                           n36572, ZN => n36073);
   U711 : INV_X1 port map( A => n36073, ZN => n3332);
   U712 : OAI22_X1 port map( A1 => n30096, A2 => n36282, B1 => n31130, B2 => 
                           n36505, ZN => n36074);
   U713 : INV_X1 port map( A => n36074, ZN => n3465);
   U714 : OAI22_X1 port map( A1 => n30093, A2 => n36315, B1 => n31116, B2 => 
                           n36606, ZN => n36075);
   U715 : INV_X1 port map( A => n36075, ZN => n3404);
   U716 : OAI22_X1 port map( A1 => n30097, A2 => n36431, B1 => n30652, B2 => 
                           n36609, ZN => n36076);
   U717 : INV_X1 port map( A => n36076, ZN => n3111);
   U718 : OAI22_X1 port map( A1 => n30093, A2 => n36489, B1 => n31117, B2 => 
                           n36606, ZN => n36077);
   U719 : INV_X1 port map( A => n36077, ZN => n3437);
   U720 : OAI22_X1 port map( A1 => n30101, A2 => n36280, B1 => n31132, B2 => 
                           n36514, ZN => n36078);
   U721 : INV_X1 port map( A => n36078, ZN => n3338);
   U722 : OAI22_X1 port map( A1 => n30099, A2 => n36441, B1 => n31071, B2 => 
                           n36572, ZN => n36079);
   U723 : INV_X1 port map( A => n36079, ZN => n3426);
   U724 : OAI22_X1 port map( A1 => n30096, A2 => n36712, B1 => n30653, B2 => 
                           n36505, ZN => n36080);
   U725 : INV_X1 port map( A => n36080, ZN => n3137);
   U726 : OAI22_X1 port map( A1 => n30097, A2 => n36282, B1 => n31129, B2 => 
                           n36609, ZN => n36081);
   U727 : INV_X1 port map( A => n36081, ZN => n3464);
   U728 : OAI22_X1 port map( A1 => n30099, A2 => n36280, B1 => n31128, B2 => 
                           n36572, ZN => n36082);
   U729 : INV_X1 port map( A => n36082, ZN => n3336);
   U730 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30109, ZN => n36726);
   U731 : OAI22_X1 port map( A1 => n30109, A2 => n36683, B1 => n30316, B2 => 
                           n36726, ZN => n36083);
   U732 : INV_X1 port map( A => n36083, ZN => n3036);
   U733 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30116, ZN => n36717);
   U734 : OAI22_X1 port map( A1 => n30116, A2 => n36683, B1 => n30312, B2 => 
                           n36717, ZN => n36084);
   U735 : INV_X1 port map( A => n36084, ZN => n3033);
   U736 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30117, ZN => n36708);
   U737 : OAI22_X1 port map( A1 => n30117, A2 => n36683, B1 => n30311, B2 => 
                           n36708, ZN => n36085);
   U738 : INV_X1 port map( A => n36085, ZN => n3032);
   U739 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30120, ZN => n36705);
   U740 : OAI22_X1 port map( A1 => n30120, A2 => n36683, B1 => n30310, B2 => 
                           n36705, ZN => n36086);
   U741 : INV_X1 port map( A => n36086, ZN => n3031);
   U742 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30123, ZN => n36703);
   U743 : OAI22_X1 port map( A1 => n30123, A2 => n36683, B1 => n30309, B2 => 
                           n36703, ZN => n36087);
   U744 : INV_X1 port map( A => n36087, ZN => n3030);
   U745 : OAI22_X1 port map( A1 => n30116, A2 => n36485, B1 => n30307, B2 => 
                           n36717, ZN => n36088);
   U746 : INV_X1 port map( A => n36088, ZN => n3193);
   U747 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30124, ZN => n36714);
   U748 : OAI22_X1 port map( A1 => n30124, A2 => n36718, B1 => n30306, B2 => 
                           n36714, ZN => n36089);
   U749 : INV_X1 port map( A => n36089, ZN => n2933);
   U750 : OAI22_X1 port map( A1 => n30117, A2 => n36485, B1 => n30305, B2 => 
                           n36708, ZN => n36090);
   U751 : INV_X1 port map( A => n36090, ZN => n3192);
   U752 : OAI22_X1 port map( A1 => n30120, A2 => n36485, B1 => n30304, B2 => 
                           n36705, ZN => n36091);
   U753 : INV_X1 port map( A => n36091, ZN => n3191);
   U754 : OAI22_X1 port map( A1 => n30123, A2 => n36427, B1 => n30303, B2 => 
                           n36703, ZN => n36092);
   U755 : INV_X1 port map( A => n36092, ZN => n3190);
   U756 : OAI22_X1 port map( A1 => n30124, A2 => n36485, B1 => n30302, B2 => 
                           n36714, ZN => n36093);
   U757 : INV_X1 port map( A => n36093, ZN => n3189);
   U758 : OAI22_X1 port map( A1 => n30109, A2 => n36427, B1 => n30301, B2 => 
                           n36726, ZN => n36094);
   U759 : INV_X1 port map( A => n36094, ZN => n3188);
   U760 : OAI22_X1 port map( A1 => n30124, A2 => n36618, B1 => n30299, B2 => 
                           n36714, ZN => n36095);
   U761 : INV_X1 port map( A => n36095, ZN => n2997);
   U762 : OAI22_X1 port map( A1 => n30116, A2 => n36783, B1 => n30297, B2 => 
                           n36717, ZN => n36096);
   U763 : INV_X1 port map( A => n36096, ZN => n3162);
   U764 : OAI22_X1 port map( A1 => n30117, A2 => n36783, B1 => n30296, B2 => 
                           n36708, ZN => n36097);
   U765 : INV_X1 port map( A => n36097, ZN => n3161);
   U766 : OAI22_X1 port map( A1 => n30120, A2 => n36783, B1 => n30295, B2 => 
                           n36705, ZN => n36098);
   U767 : INV_X1 port map( A => n36098, ZN => n3160);
   U768 : OAI22_X1 port map( A1 => n30124, A2 => n36783, B1 => n30293, B2 => 
                           n36714, ZN => n36099);
   U769 : INV_X1 port map( A => n36099, ZN => n3158);
   U770 : OAI22_X1 port map( A1 => n30124, A2 => n36662, B1 => n30291, B2 => 
                           n36714, ZN => n36100);
   U771 : INV_X1 port map( A => n36100, ZN => n2965);
   U772 : OAI22_X1 port map( A1 => n30109, A2 => n36429, B1 => n30290, B2 => 
                           n36726, ZN => n36101);
   U773 : INV_X1 port map( A => n36101, ZN => n3157);
   U774 : OAI22_X1 port map( A1 => n30116, A2 => n36712, B1 => n30288, B2 => 
                           n36717, ZN => n36102);
   U775 : INV_X1 port map( A => n36102, ZN => n3133);
   U776 : OAI22_X1 port map( A1 => n30120, A2 => n36712, B1 => n30286, B2 => 
                           n36705, ZN => n36103);
   U777 : INV_X1 port map( A => n36103, ZN => n3131);
   U778 : OAI22_X1 port map( A1 => n30123, A2 => n36712, B1 => n30285, B2 => 
                           n36703, ZN => n36104);
   U779 : INV_X1 port map( A => n36104, ZN => n3130);
   U780 : OAI22_X1 port map( A1 => n30124, A2 => n36712, B1 => n30284, B2 => 
                           n36714, ZN => n36105);
   U781 : INV_X1 port map( A => n36105, ZN => n3129);
   U782 : OAI22_X1 port map( A1 => n30109, A2 => n36712, B1 => n30280, B2 => 
                           n36726, ZN => n36106);
   U783 : INV_X1 port map( A => n36106, ZN => n3128);
   U784 : OAI22_X1 port map( A1 => n30117, A2 => n36748, B1 => n30271, B2 => 
                           n36708, ZN => n36107);
   U785 : INV_X1 port map( A => n36107, ZN => n3098);
   U786 : OAI22_X1 port map( A1 => n30116, A2 => n36433, B1 => n30270, B2 => 
                           n36717, ZN => n36108);
   U787 : INV_X1 port map( A => n36108, ZN => n3078);
   U788 : OAI22_X1 port map( A1 => n30124, A2 => n36677, B1 => n30268, B2 => 
                           n36714, ZN => n36109);
   U789 : INV_X1 port map( A => n36109, ZN => n3061);
   U790 : OAI22_X1 port map( A1 => n30123, A2 => n36748, B1 => n30265, B2 => 
                           n36703, ZN => n36110);
   U791 : INV_X1 port map( A => n36110, ZN => n3094);
   U792 : OAI22_X1 port map( A1 => n30120, A2 => n36433, B1 => n30264, B2 => 
                           n36705, ZN => n36111);
   U793 : INV_X1 port map( A => n36111, ZN => n3093);
   U794 : OAI22_X1 port map( A1 => n30117, A2 => n36420, B1 => n30252, B2 => 
                           n36708, ZN => n36112);
   U795 : INV_X1 port map( A => n36112, ZN => n3270);
   U796 : OAI22_X1 port map( A1 => n30123, A2 => n36457, B1 => n30251, B2 => 
                           n36703, ZN => n36113);
   U797 : INV_X1 port map( A => n36113, ZN => n3289);
   U798 : OAI22_X1 port map( A1 => n30124, A2 => n36457, B1 => n30250, B2 => 
                           n36714, ZN => n36114);
   U799 : INV_X1 port map( A => n36114, ZN => n3288);
   U800 : OAI22_X1 port map( A1 => n30120, A2 => n36457, B1 => n30249, B2 => 
                           n36705, ZN => n36115);
   U801 : INV_X1 port map( A => n36115, ZN => n3287);
   U802 : OAI22_X1 port map( A1 => n30116, A2 => n36420, B1 => n30248, B2 => 
                           n36717, ZN => n36116);
   U803 : INV_X1 port map( A => n36116, ZN => n3286);
   U804 : OAI22_X1 port map( A1 => n30109, A2 => n36457, B1 => n30247, B2 => 
                           n36726, ZN => n36117);
   U805 : INV_X1 port map( A => n36117, ZN => n3285);
   U806 : OAI22_X1 port map( A1 => n30109, A2 => n36674, B1 => n30238, B2 => 
                           n36726, ZN => n36118);
   U807 : INV_X1 port map( A => n36118, ZN => n3258);
   U808 : OAI22_X1 port map( A1 => n30123, A2 => n36674, B1 => n30236, B2 => 
                           n36703, ZN => n36119);
   U809 : INV_X1 port map( A => n36119, ZN => n3256);
   U810 : OAI22_X1 port map( A1 => n30116, A2 => n36674, B1 => n30235, B2 => 
                           n36717, ZN => n36120);
   U811 : INV_X1 port map( A => n36120, ZN => n3255);
   U812 : OAI22_X1 port map( A1 => n30120, A2 => n36674, B1 => n30234, B2 => 
                           n36705, ZN => n36121);
   U813 : INV_X1 port map( A => n36121, ZN => n3254);
   U814 : OAI22_X1 port map( A1 => n30117, A2 => n36422, B1 => n30233, B2 => 
                           n36708, ZN => n36122);
   U815 : INV_X1 port map( A => n36122, ZN => n3253);
   U816 : OAI22_X1 port map( A1 => n30124, A2 => n36674, B1 => n30232, B2 => 
                           n36714, ZN => n36123);
   U817 : INV_X1 port map( A => n36123, ZN => n3252);
   U818 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30085, ZN => n36710);
   U819 : OAI22_X1 port map( A1 => n30085, A2 => n36420, B1 => n30224, B2 => 
                           n36710, ZN => n36124);
   U820 : INV_X1 port map( A => n36124, ZN => n3284);
   U821 : OAI22_X1 port map( A1 => n30085, A2 => n36422, B1 => n30222, B2 => 
                           n36710, ZN => n36125);
   U822 : INV_X1 port map( A => n36125, ZN => n3251);
   U823 : OAI22_X1 port map( A1 => n30085, A2 => n36485, B1 => n30221, B2 => 
                           n36710, ZN => n36126);
   U824 : INV_X1 port map( A => n36126, ZN => n3186);
   U825 : OAI22_X1 port map( A1 => n30085, A2 => n36712, B1 => n30214, B2 => 
                           n36710, ZN => n36127);
   U826 : INV_X1 port map( A => n36127, ZN => n3124);
   U827 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30086, ZN => n36736);
   U828 : OAI22_X1 port map( A1 => n30086, A2 => n36477, B1 => n30206, B2 => 
                           n36736, ZN => n36128);
   U829 : INV_X1 port map( A => n36128, ZN => n2867);
   U830 : OAI22_X1 port map( A1 => n30086, A2 => n36701, B1 => n30200, B2 => 
                           n36736, ZN => n36129);
   U831 : INV_X1 port map( A => n36129, ZN => n2931);
   U832 : OAI22_X1 port map( A1 => n30086, A2 => n36692, B1 => n30198, B2 => 
                           n36736, ZN => n36130);
   U833 : INV_X1 port map( A => n36130, ZN => n2963);
   U834 : OAI22_X1 port map( A1 => n30085, A2 => n36579, B1 => n30197, B2 => 
                           n36710, ZN => n36131);
   U835 : INV_X1 port map( A => n36131, ZN => n3027);
   U836 : OAI22_X1 port map( A1 => n30086, A2 => n36618, B1 => n30196, B2 => 
                           n36736, ZN => n36132);
   U837 : INV_X1 port map( A => n36132, ZN => n2995);
   U838 : OAI22_X1 port map( A1 => n30086, A2 => n36683, B1 => n30195, B2 => 
                           n36736, ZN => n36133);
   U839 : INV_X1 port map( A => n36133, ZN => n3026);
   U840 : OAI22_X1 port map( A1 => n30086, A2 => n36449, B1 => n30194, B2 => 
                           n36736, ZN => n36134);
   U841 : INV_X1 port map( A => n36134, ZN => n3058);
   U842 : OAI22_X1 port map( A1 => n30086, A2 => n36748, B1 => n30186, B2 => 
                           n36736, ZN => n36135);
   U843 : INV_X1 port map( A => n36135, ZN => n3090);
   U844 : OAI22_X1 port map( A1 => n30086, A2 => n36712, B1 => n30185, B2 => 
                           n36736, ZN => n36136);
   U845 : INV_X1 port map( A => n36136, ZN => n3122);
   U846 : OAI22_X1 port map( A1 => n30086, A2 => n36485, B1 => n30182, B2 => 
                           n36736, ZN => n36137);
   U847 : INV_X1 port map( A => n36137, ZN => n3184);
   U848 : OAI22_X1 port map( A1 => n30086, A2 => n36674, B1 => n30180, B2 => 
                           n36736, ZN => n36138);
   U849 : INV_X1 port map( A => n36138, ZN => n3248);
   U850 : OAI22_X1 port map( A1 => n30086, A2 => n36457, B1 => n30179, B2 => 
                           n36736, ZN => n36139);
   U851 : INV_X1 port map( A => n36139, ZN => n3280);
   U852 : OAI22_X1 port map( A1 => n30085, A2 => n36715, B1 => n30154, B2 => 
                           n36710, ZN => n36140);
   U853 : INV_X1 port map( A => n36140, ZN => n2863);
   U854 : OAI22_X1 port map( A1 => n30085, A2 => n36718, B1 => n30152, B2 => 
                           n36710, ZN => n36141);
   U855 : INV_X1 port map( A => n36141, ZN => n2927);
   U856 : OAI22_X1 port map( A1 => n30085, A2 => n36662, B1 => n30149, B2 => 
                           n36710, ZN => n36142);
   U857 : INV_X1 port map( A => n36142, ZN => n2959);
   U858 : OAI22_X1 port map( A1 => n30085, A2 => n36398, B1 => n30147, B2 => 
                           n36710, ZN => n36143);
   U859 : INV_X1 port map( A => n36143, ZN => n2991);
   U860 : OAI22_X1 port map( A1 => n30085, A2 => n36449, B1 => n30146, B2 => 
                           n36710, ZN => n36144);
   U861 : INV_X1 port map( A => n36144, ZN => n3055);
   U862 : OAI22_X1 port map( A1 => n30116, A2 => n36751, B1 => n30947, B2 => 
                           n36717, ZN => n36145);
   U863 : INV_X1 port map( A => n36145, ZN => n2792);
   U864 : OAI22_X1 port map( A1 => n30109, A2 => n36487, B1 => n30943, B2 => 
                           n36726, ZN => n36146);
   U865 : INV_X1 port map( A => n36146, ZN => n2852);
   U866 : OAI22_X1 port map( A1 => n30120, A2 => n36584, B1 => n30940, B2 => 
                           n36705, ZN => n36147);
   U867 : INV_X1 port map( A => n36147, ZN => n2887);
   U868 : OAI22_X1 port map( A1 => n30124, A2 => n36515, B1 => n30939, B2 => 
                           n36714, ZN => n36148);
   U869 : INV_X1 port map( A => n36148, ZN => n3323);
   U870 : OAI22_X1 port map( A1 => n30117, A2 => n36788, B1 => n30952, B2 => 
                           n36708, ZN => n36149);
   U871 : INV_X1 port map( A => n36149, ZN => n2824);
   U872 : OAI22_X1 port map( A1 => n30124, A2 => n36584, B1 => n30938, B2 => 
                           n36714, ZN => n36150);
   U873 : INV_X1 port map( A => n36150, ZN => n2886);
   U874 : OAI22_X1 port map( A1 => n30117, A2 => n36472, B1 => n30937, B2 => 
                           n36708, ZN => n36151);
   U875 : INV_X1 port map( A => n36151, ZN => n2917);
   U876 : OAI22_X1 port map( A1 => n30117, A2 => n36515, B1 => n30936, B2 => 
                           n36708, ZN => n36152);
   U877 : INV_X1 port map( A => n36152, ZN => n3322);
   U878 : OAI22_X1 port map( A1 => n30120, A2 => n36515, B1 => n30935, B2 => 
                           n36705, ZN => n36153);
   U879 : INV_X1 port map( A => n36153, ZN => n3321);
   U880 : OAI22_X1 port map( A1 => n30123, A2 => n36788, B1 => n30954, B2 => 
                           n36703, ZN => n36154);
   U881 : INV_X1 port map( A => n36154, ZN => n2826);
   U882 : OAI22_X1 port map( A1 => n30123, A2 => n36472, B1 => n30932, B2 => 
                           n36703, ZN => n36155);
   U883 : INV_X1 port map( A => n36155, ZN => n2915);
   U884 : OAI22_X1 port map( A1 => n30109, A2 => n36472, B1 => n30931, B2 => 
                           n36726, ZN => n36156);
   U885 : INV_X1 port map( A => n36156, ZN => n2914);
   U886 : OAI22_X1 port map( A1 => n30116, A2 => n36472, B1 => n30929, B2 => 
                           n36717, ZN => n36157);
   U887 : INV_X1 port map( A => n36157, ZN => n2912);
   U888 : OAI22_X1 port map( A1 => n30085, A2 => n36643, B1 => n30455, B2 => 
                           n36710, ZN => n36158);
   U889 : INV_X1 port map( A => n36158, ZN => n3217);
   U890 : OAI22_X1 port map( A1 => n30086, A2 => n36643, B1 => n30454, B2 => 
                           n36736, ZN => n36159);
   U891 : INV_X1 port map( A => n36159, ZN => n3216);
   U892 : OAI22_X1 port map( A1 => n30123, A2 => n36515, B1 => n30928, B2 => 
                           n36703, ZN => n36160);
   U893 : INV_X1 port map( A => n36160, ZN => n3319);
   U894 : OAI22_X1 port map( A1 => n30086, A2 => n36280, B1 => n30436, B2 => 
                           n36736, ZN => n36161);
   U895 : INV_X1 port map( A => n36161, ZN => n3334);
   U896 : OAI22_X1 port map( A1 => n30109, A2 => n36515, B1 => n30927, B2 => 
                           n36726, ZN => n36162);
   U897 : INV_X1 port map( A => n36162, ZN => n3318);
   U898 : OAI22_X1 port map( A1 => n30086, A2 => n36469, B1 => n30435, B2 => 
                           n36736, ZN => n36163);
   U899 : INV_X1 port map( A => n36163, ZN => n3385);
   U900 : OAI22_X1 port map( A1 => n30086, A2 => n36441, B1 => n30434, B2 => 
                           n36736, ZN => n36164);
   U901 : INV_X1 port map( A => n36164, ZN => n3416);
   U902 : OAI22_X1 port map( A1 => n30086, A2 => n36327, B1 => n30432, B2 => 
                           n36736, ZN => n36165);
   U903 : INV_X1 port map( A => n36165, ZN => n3449);
   U904 : OAI22_X1 port map( A1 => n30086, A2 => n36403, B1 => n30429, B2 => 
                           n36736, ZN => n36166);
   U905 : INV_X1 port map( A => n36166, ZN => n3480);
   U906 : OAI22_X1 port map( A1 => n30085, A2 => n36425, B1 => n30426, B2 => 
                           n36710, ZN => n36167);
   U907 : INV_X1 port map( A => n36167, ZN => n3513);
   U908 : OAI22_X1 port map( A1 => n30085, A2 => n36403, B1 => n30424, B2 => 
                           n36710, ZN => n36168);
   U909 : INV_X1 port map( A => n36168, ZN => n3479);
   U910 : OAI22_X1 port map( A1 => n30085, A2 => n36327, B1 => n30423, B2 => 
                           n36710, ZN => n36169);
   U911 : INV_X1 port map( A => n36169, ZN => n3448);
   U912 : OAI22_X1 port map( A1 => n30085, A2 => n36441, B1 => n30422, B2 => 
                           n36710, ZN => n36170);
   U913 : INV_X1 port map( A => n36170, ZN => n3415);
   U914 : OAI22_X1 port map( A1 => n30085, A2 => n36469, B1 => n30421, B2 => 
                           n36710, ZN => n36171);
   U915 : INV_X1 port map( A => n36171, ZN => n3384);
   U916 : OAI22_X1 port map( A1 => n30086, A2 => n36425, B1 => n30419, B2 => 
                           n36736, ZN => n36172);
   U917 : INV_X1 port map( A => n36172, ZN => n3511);
   U918 : OAI22_X1 port map( A1 => n30116, A2 => n36515, B1 => n30925, B2 => 
                           n36717, ZN => n36173);
   U919 : INV_X1 port map( A => n36173, ZN => n3316);
   U920 : OAI22_X1 port map( A1 => n30085, A2 => n36454, B1 => n30418, B2 => 
                           n36710, ZN => n36174);
   U921 : INV_X1 port map( A => n36174, ZN => n3351);
   U922 : OAI22_X1 port map( A1 => n30123, A2 => n36643, B1 => n30923, B2 => 
                           n36703, ZN => n36175);
   U923 : INV_X1 port map( A => n36175, ZN => n3214);
   U924 : OAI22_X1 port map( A1 => n30109, A2 => n36493, B1 => n30416, B2 => 
                           n36726, ZN => n36176);
   U925 : INV_X1 port map( A => n36176, ZN => n3547);
   U926 : OAI22_X1 port map( A1 => n30116, A2 => n36493, B1 => n30415, B2 => 
                           n36717, ZN => n36177);
   U927 : INV_X1 port map( A => n36177, ZN => n3546);
   U928 : OAI22_X1 port map( A1 => n30124, A2 => n36184, B1 => n30922, B2 => 
                           n36714, ZN => n36178);
   U929 : INV_X1 port map( A => n36178, ZN => n3213);
   U930 : OAI22_X1 port map( A1 => n30123, A2 => n36493, B1 => n30412, B2 => 
                           n36703, ZN => n36179);
   U931 : INV_X1 port map( A => n36179, ZN => n3544);
   U932 : OAI22_X1 port map( A1 => n30120, A2 => n36184, B1 => n30920, B2 => 
                           n36705, ZN => n36180);
   U933 : INV_X1 port map( A => n36180, ZN => n3211);
   U934 : OAI22_X1 port map( A1 => n30124, A2 => n36493, B1 => n30411, B2 => 
                           n36714, ZN => n36181);
   U935 : INV_X1 port map( A => n36181, ZN => n3543);
   U936 : OAI22_X1 port map( A1 => n30116, A2 => n36184, B1 => n30919, B2 => 
                           n36717, ZN => n36182);
   U937 : INV_X1 port map( A => n36182, ZN => n3210);
   U938 : OAI22_X1 port map( A1 => n30120, A2 => n36493, B1 => n30409, B2 => 
                           n36705, ZN => n36183);
   U939 : INV_X1 port map( A => n36183, ZN => n3541);
   U940 : OAI22_X1 port map( A1 => n30117, A2 => n36184, B1 => n30916, B2 => 
                           n36708, ZN => n36185);
   U941 : INV_X1 port map( A => n36185, ZN => n3207);
   U942 : OAI22_X1 port map( A1 => n30120, A2 => n36398, B1 => n30407, B2 => 
                           n36705, ZN => n36186);
   U943 : INV_X1 port map( A => n36186, ZN => n3002);
   U944 : OAI22_X1 port map( A1 => n30123, A2 => n36618, B1 => n30406, B2 => 
                           n36703, ZN => n36187);
   U945 : INV_X1 port map( A => n36187, ZN => n2982);
   U946 : OAI22_X1 port map( A1 => n30109, A2 => n36643, B1 => n30915, B2 => 
                           n36726, ZN => n36188);
   U947 : INV_X1 port map( A => n36188, ZN => n3237);
   U948 : OAI22_X1 port map( A1 => n30086, A2 => n36515, B1 => n30506, B2 => 
                           n36736, ZN => n36189);
   U949 : INV_X1 port map( A => n36189, ZN => n3312);
   U950 : OAI22_X1 port map( A1 => n30085, A2 => n36515, B1 => n30507, B2 => 
                           n36710, ZN => n36190);
   U951 : INV_X1 port map( A => n36190, ZN => n3313);
   U952 : OAI22_X1 port map( A1 => n30124, A2 => n36425, B1 => n30405, B2 => 
                           n36714, ZN => n36191);
   U953 : INV_X1 port map( A => n36191, ZN => n3510);
   U954 : OAI22_X1 port map( A1 => n30109, A2 => n36398, B1 => n30404, B2 => 
                           n36726, ZN => n36192);
   U955 : INV_X1 port map( A => n36192, ZN => n3001);
   U956 : OAI22_X1 port map( A1 => n30124, A2 => n36683, B1 => n30403, B2 => 
                           n36714, ZN => n36193);
   U957 : INV_X1 port map( A => n36193, ZN => n3037);
   U958 : OAI22_X1 port map( A1 => n30117, A2 => n36441, B1 => n30401, B2 => 
                           n36708, ZN => n36194);
   U959 : INV_X1 port map( A => n36194, ZN => n3414);
   U960 : OAI22_X1 port map( A1 => n30116, A2 => n36398, B1 => n30400, B2 => 
                           n36717, ZN => n36195);
   U961 : INV_X1 port map( A => n36195, ZN => n2999);
   U962 : OAI22_X1 port map( A1 => n30109, A2 => n36425, B1 => n30399, B2 => 
                           n36726, ZN => n36196);
   U963 : INV_X1 port map( A => n36196, ZN => n3509);
   U964 : OAI22_X1 port map( A1 => n30117, A2 => n36398, B1 => n30398, B2 => 
                           n36708, ZN => n36197);
   U965 : INV_X1 port map( A => n36197, ZN => n2998);
   U966 : OAI22_X1 port map( A1 => n30109, A2 => n36441, B1 => n30397, B2 => 
                           n36726, ZN => n36198);
   U967 : INV_X1 port map( A => n36198, ZN => n3413);
   U968 : OAI22_X1 port map( A1 => n30124, A2 => n36788, B1 => n30955, B2 => 
                           n36714, ZN => n36199);
   U969 : INV_X1 port map( A => n36199, ZN => n2827);
   U970 : OAI22_X1 port map( A1 => n30116, A2 => n36403, B1 => n30395, B2 => 
                           n36717, ZN => n36200);
   U971 : INV_X1 port map( A => n36200, ZN => n3477);
   U972 : OAI22_X1 port map( A1 => n30124, A2 => n36748, B1 => n30394, B2 => 
                           n36714, ZN => n36201);
   U973 : INV_X1 port map( A => n36201, ZN => n3099);
   U974 : OAI22_X1 port map( A1 => n30117, A2 => n36282, B1 => n30393, B2 => 
                           n36708, ZN => n36202);
   U975 : INV_X1 port map( A => n36202, ZN => n3476);
   U976 : OAI22_X1 port map( A1 => n30123, A2 => n36321, B1 => n30392, B2 => 
                           n36703, ZN => n36203);
   U977 : INV_X1 port map( A => n36203, ZN => n3508);
   U978 : OAI22_X1 port map( A1 => n30120, A2 => n36321, B1 => n30391, B2 => 
                           n36705, ZN => n36204);
   U979 : INV_X1 port map( A => n36204, ZN => n3507);
   U980 : OAI22_X1 port map( A1 => n30117, A2 => n36425, B1 => n30390, B2 => 
                           n36708, ZN => n36205);
   U981 : INV_X1 port map( A => n36205, ZN => n3506);
   U982 : OAI22_X1 port map( A1 => n30116, A2 => n36425, B1 => n30389, B2 => 
                           n36717, ZN => n36206);
   U983 : INV_X1 port map( A => n36206, ZN => n3505);
   U984 : OAI22_X1 port map( A1 => n30124, A2 => n36454, B1 => n30388, B2 => 
                           n36714, ZN => n36207);
   U985 : INV_X1 port map( A => n36207, ZN => n3350);
   U986 : OAI22_X1 port map( A1 => n30116, A2 => n36315, B1 => n30387, B2 => 
                           n36717, ZN => n36208);
   U987 : INV_X1 port map( A => n36208, ZN => n3412);
   U988 : OAI22_X1 port map( A1 => n30124, A2 => n36327, B1 => n30385, B2 => 
                           n36714, ZN => n36209);
   U989 : INV_X1 port map( A => n36209, ZN => n3446);
   U990 : OAI22_X1 port map( A1 => n30124, A2 => n36282, B1 => n30384, B2 => 
                           n36714, ZN => n36210);
   U991 : INV_X1 port map( A => n36210, ZN => n3475);
   U992 : OAI22_X1 port map( A1 => n30120, A2 => n36403, B1 => n30383, B2 => 
                           n36705, ZN => n36211);
   U993 : INV_X1 port map( A => n36211, ZN => n3474);
   U994 : OAI22_X1 port map( A1 => n30123, A2 => n36315, B1 => n30381, B2 => 
                           n36703, ZN => n36212);
   U995 : INV_X1 port map( A => n36212, ZN => n3411);
   U996 : OAI22_X1 port map( A1 => n30120, A2 => n36441, B1 => n30380, B2 => 
                           n36705, ZN => n36213);
   U997 : INV_X1 port map( A => n36213, ZN => n3410);
   U998 : OAI22_X1 port map( A1 => n30116, A2 => n36327, B1 => n30379, B2 => 
                           n36717, ZN => n36214);
   U999 : INV_X1 port map( A => n36214, ZN => n3445);
   U1000 : OAI22_X1 port map( A1 => n30109, A2 => n36327, B1 => n30376, B2 => 
                           n36726, ZN => n36215);
   U1001 : INV_X1 port map( A => n36215, ZN => n3442);
   U1002 : OAI22_X1 port map( A1 => n30123, A2 => n36403, B1 => n30375, B2 => 
                           n36703, ZN => n36216);
   U1003 : INV_X1 port map( A => n36216, ZN => n3473);
   U1004 : OAI22_X1 port map( A1 => n30120, A2 => n36751, B1 => n30965, B2 => 
                           n36705, ZN => n36217);
   U1005 : INV_X1 port map( A => n36217, ZN => n2796);
   U1006 : OAI22_X1 port map( A1 => n30124, A2 => n36441, B1 => n30374, B2 => 
                           n36714, ZN => n36218);
   U1007 : INV_X1 port map( A => n36218, ZN => n3409);
   U1008 : OAI22_X1 port map( A1 => n30123, A2 => n36449, B1 => n30373, B2 => 
                           n36703, ZN => n36219);
   U1009 : INV_X1 port map( A => n36219, ZN => n3067);
   U1010 : OAI22_X1 port map( A1 => n30109, A2 => n36403, B1 => n30372, B2 => 
                           n36726, ZN => n36220);
   U1011 : INV_X1 port map( A => n36220, ZN => n3472);
   U1012 : OAI22_X1 port map( A1 => n30123, A2 => n36327, B1 => n30368, B2 => 
                           n36703, ZN => n36221);
   U1013 : INV_X1 port map( A => n36221, ZN => n3441);
   U1014 : OAI22_X1 port map( A1 => n30123, A2 => n36454, B1 => n30367, B2 => 
                           n36703, ZN => n36222);
   U1015 : INV_X1 port map( A => n36222, ZN => n3349);
   U1016 : OAI22_X1 port map( A1 => n30123, A2 => n36469, B1 => n30366, B2 => 
                           n36703, ZN => n36223);
   U1017 : INV_X1 port map( A => n36223, ZN => n3382);
   U1018 : OAI22_X1 port map( A1 => n30120, A2 => n36327, B1 => n30365, B2 => 
                           n36705, ZN => n36224);
   U1019 : INV_X1 port map( A => n36224, ZN => n3440);
   U1020 : OAI22_X1 port map( A1 => n30117, A2 => n36493, B1 => n30413, B2 => 
                           n36708, ZN => n36225);
   U1021 : INV_X1 port map( A => n36225, ZN => n3545);
   U1022 : OAI22_X1 port map( A1 => n30086, A2 => n36493, B1 => n30340, B2 => 
                           n36736, ZN => n36226);
   U1023 : INV_X1 port map( A => n36226, ZN => n3536);
   U1024 : OAI22_X1 port map( A1 => n30117, A2 => n36327, B1 => n30364, B2 => 
                           n36708, ZN => n36227);
   U1025 : INV_X1 port map( A => n36227, ZN => n3439);
   U1026 : OAI22_X1 port map( A1 => n30117, A2 => n36469, B1 => n30348, B2 => 
                           n36708, ZN => n36228);
   U1027 : INV_X1 port map( A => n36228, ZN => n3378);
   U1028 : OAI22_X1 port map( A1 => n30109, A2 => n36449, B1 => n30356, B2 => 
                           n36726, ZN => n36229);
   U1029 : INV_X1 port map( A => n36229, ZN => n3063);
   U1030 : OAI22_X1 port map( A1 => n30109, A2 => n36715, B1 => n30326, B2 => 
                           n36726, ZN => n36230);
   U1031 : INV_X1 port map( A => n36230, ZN => n2875);
   U1032 : OAI22_X1 port map( A1 => n30123, A2 => n36718, B1 => n30318, B2 => 
                           n36703, ZN => n36231);
   U1033 : INV_X1 port map( A => n36231, ZN => n2934);
   U1034 : OAI22_X1 port map( A1 => n30120, A2 => n36662, B1 => n30328, B2 => 
                           n36705, ZN => n36232);
   U1035 : INV_X1 port map( A => n36232, ZN => n2967);
   U1036 : OAI22_X1 port map( A1 => n30117, A2 => n36662, B1 => n30329, B2 => 
                           n36708, ZN => n36233);
   U1037 : INV_X1 port map( A => n36233, ZN => n2968);
   U1038 : OAI22_X1 port map( A1 => n30085, A2 => n36730, B1 => n30563, B2 => 
                           n36710, ZN => n36234);
   U1039 : INV_X1 port map( A => n36234, ZN => n2805);
   U1040 : OAI22_X1 port map( A1 => n30116, A2 => n36662, B1 => n30330, B2 => 
                           n36717, ZN => n36235);
   U1041 : INV_X1 port map( A => n36235, ZN => n2969);
   U1042 : OAI22_X1 port map( A1 => n30085, A2 => n36472, B1 => n30569, B2 => 
                           n36710, ZN => n36236);
   U1043 : INV_X1 port map( A => n36236, ZN => n2897);
   U1044 : OAI22_X1 port map( A1 => n30086, A2 => n36472, B1 => n30570, B2 => 
                           n36736, ZN => n36237);
   U1045 : INV_X1 port map( A => n36237, ZN => n2898);
   U1046 : OAI22_X1 port map( A1 => n30123, A2 => n36715, B1 => n30319, B2 => 
                           n36703, ZN => n36238);
   U1047 : INV_X1 port map( A => n36238, ZN => n2870);
   U1048 : OAI22_X1 port map( A1 => n30120, A2 => n36715, B1 => n30320, B2 => 
                           n36705, ZN => n36239);
   U1049 : INV_X1 port map( A => n36239, ZN => n2871);
   U1050 : OAI22_X1 port map( A1 => n30124, A2 => n36469, B1 => n30363, B2 => 
                           n36714, ZN => n36240);
   U1051 : INV_X1 port map( A => n36240, ZN => n3381);
   U1052 : OAI22_X1 port map( A1 => n30109, A2 => n36701, B1 => n30336, B2 => 
                           n36726, ZN => n36241);
   U1053 : INV_X1 port map( A => n36241, ZN => n2918);
   U1054 : OAI22_X1 port map( A1 => n30120, A2 => n36449, B1 => n30362, B2 => 
                           n36705, ZN => n36242);
   U1055 : INV_X1 port map( A => n36242, ZN => n3066);
   U1056 : OAI22_X1 port map( A1 => n30116, A2 => n36677, B1 => n30361, B2 => 
                           n36717, ZN => n36243);
   U1057 : INV_X1 port map( A => n36243, ZN => n3046);
   U1058 : OAI22_X1 port map( A1 => n30117, A2 => n36715, B1 => n30322, B2 => 
                           n36708, ZN => n36244);
   U1059 : INV_X1 port map( A => n36244, ZN => n2872);
   U1060 : OAI22_X1 port map( A1 => n30116, A2 => n36454, B1 => n30350, B2 => 
                           n36717, ZN => n36245);
   U1061 : INV_X1 port map( A => n36245, ZN => n3344);
   U1062 : OAI22_X1 port map( A1 => n30117, A2 => n36454, B1 => n30349, B2 => 
                           n36708, ZN => n36246);
   U1063 : INV_X1 port map( A => n36246, ZN => n3343);
   U1064 : OAI22_X1 port map( A1 => n30120, A2 => n36280, B1 => n30359, B2 => 
                           n36705, ZN => n36247);
   U1065 : INV_X1 port map( A => n36247, ZN => n3348);
   U1066 : OAI22_X1 port map( A1 => n30116, A2 => n36715, B1 => n30323, B2 => 
                           n36717, ZN => n36248);
   U1067 : INV_X1 port map( A => n36248, ZN => n2873);
   U1068 : OAI22_X1 port map( A1 => n30109, A2 => n36303, B1 => n30355, B2 => 
                           n36726, ZN => n36249);
   U1069 : INV_X1 port map( A => n36249, ZN => n3379);
   U1070 : OAI22_X1 port map( A1 => n30120, A2 => n36303, B1 => n30358, B2 => 
                           n36705, ZN => n36250);
   U1071 : INV_X1 port map( A => n36250, ZN => n3380);
   U1072 : OAI22_X1 port map( A1 => n30086, A2 => n36751, B1 => n30551, B2 => 
                           n36736, ZN => n36251);
   U1073 : INV_X1 port map( A => n36251, ZN => n2803);
   U1074 : OAI22_X1 port map( A1 => n30123, A2 => n36662, B1 => n30327, B2 => 
                           n36703, ZN => n36252);
   U1075 : INV_X1 port map( A => n36252, ZN => n2966);
   U1076 : OAI22_X1 port map( A1 => n30109, A2 => n36662, B1 => n30333, B2 => 
                           n36726, ZN => n36253);
   U1077 : INV_X1 port map( A => n36253, ZN => n2971);
   U1078 : OAI22_X1 port map( A1 => n30085, A2 => n36487, B1 => n30559, B2 => 
                           n36710, ZN => n36254);
   U1079 : INV_X1 port map( A => n36254, ZN => n2838);
   U1080 : OAI22_X1 port map( A1 => n30116, A2 => n36469, B1 => n30346, B2 => 
                           n36717, ZN => n36255);
   U1081 : INV_X1 port map( A => n36255, ZN => n3376);
   U1082 : OAI22_X1 port map( A1 => n30109, A2 => n36280, B1 => n30354, B2 => 
                           n36726, ZN => n36256);
   U1083 : INV_X1 port map( A => n36256, ZN => n3347);
   U1084 : OAI22_X1 port map( A1 => n30117, A2 => n36751, B1 => n30977, B2 => 
                           n36708, ZN => n36257);
   U1085 : INV_X1 port map( A => n36257, ZN => n2797);
   U1086 : OAI22_X1 port map( A1 => n30117, A2 => n36449, B1 => n30351, B2 => 
                           n36708, ZN => n36258);
   U1087 : INV_X1 port map( A => n36258, ZN => n3062);
   U1088 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30104, ZN => n36811);
   U1089 : OAI22_X1 port map( A1 => n30104, A2 => n36431, B1 => n30725, B2 => 
                           n36811, ZN => n36259);
   U1090 : INV_X1 port map( A => n36259, ZN => n3114);
   U1091 : OAI22_X1 port map( A1 => n30104, A2 => n36433, B1 => n30724, B2 => 
                           n36811, ZN => n36260);
   U1092 : INV_X1 port map( A => n36260, ZN => n3081);
   U1093 : OAI22_X1 port map( A1 => n30104, A2 => n36449, B1 => n30721, B2 => 
                           n36811, ZN => n36261);
   U1094 : INV_X1 port map( A => n36261, ZN => n3076);
   U1095 : OAI22_X1 port map( A1 => n30104, A2 => n36692, B1 => n30720, B2 => 
                           n36811, ZN => n36262);
   U1096 : INV_X1 port map( A => n36262, ZN => n2953);
   U1097 : OAI22_X1 port map( A1 => n30104, A2 => n36701, B1 => n30718, B2 => 
                           n36811, ZN => n36263);
   U1098 : INV_X1 port map( A => n36263, ZN => n2921);
   U1099 : OAI22_X1 port map( A1 => n30104, A2 => n36472, B1 => n30717, B2 => 
                           n36811, ZN => n36264);
   U1100 : INV_X1 port map( A => n36264, ZN => n2908);
   U1101 : OAI22_X1 port map( A1 => n30104, A2 => n36487, B1 => n30716, B2 => 
                           n36811, ZN => n36265);
   U1102 : INV_X1 port map( A => n36265, ZN => n2848);
   U1103 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30095, ZN => n36807);
   U1104 : OAI22_X1 port map( A1 => n30095, A2 => n36296, B1 => n31153, B2 => 
                           n36807, ZN => n36266);
   U1105 : INV_X1 port map( A => n36266, ZN => n3308);
   U1106 : OAI22_X1 port map( A1 => n30104, A2 => n36296, B1 => n31151, B2 => 
                           n36811, ZN => n36267);
   U1107 : INV_X1 port map( A => n36267, ZN => n3306);
   U1108 : OAI22_X1 port map( A1 => n30098, A2 => n36454, B1 => n31150, B2 => 
                           n36833, ZN => n36268);
   U1109 : INV_X1 port map( A => n36268, ZN => n3342);
   U1110 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30091, ZN => n36803);
   U1111 : OAI22_X1 port map( A1 => n30091, A2 => n36296, B1 => n31149, B2 => 
                           n36803, ZN => n36269);
   U1112 : INV_X1 port map( A => n36269, ZN => n3305);
   U1113 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30092, ZN => n36801);
   U1114 : OAI22_X1 port map( A1 => n30092, A2 => n36296, B1 => n31148, B2 => 
                           n36801, ZN => n36270);
   U1115 : INV_X1 port map( A => n36270, ZN => n3304);
   U1116 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30100, ZN => n36805);
   U1117 : OAI22_X1 port map( A1 => n30100, A2 => n36441, B1 => n31147, B2 => 
                           n36805, ZN => n36271);
   U1118 : INV_X1 port map( A => n36271, ZN => n3406);
   U1119 : OAI22_X1 port map( A1 => n30100, A2 => n36327, B1 => n31145, B2 => 
                           n36805, ZN => n36272);
   U1120 : INV_X1 port map( A => n36272, ZN => n3438);
   U1121 : OAI22_X1 port map( A1 => n30091, A2 => n36280, B1 => n31143, B2 => 
                           n36803, ZN => n36273);
   U1122 : INV_X1 port map( A => n36273, ZN => n3340);
   U1123 : OAI22_X1 port map( A1 => n30092, A2 => n36403, B1 => n31142, B2 => 
                           n36801, ZN => n36274);
   U1124 : INV_X1 port map( A => n36274, ZN => n3470);
   U1125 : OAI22_X1 port map( A1 => n30094, A2 => n36282, B1 => n31138, B2 => 
                           n36813, ZN => n36275);
   U1126 : INV_X1 port map( A => n36275, ZN => n3468);
   U1127 : OAI22_X1 port map( A1 => n30094, A2 => n36515, B1 => n31137, B2 => 
                           n36813, ZN => n36276);
   U1128 : INV_X1 port map( A => n36276, ZN => n3333);
   U1129 : OAI22_X1 port map( A1 => n30095, A2 => n36282, B1 => n31136, B2 => 
                           n36807, ZN => n36277);
   U1130 : INV_X1 port map( A => n36277, ZN => n3467);
   U1131 : OAI22_X1 port map( A1 => n30091, A2 => n36282, B1 => n31135, B2 => 
                           n36803, ZN => n36278);
   U1132 : INV_X1 port map( A => n36278, ZN => n3466);
   U1133 : OAI22_X1 port map( A1 => n30104, A2 => n36280, B1 => n31133, B2 => 
                           n36811, ZN => n36279);
   U1134 : INV_X1 port map( A => n36279, ZN => n3339);
   U1135 : OAI22_X1 port map( A1 => n30100, A2 => n36280, B1 => n31131, B2 => 
                           n36805, ZN => n36281);
   U1136 : INV_X1 port map( A => n36281, ZN => n3337);
   U1137 : OAI22_X1 port map( A1 => n30098, A2 => n36282, B1 => n31127, B2 => 
                           n36833, ZN => n36283);
   U1138 : INV_X1 port map( A => n36283, ZN => n3463);
   U1139 : OAI22_X1 port map( A1 => n30100, A2 => n36469, B1 => n31126, B2 => 
                           n36805, ZN => n36284);
   U1140 : INV_X1 port map( A => n36284, ZN => n3374);
   U1141 : OAI22_X1 port map( A1 => n30100, A2 => n36515, B1 => n31125, B2 => 
                           n36805, ZN => n36285);
   U1142 : INV_X1 port map( A => n36285, ZN => n3331);
   U1143 : OAI22_X1 port map( A1 => n30092, A2 => n36454, B1 => n31122, B2 => 
                           n36801, ZN => n36286);
   U1144 : INV_X1 port map( A => n36286, ZN => n3364);
   U1145 : OAI22_X1 port map( A1 => n30095, A2 => n36454, B1 => n31121, B2 => 
                           n36807, ZN => n36287);
   U1146 : INV_X1 port map( A => n36287, ZN => n3363);
   U1147 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30102, ZN => n36835);
   U1148 : OAI22_X1 port map( A1 => n30102, A2 => n36788, B1 => n30956, B2 => 
                           n36835, ZN => n36288);
   U1149 : INV_X1 port map( A => n36288, ZN => n2828);
   U1150 : OAI22_X1 port map( A1 => n30095, A2 => n36303, B1 => n31120, B2 => 
                           n36807, ZN => n36289);
   U1151 : INV_X1 port map( A => n36289, ZN => n3373);
   U1152 : OAI22_X1 port map( A1 => n30095, A2 => n36315, B1 => n31119, B2 => 
                           n36807, ZN => n36290);
   U1153 : INV_X1 port map( A => n36290, ZN => n3405);
   U1154 : OAI22_X1 port map( A1 => n30094, A2 => n36454, B1 => n31118, B2 => 
                           n36813, ZN => n36291);
   U1155 : INV_X1 port map( A => n36291, ZN => n3362);
   U1156 : OAI22_X1 port map( A1 => n30102, A2 => n36751, B1 => n30951, B2 => 
                           n36835, ZN => n36292);
   U1157 : INV_X1 port map( A => n36292, ZN => n2793);
   U1158 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n30115, ZN => n36799);
   U1159 : OAI22_X1 port map( A1 => n30115, A2 => n36788, B1 => n30948, B2 => 
                           n36799, ZN => n36293);
   U1160 : INV_X1 port map( A => n36293, ZN => n2822);
   U1161 : OAI22_X1 port map( A1 => n30092, A2 => n36303, B1 => n31114, B2 => 
                           n36801, ZN => n36294);
   U1162 : INV_X1 port map( A => n36294, ZN => n3371);
   U1163 : OAI22_X1 port map( A1 => n30115, A2 => n36751, B1 => n30946, B2 => 
                           n36799, ZN => n36295);
   U1164 : INV_X1 port map( A => n36295, ZN => n2791);
   U1165 : OAI22_X1 port map( A1 => n30098, A2 => n36296, B1 => n31152, B2 => 
                           n36833, ZN => n36297);
   U1166 : INV_X1 port map( A => n36297, ZN => n3307);
   U1167 : OAI22_X1 port map( A1 => n30095, A2 => n36489, B1 => n31113, B2 => 
                           n36807, ZN => n36298);
   U1168 : INV_X1 port map( A => n36298, ZN => n3436);
   U1169 : OAI22_X1 port map( A1 => n30091, A2 => n36303, B1 => n31112, B2 => 
                           n36803, ZN => n36299);
   U1170 : INV_X1 port map( A => n36299, ZN => n3370);
   U1171 : OAI22_X1 port map( A1 => n30098, A2 => n36303, B1 => n31111, B2 => 
                           n36833, ZN => n36300);
   U1172 : INV_X1 port map( A => n36300, ZN => n3369);
   U1173 : OAI22_X1 port map( A1 => n30098, A2 => n36321, B1 => n31110, B2 => 
                           n36833, ZN => n36301);
   U1174 : INV_X1 port map( A => n36301, ZN => n3501);
   U1175 : OAI22_X1 port map( A1 => n30095, A2 => n36321, B1 => n31108, B2 => 
                           n36807, ZN => n36302);
   U1176 : INV_X1 port map( A => n36302, ZN => n3500);
   U1177 : OAI22_X1 port map( A1 => n30104, A2 => n36303, B1 => n31107, B2 => 
                           n36811, ZN => n36304);
   U1178 : INV_X1 port map( A => n36304, ZN => n3367);
   U1179 : OAI22_X1 port map( A1 => n30104, A2 => n36315, B1 => n31106, B2 => 
                           n36811, ZN => n36305);
   U1180 : INV_X1 port map( A => n36305, ZN => n3403);
   U1181 : OAI22_X1 port map( A1 => n30104, A2 => n36489, B1 => n31105, B2 => 
                           n36811, ZN => n36306);
   U1182 : INV_X1 port map( A => n36306, ZN => n3435);
   U1183 : OAI22_X1 port map( A1 => n30104, A2 => n36403, B1 => n31102, B2 => 
                           n36811, ZN => n36307);
   U1184 : INV_X1 port map( A => n36307, ZN => n3493);
   U1185 : OAI22_X1 port map( A1 => n30104, A2 => n36321, B1 => n31100, B2 => 
                           n36811, ZN => n36308);
   U1186 : INV_X1 port map( A => n36308, ZN => n3499);
   U1187 : OAI22_X1 port map( A1 => n30115, A2 => n36472, B1 => n30934, B2 => 
                           n36799, ZN => n36309);
   U1188 : INV_X1 port map( A => n36309, ZN => n2916);
   U1189 : OAI22_X1 port map( A1 => n30115, A2 => n36515, B1 => n30933, B2 => 
                           n36799, ZN => n36310);
   U1190 : INV_X1 port map( A => n36310, ZN => n3320);
   U1191 : OAI22_X1 port map( A1 => n30094, A2 => n36469, B1 => n31099, B2 => 
                           n36813, ZN => n36311);
   U1192 : INV_X1 port map( A => n36311, ZN => n3394);
   U1193 : OAI22_X1 port map( A1 => n30091, A2 => n36315, B1 => n31095, B2 => 
                           n36803, ZN => n36312);
   U1194 : INV_X1 port map( A => n36312, ZN => n3402);
   U1195 : OAI22_X1 port map( A1 => n30098, A2 => n36315, B1 => n31094, B2 => 
                           n36833, ZN => n36313);
   U1196 : INV_X1 port map( A => n36313, ZN => n3401);
   U1197 : OAI22_X1 port map( A1 => n30094, A2 => n36315, B1 => n31093, B2 => 
                           n36813, ZN => n36314);
   U1198 : INV_X1 port map( A => n36314, ZN => n3400);
   U1199 : OAI22_X1 port map( A1 => n30092, A2 => n36315, B1 => n31092, B2 => 
                           n36801, ZN => n36316);
   U1200 : INV_X1 port map( A => n36316, ZN => n3399);
   U1201 : OAI22_X1 port map( A1 => n30094, A2 => n36489, B1 => n31091, B2 => 
                           n36813, ZN => n36317);
   U1202 : INV_X1 port map( A => n36317, ZN => n3433);
   U1203 : OAI22_X1 port map( A1 => n30092, A2 => n36489, B1 => n31090, B2 => 
                           n36801, ZN => n36318);
   U1204 : INV_X1 port map( A => n36318, ZN => n3432);
   U1205 : OAI22_X1 port map( A1 => n30094, A2 => n36321, B1 => n31089, B2 => 
                           n36813, ZN => n36319);
   U1206 : INV_X1 port map( A => n36319, ZN => n3497);
   U1207 : OAI22_X1 port map( A1 => n30092, A2 => n36321, B1 => n31088, B2 => 
                           n36801, ZN => n36320);
   U1208 : INV_X1 port map( A => n36320, ZN => n3496);
   U1209 : OAI22_X1 port map( A1 => n30091, A2 => n36321, B1 => n31085, B2 => 
                           n36803, ZN => n36322);
   U1210 : INV_X1 port map( A => n36322, ZN => n3495);
   U1211 : OAI22_X1 port map( A1 => n30091, A2 => n36489, B1 => n31084, B2 => 
                           n36803, ZN => n36323);
   U1212 : INV_X1 port map( A => n36323, ZN => n3431);
   U1213 : OAI22_X1 port map( A1 => n30098, A2 => n36327, B1 => n31083, B2 => 
                           n36833, ZN => n36324);
   U1214 : INV_X1 port map( A => n36324, ZN => n3461);
   U1215 : OAI22_X1 port map( A1 => n30100, A2 => n36403, B1 => n31079, B2 => 
                           n36805, ZN => n36325);
   U1216 : INV_X1 port map( A => n36325, ZN => n3490);
   U1217 : OAI22_X1 port map( A1 => n30100, A2 => n36425, B1 => n31073, B2 => 
                           n36805, ZN => n36326);
   U1218 : INV_X1 port map( A => n36326, ZN => n3522);
   U1219 : OAI22_X1 port map( A1 => n30102, A2 => n36327, B1 => n31068, B2 => 
                           n36835, ZN => n36328);
   U1220 : INV_X1 port map( A => n36328, ZN => n3457);
   U1221 : OAI22_X1 port map( A1 => n30102, A2 => n36403, B1 => n31065, B2 => 
                           n36835, ZN => n36329);
   U1222 : INV_X1 port map( A => n36329, ZN => n3489);
   U1223 : OAI22_X1 port map( A1 => n30102, A2 => n36425, B1 => n31064, B2 => 
                           n36835, ZN => n36330);
   U1224 : INV_X1 port map( A => n36330, ZN => n3520);
   U1225 : OAI22_X1 port map( A1 => n30115, A2 => n36643, B1 => n30913, B2 => 
                           n36799, ZN => n36331);
   U1226 : INV_X1 port map( A => n36331, ZN => n3235);
   U1227 : OAI22_X1 port map( A1 => n30102, A2 => n36469, B1 => n31062, B2 => 
                           n36835, ZN => n36332);
   U1228 : INV_X1 port map( A => n36332, ZN => n3392);
   U1229 : OAI22_X1 port map( A1 => n30102, A2 => n36441, B1 => n31060, B2 => 
                           n36835, ZN => n36333);
   U1230 : INV_X1 port map( A => n36333, ZN => n3424);
   U1231 : OAI22_X1 port map( A1 => n30102, A2 => n36515, B1 => n31058, B2 => 
                           n36835, ZN => n36334);
   U1232 : INV_X1 port map( A => n36334, ZN => n3328);
   U1233 : OAI22_X1 port map( A1 => n30098, A2 => n36429, B1 => n30909, B2 => 
                           n36833, ZN => n36335);
   U1234 : INV_X1 port map( A => n36335, ZN => n3149);
   U1235 : OAI22_X1 port map( A1 => n30102, A2 => n36454, B1 => n31057, B2 => 
                           n36835, ZN => n36336);
   U1236 : INV_X1 port map( A => n36336, ZN => n3360);
   U1237 : OAI22_X1 port map( A1 => n30094, A2 => n36493, B1 => n31046, B2 => 
                           n36813, ZN => n36337);
   U1238 : INV_X1 port map( A => n36337, ZN => n3534);
   U1239 : OAI22_X1 port map( A1 => n30098, A2 => n36748, B1 => n30906, B2 => 
                           n36833, ZN => n36338);
   U1240 : INV_X1 port map( A => n36338, ZN => n3086);
   U1241 : OAI22_X1 port map( A1 => n30098, A2 => n36712, B1 => n30905, B2 => 
                           n36833, ZN => n36339);
   U1242 : INV_X1 port map( A => n36339, ZN => n3119);
   U1243 : OAI22_X1 port map( A1 => n30098, A2 => n36579, B1 => n30904, B2 => 
                           n36833, ZN => n36340);
   U1244 : INV_X1 port map( A => n36340, ZN => n3021);
   U1245 : OAI22_X1 port map( A1 => n30098, A2 => n36677, B1 => n30903, B2 => 
                           n36833, ZN => n36341);
   U1246 : INV_X1 port map( A => n36341, ZN => n3050);
   U1247 : OAI22_X1 port map( A1 => n30098, A2 => n36662, B1 => n30902, B2 => 
                           n36833, ZN => n36342);
   U1248 : INV_X1 port map( A => n36342, ZN => n2958);
   U1249 : OAI22_X1 port map( A1 => n30098, A2 => n36718, B1 => n30901, B2 => 
                           n36833, ZN => n36343);
   U1250 : INV_X1 port map( A => n36343, ZN => n2926);
   U1251 : OAI22_X1 port map( A1 => n30098, A2 => n36472, B1 => n30900, B2 => 
                           n36833, ZN => n36344);
   U1252 : INV_X1 port map( A => n36344, ZN => n2911);
   U1253 : OAI22_X1 port map( A1 => n30098, A2 => n36715, B1 => n30899, B2 => 
                           n36833, ZN => n36345);
   U1254 : INV_X1 port map( A => n36345, ZN => n2862);
   U1255 : OAI22_X1 port map( A1 => n30098, A2 => n36487, B1 => n30898, B2 => 
                           n36833, ZN => n36346);
   U1256 : INV_X1 port map( A => n36346, ZN => n2851);
   U1257 : OAI22_X1 port map( A1 => n30098, A2 => n36730, B1 => n30897, B2 => 
                           n36833, ZN => n36347);
   U1258 : INV_X1 port map( A => n36347, ZN => n2819);
   U1259 : OAI22_X1 port map( A1 => n30091, A2 => n36579, B1 => n30895, B2 => 
                           n36803, ZN => n36348);
   U1260 : INV_X1 port map( A => n36348, ZN => n3020);
   U1261 : OAI22_X1 port map( A1 => n30092, A2 => n36579, B1 => n30893, B2 => 
                           n36801, ZN => n36349);
   U1262 : INV_X1 port map( A => n36349, ZN => n3019);
   U1263 : OAI22_X1 port map( A1 => n30098, A2 => n36618, B1 => n30890, B2 => 
                           n36833, ZN => n36350);
   U1264 : INV_X1 port map( A => n36350, ZN => n2986);
   U1265 : OAI22_X1 port map( A1 => n30095, A2 => n36579, B1 => n30887, B2 => 
                           n36807, ZN => n36351);
   U1266 : INV_X1 port map( A => n36351, ZN => n3017);
   U1267 : OAI22_X1 port map( A1 => n30100, A2 => n36683, B1 => n30882, B2 => 
                           n36805, ZN => n36352);
   U1268 : INV_X1 port map( A => n36352, ZN => n3045);
   U1269 : OAI22_X1 port map( A1 => n30094, A2 => n36683, B1 => n30881, B2 => 
                           n36813, ZN => n36353);
   U1270 : INV_X1 port map( A => n36353, ZN => n3044);
   U1271 : OAI22_X1 port map( A1 => n30102, A2 => n36683, B1 => n30879, B2 => 
                           n36835, ZN => n36354);
   U1272 : INV_X1 port map( A => n36354, ZN => n3042);
   U1273 : OAI22_X1 port map( A1 => n30104, A2 => n36579, B1 => n30877, B2 => 
                           n36811, ZN => n36355);
   U1274 : INV_X1 port map( A => n36355, ZN => n3015);
   U1275 : OAI22_X1 port map( A1 => n30100, A2 => n36618, B1 => n30861, B2 => 
                           n36805, ZN => n36356);
   U1276 : INV_X1 port map( A => n36356, ZN => n2984);
   U1277 : OAI22_X1 port map( A1 => n30102, A2 => n36398, B1 => n30859, B2 => 
                           n36835, ZN => n36357);
   U1278 : INV_X1 port map( A => n36357, ZN => n3013);
   U1279 : OAI22_X1 port map( A1 => n30104, A2 => n36398, B1 => n30857, B2 => 
                           n36811, ZN => n36358);
   U1280 : INV_X1 port map( A => n36358, ZN => n3011);
   U1281 : OAI22_X1 port map( A1 => n30091, A2 => n36398, B1 => n30854, B2 => 
                           n36803, ZN => n36359);
   U1282 : INV_X1 port map( A => n36359, ZN => n3010);
   U1283 : OAI22_X1 port map( A1 => n30092, A2 => n36398, B1 => n30853, B2 => 
                           n36801, ZN => n36360);
   U1284 : INV_X1 port map( A => n36360, ZN => n3009);
   U1285 : OAI22_X1 port map( A1 => n30094, A2 => n36398, B1 => n30851, B2 => 
                           n36813, ZN => n36361);
   U1286 : INV_X1 port map( A => n36361, ZN => n3007);
   U1287 : OAI22_X1 port map( A1 => n30095, A2 => n36398, B1 => n30850, B2 => 
                           n36807, ZN => n36362);
   U1288 : INV_X1 port map( A => n36362, ZN => n3006);
   U1289 : OAI22_X1 port map( A1 => n30098, A2 => n36427, B1 => n30848, B2 => 
                           n36833, ZN => n36363);
   U1290 : INV_X1 port map( A => n36363, ZN => n3174);
   U1291 : OAI22_X1 port map( A1 => n30102, A2 => n36584, B1 => n31000, B2 => 
                           n36835, ZN => n36364);
   U1292 : INV_X1 port map( A => n36364, ZN => n2889);
   U1293 : OAI22_X1 port map( A1 => n30100, A2 => n36477, B1 => n30836, B2 => 
                           n36805, ZN => n36365);
   U1294 : INV_X1 port map( A => n36365, ZN => n2859);
   U1295 : OAI22_X1 port map( A1 => n30102, A2 => n36477, B1 => n30834, B2 => 
                           n36835, ZN => n36366);
   U1296 : INV_X1 port map( A => n36366, ZN => n2857);
   U1297 : OAI22_X1 port map( A1 => n30104, A2 => n36477, B1 => n30832, B2 => 
                           n36811, ZN => n36367);
   U1298 : INV_X1 port map( A => n36367, ZN => n2855);
   U1299 : OAI22_X1 port map( A1 => n30091, A2 => n36715, B1 => n30827, B2 => 
                           n36803, ZN => n36368);
   U1300 : INV_X1 port map( A => n36368, ZN => n2885);
   U1301 : OAI22_X1 port map( A1 => n30092, A2 => n36715, B1 => n30826, B2 => 
                           n36801, ZN => n36369);
   U1302 : INV_X1 port map( A => n36369, ZN => n2884);
   U1303 : OAI22_X1 port map( A1 => n30094, A2 => n36715, B1 => n30824, B2 => 
                           n36813, ZN => n36370);
   U1304 : INV_X1 port map( A => n36370, ZN => n2882);
   U1305 : OAI22_X1 port map( A1 => n30095, A2 => n36715, B1 => n30823, B2 => 
                           n36807, ZN => n36371);
   U1306 : INV_X1 port map( A => n36371, ZN => n2881);
   U1307 : OAI22_X1 port map( A1 => n30102, A2 => n36643, B1 => n30818, B2 => 
                           n36835, ZN => n36372);
   U1308 : INV_X1 port map( A => n36372, ZN => n3233);
   U1309 : OAI22_X1 port map( A1 => n30102, A2 => n36422, B1 => n30817, B2 => 
                           n36835, ZN => n36373);
   U1310 : INV_X1 port map( A => n36373, ZN => n3244);
   U1311 : OAI22_X1 port map( A1 => n30102, A2 => n36420, B1 => n30816, B2 => 
                           n36835, ZN => n36374);
   U1312 : INV_X1 port map( A => n36374, ZN => n3277);
   U1313 : OAI22_X1 port map( A1 => n30102, A2 => n36427, B1 => n30815, B2 => 
                           n36835, ZN => n36375);
   U1314 : INV_X1 port map( A => n36375, ZN => n3176);
   U1315 : OAI22_X1 port map( A1 => n30102, A2 => n36429, B1 => n30814, B2 => 
                           n36835, ZN => n36376);
   U1316 : INV_X1 port map( A => n36376, ZN => n3147);
   U1317 : OAI22_X1 port map( A1 => n30102, A2 => n36431, B1 => n30813, B2 => 
                           n36835, ZN => n36377);
   U1318 : INV_X1 port map( A => n36377, ZN => n3117);
   U1319 : OAI22_X1 port map( A1 => n30102, A2 => n36433, B1 => n30812, B2 => 
                           n36835, ZN => n36378);
   U1320 : INV_X1 port map( A => n36378, ZN => n3084);
   U1321 : OAI22_X1 port map( A1 => n30102, A2 => n36677, B1 => n30811, B2 => 
                           n36835, ZN => n36379);
   U1322 : INV_X1 port map( A => n36379, ZN => n3048);
   U1323 : OAI22_X1 port map( A1 => n30102, A2 => n36692, B1 => n30810, B2 => 
                           n36835, ZN => n36380);
   U1324 : INV_X1 port map( A => n36380, ZN => n2956);
   U1325 : OAI22_X1 port map( A1 => n30102, A2 => n36701, B1 => n30809, B2 => 
                           n36835, ZN => n36381);
   U1326 : INV_X1 port map( A => n36381, ZN => n2924);
   U1327 : OAI22_X1 port map( A1 => n30104, A2 => n36420, B1 => n30734, B2 => 
                           n36811, ZN => n36382);
   U1328 : INV_X1 port map( A => n36382, ZN => n3274);
   U1329 : OAI22_X1 port map( A1 => n30104, A2 => n36422, B1 => n30732, B2 => 
                           n36811, ZN => n36383);
   U1330 : INV_X1 port map( A => n36383, ZN => n3241);
   U1331 : OAI22_X1 port map( A1 => n30104, A2 => n36643, B1 => n30730, B2 => 
                           n36811, ZN => n36384);
   U1332 : INV_X1 port map( A => n36384, ZN => n3232);
   U1333 : OAI22_X1 port map( A1 => n30104, A2 => n36427, B1 => n30727, B2 => 
                           n36811, ZN => n36385);
   U1334 : INV_X1 port map( A => n36385, ZN => n3179);
   U1335 : OAI22_X1 port map( A1 => n30104, A2 => n36429, B1 => n30726, B2 => 
                           n36811, ZN => n36386);
   U1336 : INV_X1 port map( A => n36386, ZN => n3144);
   U1337 : OAI22_X1 port map( A1 => n30100, A2 => n36730, B1 => n30715, B2 => 
                           n36805, ZN => n36387);
   U1338 : INV_X1 port map( A => n36387, ZN => n2816);
   U1339 : OAI22_X1 port map( A1 => n30094, A2 => n36420, B1 => n30681, B2 => 
                           n36813, ZN => n36388);
   U1340 : INV_X1 port map( A => n36388, ZN => n3272);
   U1341 : OAI22_X1 port map( A1 => n30094, A2 => n36422, B1 => n30680, B2 => 
                           n36813, ZN => n36389);
   U1342 : INV_X1 port map( A => n36389, ZN => n3238);
   U1343 : OAI22_X1 port map( A1 => n30091, A2 => n36427, B1 => n30679, B2 => 
                           n36803, ZN => n36390);
   U1344 : INV_X1 port map( A => n36390, ZN => n3181);
   U1345 : OAI22_X1 port map( A1 => n30092, A2 => n36485, B1 => n30678, B2 => 
                           n36801, ZN => n36391);
   U1346 : INV_X1 port map( A => n36391, ZN => n3205);
   U1347 : OAI22_X1 port map( A1 => n30094, A2 => n36485, B1 => n30676, B2 => 
                           n36813, ZN => n36392);
   U1348 : INV_X1 port map( A => n36392, ZN => n3203);
   U1349 : OAI22_X1 port map( A1 => n30095, A2 => n36485, B1 => n30675, B2 => 
                           n36807, ZN => n36393);
   U1350 : INV_X1 port map( A => n36393, ZN => n3202);
   U1351 : OAI22_X1 port map( A1 => n30094, A2 => n36429, B1 => n30672, B2 => 
                           n36813, ZN => n36394);
   U1352 : INV_X1 port map( A => n36394, ZN => n3142);
   U1353 : OAI22_X1 port map( A1 => n30094, A2 => n36431, B1 => n30671, B2 => 
                           n36813, ZN => n36395);
   U1354 : INV_X1 port map( A => n36395, ZN => n3112);
   U1355 : OAI22_X1 port map( A1 => n30094, A2 => n36433, B1 => n30670, B2 => 
                           n36813, ZN => n36396);
   U1356 : INV_X1 port map( A => n36396, ZN => n3079);
   U1357 : OAI22_X1 port map( A1 => n30094, A2 => n36449, B1 => n30669, B2 => 
                           n36813, ZN => n36397);
   U1358 : INV_X1 port map( A => n36397, ZN => n3074);
   U1359 : OAI22_X1 port map( A1 => n30115, A2 => n36398, B1 => n30408, B2 => 
                           n36799, ZN => n36399);
   U1360 : INV_X1 port map( A => n36399, ZN => n3003);
   U1361 : OAI22_X1 port map( A1 => n30094, A2 => n36692, B1 => n30668, B2 => 
                           n36813, ZN => n36400);
   U1362 : INV_X1 port map( A => n36400, ZN => n2951);
   U1363 : OAI22_X1 port map( A1 => n30094, A2 => n36701, B1 => n30667, B2 => 
                           n36813, ZN => n36401);
   U1364 : INV_X1 port map( A => n36401, ZN => n2919);
   U1365 : OAI22_X1 port map( A1 => n30094, A2 => n36472, B1 => n30666, B2 => 
                           n36813, ZN => n36402);
   U1366 : INV_X1 port map( A => n36402, ZN => n2906);
   U1367 : OAI22_X1 port map( A1 => n30115, A2 => n36403, B1 => n30396, B2 => 
                           n36799, ZN => n36404);
   U1368 : INV_X1 port map( A => n36404, ZN => n3478);
   U1369 : OAI22_X1 port map( A1 => n30094, A2 => n36643, B1 => n30684, B2 => 
                           n36813, ZN => n36405);
   U1370 : INV_X1 port map( A => n36405, ZN => n3227);
   U1371 : OAI22_X1 port map( A1 => n30094, A2 => n36487, B1 => n30665, B2 => 
                           n36813, ZN => n36406);
   U1372 : INV_X1 port map( A => n36406, ZN => n2846);
   U1373 : OAI22_X1 port map( A1 => n30091, A2 => n36783, B1 => n30664, B2 => 
                           n36803, ZN => n36407);
   U1374 : INV_X1 port map( A => n36407, ZN => n3173);
   U1375 : OAI22_X1 port map( A1 => n30092, A2 => n36783, B1 => n30663, B2 => 
                           n36801, ZN => n36408);
   U1376 : INV_X1 port map( A => n36408, ZN => n3172);
   U1377 : OAI22_X1 port map( A1 => n30095, A2 => n36783, B1 => n30661, B2 => 
                           n36807, ZN => n36409);
   U1378 : INV_X1 port map( A => n36409, ZN => n3170);
   U1379 : OAI22_X1 port map( A1 => n30094, A2 => n36730, B1 => n30658, B2 => 
                           n36813, ZN => n36410);
   U1380 : INV_X1 port map( A => n36410, ZN => n2814);
   U1381 : OAI22_X1 port map( A1 => n30091, A2 => n36712, B1 => n30657, B2 => 
                           n36803, ZN => n36411);
   U1382 : INV_X1 port map( A => n36411, ZN => n3141);
   U1383 : OAI22_X1 port map( A1 => n30092, A2 => n36643, B1 => n30686, B2 => 
                           n36801, ZN => n36412);
   U1384 : INV_X1 port map( A => n36412, ZN => n3229);
   U1385 : OAI22_X1 port map( A1 => n30092, A2 => n36712, B1 => n30656, B2 => 
                           n36801, ZN => n36413);
   U1386 : INV_X1 port map( A => n36413, ZN => n3140);
   U1387 : OAI22_X1 port map( A1 => n30091, A2 => n36643, B1 => n30687, B2 => 
                           n36803, ZN => n36414);
   U1388 : INV_X1 port map( A => n36414, ZN => n3230);
   U1389 : OAI22_X1 port map( A1 => n30091, A2 => n36422, B1 => n30688, B2 => 
                           n36803, ZN => n36415);
   U1390 : INV_X1 port map( A => n36415, ZN => n3239);
   U1391 : OAI22_X1 port map( A1 => n30095, A2 => n36712, B1 => n30654, B2 => 
                           n36807, ZN => n36416);
   U1392 : INV_X1 port map( A => n36416, ZN => n3138);
   U1393 : OAI22_X1 port map( A1 => n30095, A2 => n36420, B1 => n30651, B2 => 
                           n36807, ZN => n36417);
   U1394 : INV_X1 port map( A => n36417, ZN => n3271);
   U1395 : OAI22_X1 port map( A1 => n30095, A2 => n36674, B1 => n30650, B2 => 
                           n36807, ZN => n36418);
   U1396 : INV_X1 port map( A => n36418, ZN => n3269);
   U1397 : OAI22_X1 port map( A1 => n30095, A2 => n36748, B1 => n30649, B2 => 
                           n36807, ZN => n36419);
   U1398 : INV_X1 port map( A => n36419, ZN => n3109);
   U1399 : OAI22_X1 port map( A1 => n30100, A2 => n36420, B1 => n30693, B2 => 
                           n36805, ZN => n36421);
   U1400 : INV_X1 port map( A => n36421, ZN => n3273);
   U1401 : OAI22_X1 port map( A1 => n30100, A2 => n36422, B1 => n30694, B2 => 
                           n36805, ZN => n36423);
   U1402 : INV_X1 port map( A => n36423, ZN => n3240);
   U1403 : OAI22_X1 port map( A1 => n30100, A2 => n36643, B1 => n30695, B2 => 
                           n36805, ZN => n36424);
   U1404 : INV_X1 port map( A => n36424, ZN => n3231);
   U1405 : OAI22_X1 port map( A1 => n30115, A2 => n36425, B1 => n30386, B2 => 
                           n36799, ZN => n36426);
   U1406 : INV_X1 port map( A => n36426, ZN => n3504);
   U1407 : OAI22_X1 port map( A1 => n30100, A2 => n36427, B1 => n30696, B2 => 
                           n36805, ZN => n36428);
   U1408 : INV_X1 port map( A => n36428, ZN => n3180);
   U1409 : OAI22_X1 port map( A1 => n30100, A2 => n36429, B1 => n30697, B2 => 
                           n36805, ZN => n36430);
   U1410 : INV_X1 port map( A => n36430, ZN => n3143);
   U1411 : OAI22_X1 port map( A1 => n30100, A2 => n36431, B1 => n30698, B2 => 
                           n36805, ZN => n36432);
   U1412 : INV_X1 port map( A => n36432, ZN => n3113);
   U1413 : OAI22_X1 port map( A1 => n30100, A2 => n36433, B1 => n30699, B2 => 
                           n36805, ZN => n36434);
   U1414 : INV_X1 port map( A => n36434, ZN => n3080);
   U1415 : OAI22_X1 port map( A1 => n30095, A2 => n36449, B1 => n30648, B2 => 
                           n36807, ZN => n36435);
   U1416 : INV_X1 port map( A => n36435, ZN => n3073);
   U1417 : OAI22_X1 port map( A1 => n30091, A2 => n36449, B1 => n30647, B2 => 
                           n36803, ZN => n36436);
   U1418 : INV_X1 port map( A => n36436, ZN => n3072);
   U1419 : OAI22_X1 port map( A1 => n30100, A2 => n36449, B1 => n30701, B2 => 
                           n36805, ZN => n36437);
   U1420 : INV_X1 port map( A => n36437, ZN => n3075);
   U1421 : OAI22_X1 port map( A1 => n30100, A2 => n36692, B1 => n30702, B2 => 
                           n36805, ZN => n36438);
   U1422 : INV_X1 port map( A => n36438, ZN => n2952);
   U1423 : OAI22_X1 port map( A1 => n30092, A2 => n36449, B1 => n30646, B2 => 
                           n36801, ZN => n36439);
   U1424 : INV_X1 port map( A => n36439, ZN => n3071);
   U1425 : OAI22_X1 port map( A1 => n30098, A2 => n36643, B1 => n30642, B2 => 
                           n36833, ZN => n36440);
   U1426 : INV_X1 port map( A => n36440, ZN => n3225);
   U1427 : OAI22_X1 port map( A1 => n30115, A2 => n36441, B1 => n30370, B2 => 
                           n36799, ZN => n36442);
   U1428 : INV_X1 port map( A => n36442, ZN => n3408);
   U1429 : OAI22_X1 port map( A1 => n30115, A2 => n36674, B1 => n30237, B2 => 
                           n36799, ZN => n36443);
   U1430 : INV_X1 port map( A => n36443, ZN => n3257);
   U1431 : OAI22_X1 port map( A1 => n30092, A2 => n36674, B1 => n30639, B2 => 
                           n36801, ZN => n36444);
   U1432 : INV_X1 port map( A => n36444, ZN => n3266);
   U1433 : OAI22_X1 port map( A1 => n30098, A2 => n36674, B1 => n30638, B2 => 
                           n36833, ZN => n36445);
   U1434 : INV_X1 port map( A => n36445, ZN => n3265);
   U1435 : OAI22_X1 port map( A1 => n30092, A2 => n36457, B1 => n30630, B2 => 
                           n36801, ZN => n36446);
   U1436 : INV_X1 port map( A => n36446, ZN => n3300);
   U1437 : OAI22_X1 port map( A1 => n30091, A2 => n36457, B1 => n30629, B2 => 
                           n36803, ZN => n36447);
   U1438 : INV_X1 port map( A => n36447, ZN => n3299);
   U1439 : OAI22_X1 port map( A1 => n30095, A2 => n36643, B1 => n30683, B2 => 
                           n36807, ZN => n36448);
   U1440 : INV_X1 port map( A => n36448, ZN => n3226);
   U1441 : OAI22_X1 port map( A1 => n30115, A2 => n36449, B1 => n30360, B2 => 
                           n36799, ZN => n36450);
   U1442 : INV_X1 port map( A => n36450, ZN => n3065);
   U1443 : OAI22_X1 port map( A1 => n30115, A2 => n36457, B1 => n30253, B2 => 
                           n36799, ZN => n36451);
   U1444 : INV_X1 port map( A => n36451, ZN => n3290);
   U1445 : OAI22_X1 port map( A1 => n30092, A2 => n36730, B1 => n30624, B2 => 
                           n36801, ZN => n36452);
   U1446 : INV_X1 port map( A => n36452, ZN => n2812);
   U1447 : OAI22_X1 port map( A1 => n30092, A2 => n36487, B1 => n30623, B2 => 
                           n36801, ZN => n36453);
   U1448 : INV_X1 port map( A => n36453, ZN => n2844);
   U1449 : OAI22_X1 port map( A1 => n30115, A2 => n36454, B1 => n30352, B2 => 
                           n36799, ZN => n36455);
   U1450 : INV_X1 port map( A => n36455, ZN => n3345);
   U1451 : OAI22_X1 port map( A1 => n30115, A2 => n36748, B1 => n30269, B2 => 
                           n36799, ZN => n36456);
   U1452 : INV_X1 port map( A => n36456, ZN => n3097);
   U1453 : OAI22_X1 port map( A1 => n30098, A2 => n36457, B1 => n30627, B2 => 
                           n36833, ZN => n36458);
   U1454 : INV_X1 port map( A => n36458, ZN => n3298);
   U1455 : OAI22_X1 port map( A1 => n30100, A2 => n36701, B1 => n30712, B2 => 
                           n36805, ZN => n36459);
   U1456 : INV_X1 port map( A => n36459, ZN => n2920);
   U1457 : OAI22_X1 port map( A1 => n30092, A2 => n36662, B1 => n30620, B2 => 
                           n36801, ZN => n36460);
   U1458 : INV_X1 port map( A => n36460, ZN => n2980);
   U1459 : OAI22_X1 port map( A1 => n30100, A2 => n36472, B1 => n30713, B2 => 
                           n36805, ZN => n36461);
   U1460 : INV_X1 port map( A => n36461, ZN => n2907);
   U1461 : OAI22_X1 port map( A1 => n30095, A2 => n36472, B1 => n30596, B2 => 
                           n36807, ZN => n36462);
   U1462 : INV_X1 port map( A => n36462, ZN => n2900);
   U1463 : OAI22_X1 port map( A1 => n30092, A2 => n36472, B1 => n30622, B2 => 
                           n36801, ZN => n36463);
   U1464 : INV_X1 port map( A => n36463, ZN => n2904);
   U1465 : OAI22_X1 port map( A1 => n30092, A2 => n36718, B1 => n30621, B2 => 
                           n36801, ZN => n36464);
   U1466 : INV_X1 port map( A => n36464, ZN => n2948);
   U1467 : OAI22_X1 port map( A1 => n30115, A2 => n36712, B1 => n30278, B2 => 
                           n36799, ZN => n36465);
   U1468 : INV_X1 port map( A => n36465, ZN => n3126);
   U1469 : OAI22_X1 port map( A1 => n30091, A2 => n36718, B1 => n30614, B2 => 
                           n36803, ZN => n36466);
   U1470 : INV_X1 port map( A => n36466, ZN => n2947);
   U1471 : OAI22_X1 port map( A1 => n30092, A2 => n36748, B1 => n30619, B2 => 
                           n36801, ZN => n36467);
   U1472 : INV_X1 port map( A => n36467, ZN => n3107);
   U1473 : OAI22_X1 port map( A1 => n30091, A2 => n36730, B1 => n30617, B2 => 
                           n36803, ZN => n36468);
   U1474 : INV_X1 port map( A => n36468, ZN => n2811);
   U1475 : OAI22_X1 port map( A1 => n30115, A2 => n36469, B1 => n30345, B2 => 
                           n36799, ZN => n36470);
   U1476 : INV_X1 port map( A => n36470, ZN => n3375);
   U1477 : OAI22_X1 port map( A1 => n30091, A2 => n36487, B1 => n30616, B2 => 
                           n36803, ZN => n36471);
   U1478 : INV_X1 port map( A => n36471, ZN => n2843);
   U1479 : OAI22_X1 port map( A1 => n30091, A2 => n36472, B1 => n30615, B2 => 
                           n36803, ZN => n36473);
   U1480 : INV_X1 port map( A => n36473, ZN => n2903);
   U1481 : OAI22_X1 port map( A1 => n30115, A2 => n36783, B1 => n30298, B2 => 
                           n36799, ZN => n36474);
   U1482 : INV_X1 port map( A => n36474, ZN => n3163);
   U1483 : OAI22_X1 port map( A1 => n30095, A2 => n36487, B1 => n30608, B2 => 
                           n36807, ZN => n36475);
   U1484 : INV_X1 port map( A => n36475, ZN => n2842);
   U1485 : OAI22_X1 port map( A1 => n30091, A2 => n36748, B1 => n30612, B2 => 
                           n36803, ZN => n36476);
   U1486 : INV_X1 port map( A => n36476, ZN => n3106);
   U1487 : OAI22_X1 port map( A1 => n30115, A2 => n36477, B1 => n30324, B2 => 
                           n36799, ZN => n36478);
   U1488 : INV_X1 port map( A => n36478, ZN => n2854);
   U1489 : OAI22_X1 port map( A1 => n30095, A2 => n36662, B1 => n30611, B2 => 
                           n36807, ZN => n36479);
   U1490 : INV_X1 port map( A => n36479, ZN => n2978);
   U1491 : OAI22_X1 port map( A1 => n30115, A2 => n36718, B1 => n30337, B2 => 
                           n36799, ZN => n36480);
   U1492 : INV_X1 port map( A => n36480, ZN => n2938);
   U1493 : OAI22_X1 port map( A1 => n30095, A2 => n36730, B1 => n30603, B2 => 
                           n36807, ZN => n36481);
   U1494 : INV_X1 port map( A => n36481, ZN => n2808);
   U1495 : OAI22_X1 port map( A1 => n30091, A2 => n36662, B1 => n30613, B2 => 
                           n36803, ZN => n36482);
   U1496 : INV_X1 port map( A => n36482, ZN => n2979);
   U1497 : OAI22_X1 port map( A1 => n30115, A2 => n36692, B1 => n30331, B2 => 
                           n36799, ZN => n36483);
   U1498 : INV_X1 port map( A => n36483, ZN => n2950);
   U1499 : OAI22_X1 port map( A1 => n30115, A2 => n36683, B1 => n30313, B2 => 
                           n36799, ZN => n36484);
   U1500 : INV_X1 port map( A => n36484, ZN => n3034);
   U1501 : OAI22_X1 port map( A1 => n30115, A2 => n36485, B1 => n30308, B2 => 
                           n36799, ZN => n36486);
   U1502 : INV_X1 port map( A => n36486, ZN => n3194);
   U1503 : OAI22_X1 port map( A1 => n30100, A2 => n36487, B1 => n30714, B2 => 
                           n36805, ZN => n36488);
   U1504 : INV_X1 port map( A => n36488, ZN => n2847);
   U1505 : OAI22_X1 port map( A1 => n30115, A2 => n36489, B1 => n30378, B2 => 
                           n36799, ZN => n36490);
   U1506 : INV_X1 port map( A => n36490, ZN => n3444);
   U1507 : OAI22_X1 port map( A1 => n30104, A2 => n36730, B1 => n30710, B2 => 
                           n36811, ZN => n36491);
   U1508 : INV_X1 port map( A => n36491, ZN => n2815);
   U1509 : OAI22_X1 port map( A1 => n30095, A2 => n36718, B1 => n30599, B2 => 
                           n36807, ZN => n36492);
   U1510 : INV_X1 port map( A => n36492, ZN => n2944);
   U1511 : CLKBUF_X1 port map( A => n36493, Z => n36503);
   U1512 : OAI22_X1 port map( A1 => n30104, A2 => n36503, B1 => n31039, B2 => 
                           n36811, ZN => n36494);
   U1513 : INV_X1 port map( A => n36494, ZN => n3527);
   U1514 : OAI22_X1 port map( A1 => n30095, A2 => n36503, B1 => n31040, B2 => 
                           n36807, ZN => n36495);
   U1515 : INV_X1 port map( A => n36495, ZN => n3528);
   U1516 : OAI22_X1 port map( A1 => n30098, A2 => n36503, B1 => n31042, B2 => 
                           n36833, ZN => n36496);
   U1517 : INV_X1 port map( A => n36496, ZN => n3530);
   U1518 : OAI22_X1 port map( A1 => n30102, A2 => n36503, B1 => n31043, B2 => 
                           n36835, ZN => n36497);
   U1519 : INV_X1 port map( A => n36497, ZN => n3531);
   U1520 : OAI22_X1 port map( A1 => n30091, A2 => n36503, B1 => n31044, B2 => 
                           n36803, ZN => n36498);
   U1521 : INV_X1 port map( A => n36498, ZN => n3532);
   U1522 : OAI22_X1 port map( A1 => n30085, A2 => n36503, B1 => n30343, B2 => 
                           n36710, ZN => n36499);
   U1523 : INV_X1 port map( A => n36499, ZN => n3539);
   U1524 : OAI22_X1 port map( A1 => n30100, A2 => n36503, B1 => n31041, B2 => 
                           n36805, ZN => n36500);
   U1525 : INV_X1 port map( A => n36500, ZN => n3529);
   U1526 : OAI22_X1 port map( A1 => n30115, A2 => n36503, B1 => n30414, B2 => 
                           n36799, ZN => n36501);
   U1527 : INV_X1 port map( A => n36501, ZN => n3526);
   U1528 : OAI22_X1 port map( A1 => n30092, A2 => n36503, B1 => n31045, B2 => 
                           n36801, ZN => n36502);
   U1529 : INV_X1 port map( A => n36502, ZN => n3533);
   U1530 : OAI22_X1 port map( A1 => n30088, A2 => n36503, B1 => n30344, B2 => 
                           n36535, ZN => n36504);
   U1531 : INV_X1 port map( A => n36504, ZN => n3540);
   U1532 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31264, ZN => n36880);
   U1533 : CLKBUF_X1 port map( A => n36880, Z => n36866);
   U1534 : CLKBUF_X1 port map( A => n36505, Z => n36698);
   U1535 : OAI22_X1 port map( A1 => n30096, A2 => n36866, B1 => n30978, B2 => 
                           n36698, ZN => n36506);
   U1536 : INV_X1 port map( A => n36506, ZN => n2571);
   U1537 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31261, ZN => n36872);
   U1538 : OAI22_X1 port map( A1 => n30096, A2 => n36872, B1 => n30979, B2 => 
                           n36698, ZN => n36507);
   U1539 : INV_X1 port map( A => n36507, ZN => n2692);
   U1540 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31259, ZN => n36875);
   U1541 : CLKBUF_X1 port map( A => n36875, Z => n36896);
   U1542 : CLKBUF_X1 port map( A => n36508, Z => n36700);
   U1543 : OAI22_X1 port map( A1 => n30103, A2 => n36896, B1 => n30980, B2 => 
                           n36700, ZN => n36509);
   U1544 : INV_X1 port map( A => n36509, ZN => n2727);
   U1545 : OAI22_X1 port map( A1 => n30103, A2 => n36866, B1 => n30983, B2 => 
                           n36700, ZN => n36510);
   U1546 : INV_X1 port map( A => n36510, ZN => n2572);
   U1547 : CLKBUF_X1 port map( A => n36872, Z => n36894);
   U1548 : OAI22_X1 port map( A1 => n30090, A2 => n36894, B1 => n30985, B2 => 
                           n36511, ZN => n36512);
   U1549 : INV_X1 port map( A => n36512, ZN => n2662);
   U1550 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31262, ZN => n36887);
   U1551 : CLKBUF_X1 port map( A => n36887, Z => n36878);
   U1552 : OAI22_X1 port map( A1 => n30096, A2 => n36878, B1 => n30986, B2 => 
                           n36698, ZN => n36513);
   U1553 : INV_X1 port map( A => n36513, ZN => n2634);
   U1554 : CLKBUF_X1 port map( A => n36514, Z => n36676);
   U1555 : OAI22_X1 port map( A1 => n30101, A2 => n36515, B1 => n31086, B2 => 
                           n36676, ZN => n36516);
   U1556 : INV_X1 port map( A => n36516, ZN => n3330);
   U1557 : OAI22_X1 port map( A1 => n30103, A2 => n36878, B1 => n30987, B2 => 
                           n36700, ZN => n36517);
   U1558 : INV_X1 port map( A => n36517, ZN => n2635);
   U1559 : OAI22_X1 port map( A1 => n30090, A2 => n36878, B1 => n30988, B2 => 
                           n36511, ZN => n36518);
   U1560 : INV_X1 port map( A => n36518, ZN => n2636);
   U1561 : OAI22_X1 port map( A1 => n30112, A2 => n36887, B1 => n30974, B2 => 
                           n36519, ZN => n36520);
   U1562 : INV_X1 port map( A => n36520, ZN => n2661);
   U1563 : OAI22_X1 port map( A1 => n30090, A2 => n36715, B1 => n30173, B2 => 
                           n36511, ZN => n36521);
   U1564 : INV_X1 port map( A => n36521, ZN => n2864);
   U1565 : OAI22_X1 port map( A1 => n30089, A2 => n36783, B1 => n30175, B2 => 
                           n36522, ZN => n36523);
   U1566 : INV_X1 port map( A => n36523, ZN => n3151);
   U1567 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31265, ZN => n36884);
   U1568 : OAI22_X1 port map( A1 => n30112, A2 => n36884, B1 => n30141, B2 => 
                           n36519, ZN => n36524);
   U1569 : INV_X1 port map( A => n36524, ZN => n2548);
   U1570 : OAI22_X1 port map( A1 => n30107, A2 => n36584, B1 => n31008, B2 => 
                           n36525, ZN => n36526);
   U1571 : INV_X1 port map( A => n36526, ZN => n2890);
   U1572 : OAI22_X1 port map( A1 => n30112, A2 => n36875, B1 => n31004, B2 => 
                           n36519, ZN => n36527);
   U1573 : INV_X1 port map( A => n36527, ZN => n2734);
   U1574 : OAI22_X1 port map( A1 => n30096, A2 => n36896, B1 => n31003, B2 => 
                           n36698, ZN => n36528);
   U1575 : INV_X1 port map( A => n36528, ZN => n2733);
   U1576 : OAI22_X1 port map( A1 => n30090, A2 => n36896, B1 => n31001, B2 => 
                           n36511, ZN => n36529);
   U1577 : INV_X1 port map( A => n36529, ZN => n2731);
   U1578 : OAI22_X1 port map( A1 => n30112, A2 => n36894, B1 => n30992, B2 => 
                           n36519, ZN => n36530);
   U1579 : INV_X1 port map( A => n36530, ZN => n2665);
   U1580 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31258, ZN => n36889);
   U1581 : OAI22_X1 port map( A1 => n30089, A2 => n36889, B1 => n30148, B2 => 
                           n36522, ZN => n36531);
   U1582 : INV_X1 port map( A => n36531, ZN => n2769);
   U1583 : OAI22_X1 port map( A1 => n30103, A2 => n36894, B1 => n30991, B2 => 
                           n36700, ZN => n36532);
   U1584 : INV_X1 port map( A => n36532, ZN => n2664);
   U1585 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31260, ZN => n36863);
   U1586 : OAI22_X1 port map( A1 => n30089, A2 => n36863, B1 => n30150, B2 => 
                           n36522, ZN => n36533);
   U1587 : INV_X1 port map( A => n36533, ZN => n2705);
   U1588 : OAI22_X1 port map( A1 => n30089, A2 => n36718, B1 => n30181, B2 => 
                           n36522, ZN => n36534);
   U1589 : INV_X1 port map( A => n36534, ZN => n2929);
   U1590 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n31263, ZN => n36851);
   U1591 : CLKBUF_X1 port map( A => n36851, Z => n36892);
   U1592 : OAI22_X1 port map( A1 => n30088, A2 => n36892, B1 => n30188, B2 => 
                           n36535, ZN => n36536);
   U1593 : INV_X1 port map( A => n36536, ZN => n2611);
   U1594 : OAI22_X1 port map( A1 => n30089, A2 => n36851, B1 => n30151, B2 => 
                           n36522, ZN => n36537);
   U1595 : INV_X1 port map( A => n36537, ZN => n2609);
   U1596 : OAI22_X1 port map( A1 => n30108, A2 => n36584, B1 => n31015, B2 => 
                           n36538, ZN => n36539);
   U1597 : INV_X1 port map( A => n36539, ZN => n2892);
   U1598 : CLKBUF_X1 port map( A => n36863, Z => n36857);
   U1599 : OAI22_X1 port map( A1 => n30088, A2 => n36857, B1 => n30189, B2 => 
                           n36535, ZN => n36540);
   U1600 : INV_X1 port map( A => n36540, ZN => n2707);
   U1601 : CLKBUF_X1 port map( A => n36889, Z => n36870);
   U1602 : OAI22_X1 port map( A1 => n30088, A2 => n36870, B1 => n30190, B2 => 
                           n36535, ZN => n36541);
   U1603 : INV_X1 port map( A => n36541, ZN => n2771);
   U1604 : OAI22_X1 port map( A1 => n30088, A2 => n36872, B1 => n30566, B2 => 
                           n36535, ZN => n36542);
   U1605 : INV_X1 port map( A => n36542, ZN => n2679);
   U1606 : OAI22_X1 port map( A1 => n30087, A2 => n36875, B1 => n30535, B2 => 
                           n36543, ZN => n36544);
   U1607 : INV_X1 port map( A => n36544, ZN => n2738);
   U1608 : OAI22_X1 port map( A1 => n30087, A2 => n36887, B1 => n30533, B2 => 
                           n36543, ZN => n36545);
   U1609 : INV_X1 port map( A => n36545, ZN => n2640);
   U1610 : OAI22_X1 port map( A1 => n30087, A2 => n36880, B1 => n30532, B2 => 
                           n36543, ZN => n36546);
   U1611 : INV_X1 port map( A => n36546, ZN => n2577);
   U1612 : OAI22_X1 port map( A1 => n30090, A2 => n36863, B1 => n30282, B2 => 
                           n36511, ZN => n36547);
   U1613 : INV_X1 port map( A => n36547, ZN => n2715);
   U1614 : OAI22_X1 port map( A1 => n30090, A2 => n36851, B1 => n30283, B2 => 
                           n36511, ZN => n36548);
   U1615 : INV_X1 port map( A => n36548, ZN => n2619);
   U1616 : OAI22_X1 port map( A1 => n30108, A2 => n36887, B1 => n30540, B2 => 
                           n36538, ZN => n36549);
   U1617 : INV_X1 port map( A => n36549, ZN => n2642);
   U1618 : OAI22_X1 port map( A1 => n30106, A2 => n36875, B1 => n30527, B2 => 
                           n36550, ZN => n36551);
   U1619 : INV_X1 port map( A => n36551, ZN => n2737);
   U1620 : CLKBUF_X1 port map( A => n36884, Z => n36882);
   U1621 : OAI22_X1 port map( A1 => n30087, A2 => n36882, B1 => n30281, B2 => 
                           n36543, ZN => n36552);
   U1622 : INV_X1 port map( A => n36552, ZN => n2534);
   U1623 : OAI22_X1 port map( A1 => n30089, A2 => n36866, B1 => n30545, B2 => 
                           n36522, ZN => n36553);
   U1624 : INV_X1 port map( A => n36553, ZN => n2579);
   U1625 : OAI22_X1 port map( A1 => n30089, A2 => n36878, B1 => n30546, B2 => 
                           n36522, ZN => n36554);
   U1626 : INV_X1 port map( A => n36554, ZN => n2643);
   U1627 : OAI22_X1 port map( A1 => n30089, A2 => n36872, B1 => n30547, B2 => 
                           n36522, ZN => n36555);
   U1628 : INV_X1 port map( A => n36555, ZN => n2676);
   U1629 : OAI22_X1 port map( A1 => n30106, A2 => n36872, B1 => n30526, B2 => 
                           n36550, ZN => n36556);
   U1630 : INV_X1 port map( A => n36556, ZN => n2672);
   U1631 : OAI22_X1 port map( A1 => n30106, A2 => n36887, B1 => n30525, B2 => 
                           n36550, ZN => n36557);
   U1632 : INV_X1 port map( A => n36557, ZN => n2639);
   U1633 : OAI22_X1 port map( A1 => n30106, A2 => n36880, B1 => n30524, B2 => 
                           n36550, ZN => n36558);
   U1634 : INV_X1 port map( A => n36558, ZN => n2576);
   U1635 : OAI22_X1 port map( A1 => n30090, A2 => n36730, B1 => n30523, B2 => 
                           n36511, ZN => n36559);
   U1636 : INV_X1 port map( A => n36559, ZN => n2801);
   U1637 : OAI22_X1 port map( A1 => n30089, A2 => n36875, B1 => n30548, B2 => 
                           n36522, ZN => n36560);
   U1638 : INV_X1 port map( A => n36560, ZN => n2740);
   U1639 : OAI22_X1 port map( A1 => n30107, A2 => n36875, B1 => n30520, B2 => 
                           n36525, ZN => n36561);
   U1640 : INV_X1 port map( A => n36561, ZN => n2736);
   U1641 : OAI22_X1 port map( A1 => n30107, A2 => n36872, B1 => n30519, B2 => 
                           n36525, ZN => n36562);
   U1642 : INV_X1 port map( A => n36562, ZN => n2671);
   U1643 : OAI22_X1 port map( A1 => n30107, A2 => n36887, B1 => n30518, B2 => 
                           n36525, ZN => n36563);
   U1644 : INV_X1 port map( A => n36563, ZN => n2638);
   U1645 : OAI22_X1 port map( A1 => n30107, A2 => n36880, B1 => n30517, B2 => 
                           n36525, ZN => n36564);
   U1646 : INV_X1 port map( A => n36564, ZN => n2575);
   U1647 : OAI22_X1 port map( A1 => n30112, A2 => n36783, B1 => n30289, B2 => 
                           n36519, ZN => n36565);
   U1648 : INV_X1 port map( A => n36565, ZN => n3156);
   U1649 : OAI22_X1 port map( A1 => n30108, A2 => n36875, B1 => n30513, B2 => 
                           n36538, ZN => n36566);
   U1650 : INV_X1 port map( A => n36566, ZN => n2735);
   U1651 : OAI22_X1 port map( A1 => n30108, A2 => n36872, B1 => n30511, B2 => 
                           n36538, ZN => n36567);
   U1652 : INV_X1 port map( A => n36567, ZN => n2670);
   U1653 : OAI22_X1 port map( A1 => n30108, A2 => n36880, B1 => n30510, B2 => 
                           n36538, ZN => n36568);
   U1654 : INV_X1 port map( A => n36568, ZN => n2574);
   U1655 : OAI22_X1 port map( A1 => n30088, A2 => n36887, B1 => n30554, B2 => 
                           n36535, ZN => n36569);
   U1656 : INV_X1 port map( A => n36569, ZN => n2645);
   U1657 : OAI22_X1 port map( A1 => n30089, A2 => n36884, B1 => n30277, B2 => 
                           n36522, ZN => n36570);
   U1658 : INV_X1 port map( A => n36570, ZN => n2553);
   U1659 : OAI22_X1 port map( A1 => n30103, A2 => n36643, B1 => n30914, B2 => 
                           n36700, ZN => n36571);
   U1660 : INV_X1 port map( A => n36571, ZN => n3236);
   U1661 : CLKBUF_X1 port map( A => n36572, Z => n36687);
   U1662 : OAI22_X1 port map( A1 => n30099, A2 => n36870, B1 => n30889, B2 => 
                           n36687, ZN => n36573);
   U1663 : INV_X1 port map( A => n36573, ZN => n2765);
   U1664 : OAI22_X1 port map( A1 => n30088, A2 => n36880, B1 => n30561, B2 => 
                           n36535, ZN => n36574);
   U1665 : INV_X1 port map( A => n36574, ZN => n2581);
   U1666 : OAI22_X1 port map( A1 => n30088, A2 => n36751, B1 => n30562, B2 => 
                           n36535, ZN => n36575);
   U1667 : INV_X1 port map( A => n36575, ZN => n2804);
   U1668 : OAI22_X1 port map( A1 => n30101, A2 => n36870, B1 => n30886, B2 => 
                           n36676, ZN => n36576);
   U1669 : INV_X1 port map( A => n36576, ZN => n2763);
   U1670 : OAI22_X1 port map( A1 => n30107, A2 => n36715, B1 => n30501, B2 => 
                           n36525, ZN => n36577);
   U1671 : INV_X1 port map( A => n36577, ZN => n2878);
   U1672 : OAI22_X1 port map( A1 => n30103, A2 => n36870, B1 => n30884, B2 => 
                           n36700, ZN => n36578);
   U1673 : INV_X1 port map( A => n36578, ZN => n2761);
   U1674 : OAI22_X1 port map( A1 => n30099, A2 => n36579, B1 => n30883, B2 => 
                           n36687, ZN => n36580);
   U1675 : INV_X1 port map( A => n36580, ZN => n3016);
   U1676 : OAI22_X1 port map( A1 => n30088, A2 => n36875, B1 => n30567, B2 => 
                           n36535, ZN => n36581);
   U1677 : INV_X1 port map( A => n36581, ZN => n2743);
   U1678 : OAI22_X1 port map( A1 => n30106, A2 => n36884, B1 => n30497, B2 => 
                           n36550, ZN => n36582);
   U1679 : INV_X1 port map( A => n36582, ZN => n2558);
   U1680 : OAI22_X1 port map( A1 => n30107, A2 => n36643, B1 => n30496, B2 => 
                           n36525, ZN => n36583);
   U1681 : INV_X1 port map( A => n36583, ZN => n3223);
   U1682 : OAI22_X1 port map( A1 => n30087, A2 => n36584, B1 => n30571, B2 => 
                           n36543, ZN => n36585);
   U1683 : INV_X1 port map( A => n36585, ZN => n2899);
   U1684 : CLKBUF_X1 port map( A => n36586, Z => n36638);
   U1685 : OAI22_X1 port map( A1 => n30105, A2 => n36880, B1 => n30574, B2 => 
                           n36638, ZN => n36587);
   U1686 : INV_X1 port map( A => n36587, ZN => n2584);
   U1687 : OAI22_X1 port map( A1 => n30105, A2 => n36872, B1 => n30575, B2 => 
                           n36638, ZN => n36588);
   U1688 : INV_X1 port map( A => n36588, ZN => n2680);
   U1689 : OAI22_X1 port map( A1 => n30107, A2 => n36863, B1 => n30491, B2 => 
                           n36525, ZN => n36589);
   U1690 : INV_X1 port map( A => n36589, ZN => n2718);
   U1691 : OAI22_X1 port map( A1 => n30105, A2 => n36718, B1 => n30576, B2 => 
                           n36638, ZN => n36590);
   U1692 : INV_X1 port map( A => n36590, ZN => n2943);
   U1693 : OAI22_X1 port map( A1 => n30106, A2 => n36863, B1 => n30490, B2 => 
                           n36550, ZN => n36591);
   U1694 : INV_X1 port map( A => n36591, ZN => n2717);
   U1695 : OAI22_X1 port map( A1 => n30106, A2 => n36889, B1 => n30488, B2 => 
                           n36550, ZN => n36592);
   U1696 : INV_X1 port map( A => n36592, ZN => n2782);
   U1697 : OAI22_X1 port map( A1 => n30108, A2 => n36643, B1 => n30486, B2 => 
                           n36538, ZN => n36593);
   U1698 : INV_X1 port map( A => n36593, ZN => n3222);
   U1699 : OAI22_X1 port map( A1 => n30106, A2 => n36715, B1 => n30485, B2 => 
                           n36550, ZN => n36594);
   U1700 : INV_X1 port map( A => n36594, ZN => n2877);
   U1701 : OAI22_X1 port map( A1 => n30105, A2 => n36851, B1 => n30577, B2 => 
                           n36638, ZN => n36595);
   U1702 : INV_X1 port map( A => n36595, ZN => n2623);
   U1703 : OAI22_X1 port map( A1 => n30105, A2 => n36875, B1 => n30578, B2 => 
                           n36638, ZN => n36596);
   U1704 : INV_X1 port map( A => n36596, ZN => n2744);
   U1705 : OAI22_X1 port map( A1 => n30088, A2 => n36884, B1 => n30272, B2 => 
                           n36535, ZN => n36597);
   U1706 : INV_X1 port map( A => n36597, ZN => n2552);
   U1707 : OAI22_X1 port map( A1 => n30108, A2 => n36889, B1 => n30480, B2 => 
                           n36538, ZN => n36598);
   U1708 : INV_X1 port map( A => n36598, ZN => n2781);
   U1709 : OAI22_X1 port map( A1 => n30105, A2 => n36715, B1 => n30581, B2 => 
                           n36638, ZN => n36599);
   U1710 : INV_X1 port map( A => n36599, ZN => n2879);
   U1711 : OAI22_X1 port map( A1 => n30105, A2 => n36643, B1 => n30582, B2 => 
                           n36638, ZN => n36600);
   U1712 : INV_X1 port map( A => n36600, ZN => n3224);
   U1713 : OAI22_X1 port map( A1 => n30105, A2 => n36889, B1 => n30584, B2 => 
                           n36638, ZN => n36601);
   U1714 : INV_X1 port map( A => n36601, ZN => n2783);
   U1715 : OAI22_X1 port map( A1 => n30106, A2 => n36683, B1 => n30479, B2 => 
                           n36550, ZN => n36602);
   U1716 : INV_X1 port map( A => n36602, ZN => n3039);
   U1717 : OAI22_X1 port map( A1 => n30105, A2 => n36863, B1 => n30585, B2 => 
                           n36638, ZN => n36603);
   U1718 : INV_X1 port map( A => n36603, ZN => n2719);
   U1719 : OAI22_X1 port map( A1 => n30105, A2 => n36887, B1 => n30589, B2 => 
                           n36638, ZN => n36604);
   U1720 : INV_X1 port map( A => n36604, ZN => n2648);
   U1721 : OAI22_X1 port map( A1 => n30107, A2 => n36884, B1 => n30478, B2 => 
                           n36525, ZN => n36605);
   U1722 : INV_X1 port map( A => n36605, ZN => n2557);
   U1723 : CLKBUF_X1 port map( A => n36606, Z => n36696);
   U1724 : OAI22_X1 port map( A1 => n30093, A2 => n36889, B1 => n30869, B2 => 
                           n36696, ZN => n36607);
   U1725 : INV_X1 port map( A => n36607, ZN => n2788);
   U1726 : OAI22_X1 port map( A1 => n30107, A2 => n36851, B1 => n30476, B2 => 
                           n36525, ZN => n36608);
   U1727 : INV_X1 port map( A => n36608, ZN => n2622);
   U1728 : CLKBUF_X1 port map( A => n36609, Z => n36694);
   U1729 : OAI22_X1 port map( A1 => n30097, A2 => n36889, B1 => n30866, B2 => 
                           n36694, ZN => n36610);
   U1730 : INV_X1 port map( A => n36610, ZN => n2785);
   U1731 : OAI22_X1 port map( A1 => n30106, A2 => n36674, B1 => n30470, B2 => 
                           n36550, ZN => n36611);
   U1732 : INV_X1 port map( A => n36611, ZN => n3261);
   U1733 : OAI22_X1 port map( A1 => n30108, A2 => n36863, B1 => n30468, B2 => 
                           n36538, ZN => n36612);
   U1734 : INV_X1 port map( A => n36612, ZN => n2716);
   U1735 : OAI22_X1 port map( A1 => n30099, A2 => n36618, B1 => n30862, B2 => 
                           n36687, ZN => n36613);
   U1736 : INV_X1 port map( A => n36613, ZN => n2985);
   U1737 : OAI22_X1 port map( A1 => n30112, A2 => n36863, B1 => n30262, B2 => 
                           n36519, ZN => n36614);
   U1738 : INV_X1 port map( A => n36614, ZN => n2710);
   U1739 : OAI22_X1 port map( A1 => n30106, A2 => n36851, B1 => n30466, B2 => 
                           n36550, ZN => n36615);
   U1740 : INV_X1 port map( A => n36615, ZN => n2621);
   U1741 : OAI22_X1 port map( A1 => n30108, A2 => n36851, B1 => n30465, B2 => 
                           n36538, ZN => n36616);
   U1742 : INV_X1 port map( A => n36616, ZN => n2620);
   U1743 : OAI22_X1 port map( A1 => n30108, A2 => n36662, B1 => n30463, B2 => 
                           n36538, ZN => n36617);
   U1744 : INV_X1 port map( A => n36617, ZN => n2972);
   U1745 : OAI22_X1 port map( A1 => n30101, A2 => n36618, B1 => n30860, B2 => 
                           n36676, ZN => n36619);
   U1746 : INV_X1 port map( A => n36619, ZN => n2983);
   U1747 : OAI22_X1 port map( A1 => n30107, A2 => n36889, B1 => n30460, B2 => 
                           n36525, ZN => n36620);
   U1748 : INV_X1 port map( A => n36620, ZN => n2780);
   U1749 : OAI22_X1 port map( A1 => n30108, A2 => n36884, B1 => n30459, B2 => 
                           n36538, ZN => n36621);
   U1750 : INV_X1 port map( A => n36621, ZN => n2556);
   U1751 : OAI22_X1 port map( A1 => n30088, A2 => n36643, B1 => n30458, B2 => 
                           n36535, ZN => n36622);
   U1752 : INV_X1 port map( A => n36622, ZN => n3220);
   U1753 : OAI22_X1 port map( A1 => n30089, A2 => n36643, B1 => n30456, B2 => 
                           n36522, ZN => n36623);
   U1754 : INV_X1 port map( A => n36623, ZN => n3218);
   U1755 : OAI22_X1 port map( A1 => n30090, A2 => n36884, B1 => n30300, B2 => 
                           n36511, ZN => n36624);
   U1756 : INV_X1 port map( A => n36624, ZN => n2555);
   U1757 : OAI22_X1 port map( A1 => n30090, A2 => n36643, B1 => n30453, B2 => 
                           n36511, ZN => n36625);
   U1758 : INV_X1 port map( A => n36625, ZN => n3215);
   U1759 : OAI22_X1 port map( A1 => n30099, A2 => n36643, B1 => n30846, B2 => 
                           n36687, ZN => n36626);
   U1760 : INV_X1 port map( A => n36626, ZN => n3234);
   U1761 : OAI22_X1 port map( A1 => n30112, A2 => n36851, B1 => n30256, B2 => 
                           n36519, ZN => n36627);
   U1762 : INV_X1 port map( A => n36627, ZN => n2615);
   U1763 : OAI22_X1 port map( A1 => n30101, A2 => n36875, B1 => n30842, B2 => 
                           n36676, ZN => n36628);
   U1764 : INV_X1 port map( A => n36628, ZN => n2753);
   U1765 : OAI22_X1 port map( A1 => n30096, A2 => n36715, B1 => n30822, B2 => 
                           n36698, ZN => n36629);
   U1766 : INV_X1 port map( A => n36629, ZN => n2880);
   U1767 : OAI22_X1 port map( A1 => n30097, A2 => n36875, B1 => n30821, B2 => 
                           n36694, ZN => n36630);
   U1768 : INV_X1 port map( A => n36630, ZN => n2752);
   U1769 : OAI22_X1 port map( A1 => n30099, A2 => n36875, B1 => n30819, B2 => 
                           n36687, ZN => n36631);
   U1770 : INV_X1 port map( A => n36631, ZN => n2750);
   U1771 : OAI22_X1 port map( A1 => n30103, A2 => n36857, B1 => n30744, B2 => 
                           n36700, ZN => n36632);
   U1772 : INV_X1 port map( A => n36632, ZN => n2699);
   U1773 : OAI22_X1 port map( A1 => n30093, A2 => n36887, B1 => n30735, B2 => 
                           n36696, ZN => n36633);
   U1774 : INV_X1 port map( A => n36633, ZN => n2655);
   U1775 : OAI22_X1 port map( A1 => n30103, A2 => n36884, B1 => n30791, B2 => 
                           n36700, ZN => n36634);
   U1776 : INV_X1 port map( A => n36634, ZN => n2561);
   U1777 : OAI22_X1 port map( A1 => n30093, A2 => n36875, B1 => n30690, B2 => 
                           n36696, ZN => n36635);
   U1778 : INV_X1 port map( A => n36635, ZN => n2746);
   U1779 : OAI22_X1 port map( A1 => n30087, A2 => n36892, B1 => n30228, B2 => 
                           n36543, ZN => n36636);
   U1780 : INV_X1 port map( A => n36636, ZN => n2613);
   U1781 : OAI22_X1 port map( A1 => n30099, A2 => n36857, B1 => n30711, B2 => 
                           n36687, ZN => n36637);
   U1782 : INV_X1 port map( A => n36637, ZN => n2697);
   U1783 : OAI22_X1 port map( A1 => n30105, A2 => n36884, B1 => n30593, B2 => 
                           n36638, ZN => n36639);
   U1784 : INV_X1 port map( A => n36639, ZN => n2559);
   U1785 : OAI22_X1 port map( A1 => n30101, A2 => n36882, B1 => n30808, B2 => 
                           n36676, ZN => n36640);
   U1786 : INV_X1 port map( A => n36640, ZN => n2541);
   U1787 : OAI22_X1 port map( A1 => n30101, A2 => n36880, B1 => n30807, B2 => 
                           n36676, ZN => n36641);
   U1788 : INV_X1 port map( A => n36641, ZN => n2594);
   U1789 : OAI22_X1 port map( A1 => n30101, A2 => n36892, B1 => n30806, B2 => 
                           n36676, ZN => n36642);
   U1790 : INV_X1 port map( A => n36642, ZN => n2600);
   U1791 : OAI22_X1 port map( A1 => n30093, A2 => n36643, B1 => n30685, B2 => 
                           n36696, ZN => n36644);
   U1792 : INV_X1 port map( A => n36644, ZN => n3228);
   U1793 : OAI22_X1 port map( A1 => n30101, A2 => n36887, B1 => n30805, B2 => 
                           n36676, ZN => n36645);
   U1794 : INV_X1 port map( A => n36645, ZN => n2658);
   U1795 : OAI22_X1 port map( A1 => n30096, A2 => n36718, B1 => n30600, B2 => 
                           n36698, ZN => n36646);
   U1796 : INV_X1 port map( A => n36646, ZN => n2945);
   U1797 : OAI22_X1 port map( A1 => n30101, A2 => n36872, B1 => n30804, B2 => 
                           n36676, ZN => n36647);
   U1798 : INV_X1 port map( A => n36647, ZN => n2690);
   U1799 : OAI22_X1 port map( A1 => n30090, A2 => n36889, B1 => n30242, B2 => 
                           n36511, ZN => n36648);
   U1800 : INV_X1 port map( A => n36648, ZN => n2776);
   U1801 : OAI22_X1 port map( A1 => n30099, A2 => n36882, B1 => n30802, B2 => 
                           n36687, ZN => n36649);
   U1802 : INV_X1 port map( A => n36649, ZN => n2539);
   U1803 : OAI22_X1 port map( A1 => n30097, A2 => n36882, B1 => n30801, B2 => 
                           n36694, ZN => n36650);
   U1804 : INV_X1 port map( A => n36650, ZN => n2538);
   U1805 : OAI22_X1 port map( A1 => n30096, A2 => n36882, B1 => n30800, B2 => 
                           n36698, ZN => n36651);
   U1806 : INV_X1 port map( A => n36651, ZN => n2537);
   U1807 : OAI22_X1 port map( A1 => n30112, A2 => n36889, B1 => n30240, B2 => 
                           n36519, ZN => n36652);
   U1808 : INV_X1 port map( A => n36652, ZN => n2774);
   U1809 : OAI22_X1 port map( A1 => n30097, A2 => n36718, B1 => n30601, B2 => 
                           n36694, ZN => n36653);
   U1810 : INV_X1 port map( A => n36653, ZN => n2946);
   U1811 : OAI22_X1 port map( A1 => n30112, A2 => n36674, B1 => n30239, B2 => 
                           n36519, ZN => n36654);
   U1812 : INV_X1 port map( A => n36654, ZN => n3259);
   U1813 : OAI22_X1 port map( A1 => n30097, A2 => n36857, B1 => n30709, B2 => 
                           n36694, ZN => n36655);
   U1814 : INV_X1 port map( A => n36655, ZN => n2696);
   U1815 : OAI22_X1 port map( A1 => n30097, A2 => n36887, B1 => n30728, B2 => 
                           n36694, ZN => n36656);
   U1816 : INV_X1 port map( A => n36656, ZN => n2651);
   U1817 : OAI22_X1 port map( A1 => n30099, A2 => n36887, B1 => n30729, B2 => 
                           n36687, ZN => n36657);
   U1818 : INV_X1 port map( A => n36657, ZN => n2652);
   U1819 : OAI22_X1 port map( A1 => n30093, A2 => n36884, B1 => n30797, B2 => 
                           n36696, ZN => n36658);
   U1820 : INV_X1 port map( A => n36658, ZN => n2565);
   U1821 : OAI22_X1 port map( A1 => n30096, A2 => n36857, B1 => n30708, B2 => 
                           n36698, ZN => n36659);
   U1822 : INV_X1 port map( A => n36659, ZN => n2695);
   U1823 : OAI22_X1 port map( A1 => n30101, A2 => n36857, B1 => n30794, B2 => 
                           n36676, ZN => n36660);
   U1824 : INV_X1 port map( A => n36660, ZN => n2701);
   U1825 : OAI22_X1 port map( A1 => n30087, A2 => n36674, B1 => n30210, B2 => 
                           n36543, ZN => n36661);
   U1826 : INV_X1 port map( A => n36661, ZN => n3250);
   U1827 : OAI22_X1 port map( A1 => n30097, A2 => n36662, B1 => n30610, B2 => 
                           n36694, ZN => n36663);
   U1828 : INV_X1 port map( A => n36663, ZN => n2977);
   U1829 : OAI22_X1 port map( A1 => n30087, A2 => n36889, B1 => n30220, B2 => 
                           n36543, ZN => n36664);
   U1830 : INV_X1 port map( A => n36664, ZN => n2773);
   U1831 : OAI22_X1 port map( A1 => n30093, A2 => n36863, B1 => n30705, B2 => 
                           n36696, ZN => n36665);
   U1832 : INV_X1 port map( A => n36665, ZN => n2723);
   U1833 : OAI22_X1 port map( A1 => n30088, A2 => n36677, B1 => n30207, B2 => 
                           n36535, ZN => n36666);
   U1834 : INV_X1 port map( A => n36666, ZN => n3059);
   U1835 : OAI22_X1 port map( A1 => n30112, A2 => n36866, B1 => n30970, B2 => 
                           n36519, ZN => n36667);
   U1836 : INV_X1 port map( A => n36667, ZN => n2569);
   U1837 : OAI22_X1 port map( A1 => n30097, A2 => n36674, B1 => n30637, B2 => 
                           n36694, ZN => n36668);
   U1838 : INV_X1 port map( A => n36668, ZN => n3264);
   U1839 : OAI22_X1 port map( A1 => n30090, A2 => n36880, B1 => n30963, B2 => 
                           n36511, ZN => n36669);
   U1840 : INV_X1 port map( A => n36669, ZN => n2596);
   U1841 : OAI22_X1 port map( A1 => n30093, A2 => n36718, B1 => n30633, B2 => 
                           n36696, ZN => n36670);
   U1842 : INV_X1 port map( A => n36670, ZN => n2949);
   U1843 : OAI22_X1 port map( A1 => n30097, A2 => n36872, B1 => n30737, B2 => 
                           n36694, ZN => n36671);
   U1844 : INV_X1 port map( A => n36671, ZN => n2682);
   U1845 : OAI22_X1 port map( A1 => n30099, A2 => n36880, B1 => n30751, B2 => 
                           n36687, ZN => n36672);
   U1846 : INV_X1 port map( A => n36672, ZN => n2590);
   U1847 : OAI22_X1 port map( A1 => n30103, A2 => n36892, B1 => n30766, B2 => 
                           n36700, ZN => n36673);
   U1848 : INV_X1 port map( A => n36673, ZN => n2604);
   U1849 : OAI22_X1 port map( A1 => n30096, A2 => n36674, B1 => n30641, B2 => 
                           n36698, ZN => n36675);
   U1850 : INV_X1 port map( A => n36675, ZN => n3268);
   U1851 : OAI22_X1 port map( A1 => n30101, A2 => n36677, B1 => n30785, B2 => 
                           n36676, ZN => n36678);
   U1852 : INV_X1 port map( A => n36678, ZN => n3047);
   U1853 : OAI22_X1 port map( A1 => n30087, A2 => n36857, B1 => n30208, B2 => 
                           n36543, ZN => n36679);
   U1854 : INV_X1 port map( A => n36679, ZN => n2708);
   U1855 : OAI22_X1 port map( A1 => n30096, A2 => n36889, B1 => n30618, B2 => 
                           n36698, ZN => n36680);
   U1856 : INV_X1 port map( A => n36680, ZN => n2784);
   U1857 : OAI22_X1 port map( A1 => n30087, A2 => n36872, B1 => n30534, B2 => 
                           n36543, ZN => n36681);
   U1858 : INV_X1 port map( A => n36681, ZN => n2673);
   U1859 : OAI22_X1 port map( A1 => n30099, A2 => n36872, B1 => n30738, B2 => 
                           n36687, ZN => n36682);
   U1860 : INV_X1 port map( A => n36682, ZN => n2683);
   U1861 : OAI22_X1 port map( A1 => n30087, A2 => n36683, B1 => n30223, B2 => 
                           n36543, ZN => n36684);
   U1862 : INV_X1 port map( A => n36684, ZN => n3029);
   U1863 : OAI22_X1 port map( A1 => n30112, A2 => n36715, B1 => n30325, B2 => 
                           n36519, ZN => n36685);
   U1864 : INV_X1 port map( A => n36685, ZN => n2874);
   U1865 : OAI22_X1 port map( A1 => n30093, A2 => n36872, B1 => n30742, B2 => 
                           n36696, ZN => n36686);
   U1866 : INV_X1 port map( A => n36686, ZN => n2687);
   U1867 : OAI22_X1 port map( A1 => n30099, A2 => n36851, B1 => n30763, B2 => 
                           n36687, ZN => n36688);
   U1868 : INV_X1 port map( A => n36688, ZN => n2629);
   U1869 : OAI22_X1 port map( A1 => n30097, A2 => n36851, B1 => n30762, B2 => 
                           n36694, ZN => n36689);
   U1870 : INV_X1 port map( A => n36689, ZN => n2628);
   U1871 : OAI22_X1 port map( A1 => n30093, A2 => n36880, B1 => n30746, B2 => 
                           n36696, ZN => n36690);
   U1872 : INV_X1 port map( A => n36690, ZN => n2586);
   U1873 : OAI22_X1 port map( A1 => n30093, A2 => n36730, B1 => n30636, B2 => 
                           n36696, ZN => n36691);
   U1874 : INV_X1 port map( A => n36691, ZN => n2813);
   U1875 : OAI22_X1 port map( A1 => n30103, A2 => n36692, B1 => n30756, B2 => 
                           n36700, ZN => n36693);
   U1876 : INV_X1 port map( A => n36693, ZN => n2954);
   U1877 : OAI22_X1 port map( A1 => n30097, A2 => n36880, B1 => n30750, B2 => 
                           n36694, ZN => n36695);
   U1878 : INV_X1 port map( A => n36695, ZN => n2589);
   U1879 : OAI22_X1 port map( A1 => n30093, A2 => n36851, B1 => n30758, B2 => 
                           n36696, ZN => n36697);
   U1880 : INV_X1 port map( A => n36697, ZN => n2624);
   U1881 : OAI22_X1 port map( A1 => n30096, A2 => n36851, B1 => n30761, B2 => 
                           n36698, ZN => n36699);
   U1882 : INV_X1 port map( A => n36699, ZN => n2627);
   U1883 : OAI22_X1 port map( A1 => n30103, A2 => n36701, B1 => n30755, B2 => 
                           n36700, ZN => n36702);
   U1884 : INV_X1 port map( A => n36702, ZN => n2922);
   U1885 : OAI22_X1 port map( A1 => n30123, A2 => n36889, B1 => n31163, B2 => 
                           n36703, ZN => n36704);
   U1886 : INV_X1 port map( A => n36704, ZN => n2767);
   U1887 : OAI22_X1 port map( A1 => n30120, A2 => n36718, B1 => n30334, B2 => 
                           n36705, ZN => n36706);
   U1888 : INV_X1 port map( A => n36706, ZN => n2936);
   U1889 : OAI22_X1 port map( A1 => n30123, A2 => n36783, B1 => n30294, B2 => 
                           n36703, ZN => n36707);
   U1890 : INV_X1 port map( A => n36707, ZN => n3159);
   U1891 : OAI22_X1 port map( A1 => n30117, A2 => n36718, B1 => n30335, B2 => 
                           n36708, ZN => n36709);
   U1892 : INV_X1 port map( A => n36709, ZN => n2937);
   U1893 : OAI22_X1 port map( A1 => n30085, A2 => n36884, B1 => n30292, B2 => 
                           n36710, ZN => n36711);
   U1894 : INV_X1 port map( A => n36711, ZN => n2554);
   U1895 : OAI22_X1 port map( A1 => n30117, A2 => n36712, B1 => n30287, B2 => 
                           n36708, ZN => n36713);
   U1896 : INV_X1 port map( A => n36713, ZN => n3132);
   U1897 : OAI22_X1 port map( A1 => n30124, A2 => n36715, B1 => n30317, B2 => 
                           n36714, ZN => n36716);
   U1898 : INV_X1 port map( A => n36716, ZN => n2869);
   U1899 : OAI22_X1 port map( A1 => n30116, A2 => n36718, B1 => n30321, B2 => 
                           n36717, ZN => n36719);
   U1900 : INV_X1 port map( A => n36719, ZN => n2935);
   U1901 : OAI22_X1 port map( A1 => n30117, A2 => n36889, B1 => n30243, B2 => 
                           n36708, ZN => n36720);
   U1902 : INV_X1 port map( A => n36720, ZN => n2777);
   U1903 : OAI22_X1 port map( A1 => n30117, A2 => n36878, B1 => n30981, B2 => 
                           n36708, ZN => n36721);
   U1904 : INV_X1 port map( A => n36721, ZN => n2632);
   U1905 : OAI22_X1 port map( A1 => n30120, A2 => n36878, B1 => n30982, B2 => 
                           n36705, ZN => n36722);
   U1906 : INV_X1 port map( A => n36722, ZN => n2633);
   U1907 : OAI22_X1 port map( A1 => n30120, A2 => n36870, B1 => n30244, B2 => 
                           n36705, ZN => n36723);
   U1908 : INV_X1 port map( A => n36723, ZN => n2758);
   U1909 : OAI22_X1 port map( A1 => n30116, A2 => n36878, B1 => n30976, B2 => 
                           n36717, ZN => n36724);
   U1910 : INV_X1 port map( A => n36724, ZN => n2631);
   U1911 : OAI22_X1 port map( A1 => n30120, A2 => n36875, B1 => n30949, B2 => 
                           n36705, ZN => n36725);
   U1912 : INV_X1 port map( A => n36725, ZN => n2756);
   U1913 : OAI22_X1 port map( A1 => n30109, A2 => n36889, B1 => n30245, B2 => 
                           n36726, ZN => n36727);
   U1914 : INV_X1 port map( A => n36727, ZN => n2778);
   U1915 : OAI22_X1 port map( A1 => n30116, A2 => n36788, B1 => n30950, B2 => 
                           n36717, ZN => n36728);
   U1916 : INV_X1 port map( A => n36728, ZN => n2823);
   U1917 : OAI22_X1 port map( A1 => n30116, A2 => n36889, B1 => n30246, B2 => 
                           n36717, ZN => n36729);
   U1918 : INV_X1 port map( A => n36729, ZN => n2779);
   U1919 : OAI22_X1 port map( A1 => n30109, A2 => n36730, B1 => n30941, B2 => 
                           n36726, ZN => n36731);
   U1920 : INV_X1 port map( A => n36731, ZN => n2820);
   U1921 : OAI22_X1 port map( A1 => n30109, A2 => n36851, B1 => n30255, B2 => 
                           n36726, ZN => n36732);
   U1922 : INV_X1 port map( A => n36732, ZN => n2614);
   U1923 : OAI22_X1 port map( A1 => n30109, A2 => n36866, B1 => n30973, B2 => 
                           n36726, ZN => n36733);
   U1924 : INV_X1 port map( A => n36733, ZN => n2570);
   U1925 : OAI22_X1 port map( A1 => n30120, A2 => n36788, B1 => n30953, B2 => 
                           n36705, ZN => n36734);
   U1926 : INV_X1 port map( A => n36734, ZN => n2825);
   U1927 : OAI22_X1 port map( A1 => n30109, A2 => n36894, B1 => n30990, B2 => 
                           n36726, ZN => n36735);
   U1928 : INV_X1 port map( A => n36735, ZN => n2663);
   U1929 : OAI22_X1 port map( A1 => n30086, A2 => n36884, B1 => n30258, B2 => 
                           n36736, ZN => n36737);
   U1930 : INV_X1 port map( A => n36737, ZN => n2551);
   U1931 : OAI22_X1 port map( A1 => n30116, A2 => n36851, B1 => n30259, B2 => 
                           n36717, ZN => n36738);
   U1932 : INV_X1 port map( A => n36738, ZN => n2617);
   U1933 : OAI22_X1 port map( A1 => n30086, A2 => n36863, B1 => n30227, B2 => 
                           n36736, ZN => n36739);
   U1934 : INV_X1 port map( A => n36739, ZN => n2709);
   U1935 : OAI22_X1 port map( A1 => n30117, A2 => n36851, B1 => n30260, B2 => 
                           n36708, ZN => n36740);
   U1936 : INV_X1 port map( A => n36740, ZN => n2606);
   U1937 : OAI22_X1 port map( A1 => n30120, A2 => n36851, B1 => n30261, B2 => 
                           n36705, ZN => n36741);
   U1938 : INV_X1 port map( A => n36741, ZN => n2618);
   U1939 : OAI22_X1 port map( A1 => n30109, A2 => n36863, B1 => n30263, B2 => 
                           n36726, ZN => n36742);
   U1940 : INV_X1 port map( A => n36742, ZN => n2711);
   U1941 : OAI22_X1 port map( A1 => n30117, A2 => n36875, B1 => n30959, B2 => 
                           n36708, ZN => n36743);
   U1942 : INV_X1 port map( A => n36743, ZN => n2757);
   U1943 : OAI22_X1 port map( A1 => n30085, A2 => n36851, B1 => n30163, B2 => 
                           n36710, ZN => n36744);
   U1944 : INV_X1 port map( A => n36744, ZN => n2610);
   U1945 : OAI22_X1 port map( A1 => n30085, A2 => n36863, B1 => n30156, B2 => 
                           n36710, ZN => n36745);
   U1946 : INV_X1 port map( A => n36745, ZN => n2706);
   U1947 : OAI22_X1 port map( A1 => n30085, A2 => n36870, B1 => n30155, B2 => 
                           n36710, ZN => n36746);
   U1948 : INV_X1 port map( A => n36746, ZN => n2770);
   U1949 : OAI22_X1 port map( A1 => n30109, A2 => n36748, B1 => n30266, B2 => 
                           n36726, ZN => n36747);
   U1950 : INV_X1 port map( A => n36747, ZN => n3095);
   U1951 : OAI22_X1 port map( A1 => n30085, A2 => n36748, B1 => n30153, B2 => 
                           n36710, ZN => n36749);
   U1952 : INV_X1 port map( A => n36749, ZN => n3087);
   U1953 : OAI22_X1 port map( A1 => n30124, A2 => n36751, B1 => n30960, B2 => 
                           n36714, ZN => n36750);
   U1954 : INV_X1 port map( A => n36750, ZN => n2794);
   U1955 : OAI22_X1 port map( A1 => n30123, A2 => n36751, B1 => n30964, B2 => 
                           n36703, ZN => n36752);
   U1956 : INV_X1 port map( A => n36752, ZN => n2795);
   U1957 : OAI22_X1 port map( A1 => n30116, A2 => n36894, B1 => n30995, B2 => 
                           n36717, ZN => n36753);
   U1958 : INV_X1 port map( A => n36753, ZN => n2667);
   U1959 : OAI22_X1 port map( A1 => n30124, A2 => n36884, B1 => n30145, B2 => 
                           n36714, ZN => n36754);
   U1960 : INV_X1 port map( A => n36754, ZN => n2550);
   U1961 : OAI22_X1 port map( A1 => n30116, A2 => n36896, B1 => n30996, B2 => 
                           n36717, ZN => n36755);
   U1962 : INV_X1 port map( A => n36755, ZN => n2728);
   U1963 : OAI22_X1 port map( A1 => n30085, A2 => n36783, B1 => n30217, B2 => 
                           n36710, ZN => n36756);
   U1964 : INV_X1 port map( A => n36756, ZN => n3154);
   U1965 : OAI22_X1 port map( A1 => n30123, A2 => n36863, B1 => n30144, B2 => 
                           n36703, ZN => n36757);
   U1966 : INV_X1 port map( A => n36757, ZN => n2704);
   U1967 : OAI22_X1 port map( A1 => n30120, A2 => n36894, B1 => n30997, B2 => 
                           n36705, ZN => n36758);
   U1968 : INV_X1 port map( A => n36758, ZN => n2668);
   U1969 : OAI22_X1 port map( A1 => n30124, A2 => n36889, B1 => n30143, B2 => 
                           n36714, ZN => n36759);
   U1970 : INV_X1 port map( A => n36759, ZN => n2768);
   U1971 : OAI22_X1 port map( A1 => n30086, A2 => n36851, B1 => n30215, B2 => 
                           n36736, ZN => n36760);
   U1972 : INV_X1 port map( A => n36760, ZN => n2612);
   U1973 : OAI22_X1 port map( A1 => n30109, A2 => n36896, B1 => n30999, B2 => 
                           n36726, ZN => n36761);
   U1974 : INV_X1 port map( A => n36761, ZN => n2730);
   U1975 : OAI22_X1 port map( A1 => n30117, A2 => n36882, B1 => n30142, B2 => 
                           n36708, ZN => n36762);
   U1976 : INV_X1 port map( A => n36762, ZN => n2549);
   U1977 : OAI22_X1 port map( A1 => n30117, A2 => n36894, B1 => n31005, B2 => 
                           n36708, ZN => n36763);
   U1978 : INV_X1 port map( A => n36763, ZN => n2669);
   U1979 : OAI22_X1 port map( A1 => n30085, A2 => n36896, B1 => n30572, B2 => 
                           n36710, ZN => n36764);
   U1980 : INV_X1 port map( A => n36764, ZN => n2726);
   U1981 : OAI22_X1 port map( A1 => n30120, A2 => n36863, B1 => n30273, B2 => 
                           n36705, ZN => n36765);
   U1982 : INV_X1 port map( A => n36765, ZN => n2712);
   U1983 : OAI22_X1 port map( A1 => n30117, A2 => n36863, B1 => n30274, B2 => 
                           n36708, ZN => n36766);
   U1984 : INV_X1 port map( A => n36766, ZN => n2713);
   U1985 : OAI22_X1 port map( A1 => n30123, A2 => n36882, B1 => n30140, B2 => 
                           n36703, ZN => n36767);
   U1986 : INV_X1 port map( A => n36767, ZN => n2547);
   U1987 : OAI22_X1 port map( A1 => n30120, A2 => n36884, B1 => n30139, B2 => 
                           n36705, ZN => n36768);
   U1988 : INV_X1 port map( A => n36768, ZN => n2546);
   U1989 : OAI22_X1 port map( A1 => n30120, A2 => n36866, B1 => n30993, B2 => 
                           n36705, ZN => n36769);
   U1990 : INV_X1 port map( A => n36769, ZN => n2573);
   U1991 : OAI22_X1 port map( A1 => n30086, A2 => n36880, B1 => n30568, B2 => 
                           n36736, ZN => n36770);
   U1992 : INV_X1 port map( A => n36770, ZN => n2582);
   U1993 : OAI22_X1 port map( A1 => n30123, A2 => n36880, B1 => n30557, B2 => 
                           n36703, ZN => n36771);
   U1994 : INV_X1 port map( A => n36771, ZN => n2580);
   U1995 : OAI22_X1 port map( A1 => n30124, A2 => n36851, B1 => n30138, B2 => 
                           n36714, ZN => n36772);
   U1996 : INV_X1 port map( A => n36772, ZN => n2608);
   U1997 : OAI22_X1 port map( A1 => n30123, A2 => n36851, B1 => n30137, B2 => 
                           n36703, ZN => n36773);
   U1998 : INV_X1 port map( A => n36773, ZN => n2607);
   U1999 : OAI22_X1 port map( A1 => n30124, A2 => n36863, B1 => n30136, B2 => 
                           n36714, ZN => n36774);
   U2000 : INV_X1 port map( A => n36774, ZN => n2703);
   U2001 : OAI22_X1 port map( A1 => n30116, A2 => n36857, B1 => n30275, B2 => 
                           n36717, ZN => n36775);
   U2002 : INV_X1 port map( A => n36775, ZN => n2694);
   U2003 : OAI22_X1 port map( A1 => n30124, A2 => n36896, B1 => n30539, B2 => 
                           n36714, ZN => n36776);
   U2004 : INV_X1 port map( A => n36776, ZN => n2739);
   U2005 : OAI22_X1 port map( A1 => n30109, A2 => n36884, B1 => n30135, B2 => 
                           n36726, ZN => n36777);
   U2006 : INV_X1 port map( A => n36777, ZN => n2545);
   U2007 : OAI22_X1 port map( A1 => n30085, A2 => n36887, B1 => n30564, B2 => 
                           n36710, ZN => n36778);
   U2008 : INV_X1 port map( A => n36778, ZN => n2647);
   U2009 : OAI22_X1 port map( A1 => n30086, A2 => n36894, B1 => n30549, B2 => 
                           n36736, ZN => n36779);
   U2010 : INV_X1 port map( A => n36779, ZN => n2677);
   U2011 : OAI22_X1 port map( A1 => n30116, A2 => n36884, B1 => n30134, B2 => 
                           n36717, ZN => n36780);
   U2012 : INV_X1 port map( A => n36780, ZN => n2544);
   U2013 : OAI22_X1 port map( A1 => n30124, A2 => n36894, B1 => n30538, B2 => 
                           n36714, ZN => n36781);
   U2014 : INV_X1 port map( A => n36781, ZN => n2674);
   U2015 : OAI22_X1 port map( A1 => n30123, A2 => n36887, B1 => n30558, B2 => 
                           n36703, ZN => n36782);
   U2016 : INV_X1 port map( A => n36782, ZN => n2646);
   U2017 : OAI22_X1 port map( A1 => n30086, A2 => n36783, B1 => n30183, B2 => 
                           n36736, ZN => n36784);
   U2018 : INV_X1 port map( A => n36784, ZN => n3152);
   U2019 : OAI22_X1 port map( A1 => n30086, A2 => n36878, B1 => n30553, B2 => 
                           n36736, ZN => n36785);
   U2020 : INV_X1 port map( A => n36785, ZN => n2644);
   U2021 : OAI22_X1 port map( A1 => n30109, A2 => n36887, B1 => n30972, B2 => 
                           n36726, ZN => n36786);
   U2022 : INV_X1 port map( A => n36786, ZN => n2660);
   U2023 : OAI22_X1 port map( A1 => n30085, A2 => n36880, B1 => n30573, B2 => 
                           n36710, ZN => n36787);
   U2024 : INV_X1 port map( A => n36787, ZN => n2583);
   U2025 : OAI22_X1 port map( A1 => n30086, A2 => n36788, B1 => n30552, B2 => 
                           n36736, ZN => n36789);
   U2026 : INV_X1 port map( A => n36789, ZN => n2837);
   U2027 : OAI22_X1 port map( A1 => n30117, A2 => n36866, B1 => n30967, B2 => 
                           n36708, ZN => n36790);
   U2028 : INV_X1 port map( A => n36790, ZN => n2566);
   U2029 : OAI22_X1 port map( A1 => n30086, A2 => n36889, B1 => n30212, B2 => 
                           n36736, ZN => n36791);
   U2030 : INV_X1 port map( A => n36791, ZN => n2772);
   U2031 : OAI22_X1 port map( A1 => n30124, A2 => n36887, B1 => n30537, B2 => 
                           n36714, ZN => n36792);
   U2032 : INV_X1 port map( A => n36792, ZN => n2641);
   U2033 : OAI22_X1 port map( A1 => n30116, A2 => n36866, B1 => n30968, B2 => 
                           n36717, ZN => n36793);
   U2034 : INV_X1 port map( A => n36793, ZN => n2567);
   U2035 : OAI22_X1 port map( A1 => n30123, A2 => n36875, B1 => n30560, B2 => 
                           n36703, ZN => n36794);
   U2036 : INV_X1 port map( A => n36794, ZN => n2742);
   U2037 : OAI22_X1 port map( A1 => n30123, A2 => n36894, B1 => n30541, B2 => 
                           n36703, ZN => n36795);
   U2038 : INV_X1 port map( A => n36795, ZN => n2675);
   U2039 : OAI22_X1 port map( A1 => n30085, A2 => n36872, B1 => n30555, B2 => 
                           n36710, ZN => n36796);
   U2040 : INV_X1 port map( A => n36796, ZN => n2678);
   U2041 : OAI22_X1 port map( A1 => n30086, A2 => n36896, B1 => n30550, B2 => 
                           n36736, ZN => n36797);
   U2042 : INV_X1 port map( A => n36797, ZN => n2741);
   U2043 : OAI22_X1 port map( A1 => n30124, A2 => n36866, B1 => n30536, B2 => 
                           n36714, ZN => n36798);
   U2044 : INV_X1 port map( A => n36798, ZN => n2578);
   U2045 : OAI22_X1 port map( A1 => n30115, A2 => n36889, B1 => n30241, B2 => 
                           n36799, ZN => n36800);
   U2046 : INV_X1 port map( A => n36800, ZN => n2775);
   U2047 : OAI22_X1 port map( A1 => n30092, A2 => n36892, B1 => n30772, B2 => 
                           n36801, ZN => n36802);
   U2048 : INV_X1 port map( A => n36802, ZN => n2602);
   U2049 : OAI22_X1 port map( A1 => n30091, A2 => n36892, B1 => n30771, B2 => 
                           n36803, ZN => n36804);
   U2050 : INV_X1 port map( A => n36804, ZN => n2603);
   U2051 : OAI22_X1 port map( A1 => n30100, A2 => n36892, B1 => n30765, B2 => 
                           n36805, ZN => n36806);
   U2052 : INV_X1 port map( A => n36806, ZN => n2605);
   U2053 : OAI22_X1 port map( A1 => n30095, A2 => n36851, B1 => n30760, B2 => 
                           n36807, ZN => n36808);
   U2054 : INV_X1 port map( A => n36808, ZN => n2626);
   U2055 : OAI22_X1 port map( A1 => n30091, A2 => n36863, B1 => n30703, B2 => 
                           n36803, ZN => n36809);
   U2056 : INV_X1 port map( A => n36809, ZN => n2721);
   U2057 : OAI22_X1 port map( A1 => n30092, A2 => n36863, B1 => n30704, B2 => 
                           n36801, ZN => n36810);
   U2058 : INV_X1 port map( A => n36810, ZN => n2722);
   U2059 : OAI22_X1 port map( A1 => n30104, A2 => n36887, B1 => n30731, B2 => 
                           n36811, ZN => n36812);
   U2060 : INV_X1 port map( A => n36812, ZN => n2653);
   U2061 : CLKBUF_X1 port map( A => n36813, Z => n36855);
   U2062 : OAI22_X1 port map( A1 => n30094, A2 => n36863, B1 => n30706, B2 => 
                           n36855, ZN => n36814);
   U2063 : INV_X1 port map( A => n36814, ZN => n2724);
   U2064 : OAI22_X1 port map( A1 => n30091, A2 => n36887, B1 => n30733, B2 => 
                           n36803, ZN => n36815);
   U2065 : INV_X1 port map( A => n36815, ZN => n2654);
   U2066 : OAI22_X1 port map( A1 => n30095, A2 => n36863, B1 => n30707, B2 => 
                           n36807, ZN => n36816);
   U2067 : INV_X1 port map( A => n36816, ZN => n2725);
   U2068 : OAI22_X1 port map( A1 => n30094, A2 => n36851, B1 => n30759, B2 => 
                           n36855, ZN => n36817);
   U2069 : INV_X1 port map( A => n36817, ZN => n2625);
   U2070 : OAI22_X1 port map( A1 => n30095, A2 => n36872, B1 => n30736, B2 => 
                           n36807, ZN => n36818);
   U2071 : INV_X1 port map( A => n36818, ZN => n2681);
   U2072 : OAI22_X1 port map( A1 => n30100, A2 => n36872, B1 => n30739, B2 => 
                           n36805, ZN => n36819);
   U2073 : INV_X1 port map( A => n36819, ZN => n2684);
   U2074 : OAI22_X1 port map( A1 => n30100, A2 => n36880, B1 => n30754, B2 => 
                           n36805, ZN => n36820);
   U2075 : INV_X1 port map( A => n36820, ZN => n2592);
   U2076 : OAI22_X1 port map( A1 => n30091, A2 => n36880, B1 => n30753, B2 => 
                           n36803, ZN => n36821);
   U2077 : INV_X1 port map( A => n36821, ZN => n2591);
   U2078 : OAI22_X1 port map( A1 => n30095, A2 => n36887, B1 => n30723, B2 => 
                           n36807, ZN => n36822);
   U2079 : INV_X1 port map( A => n36822, ZN => n2650);
   U2080 : OAI22_X1 port map( A1 => n30100, A2 => n36887, B1 => n30752, B2 => 
                           n36805, ZN => n36823);
   U2081 : INV_X1 port map( A => n36823, ZN => n2656);
   U2082 : OAI22_X1 port map( A1 => n30104, A2 => n36872, B1 => n30740, B2 => 
                           n36811, ZN => n36824);
   U2083 : INV_X1 port map( A => n36824, ZN => n2685);
   U2084 : OAI22_X1 port map( A1 => n30091, A2 => n36872, B1 => n30741, B2 => 
                           n36803, ZN => n36825);
   U2085 : INV_X1 port map( A => n36825, ZN => n2686);
   U2086 : OAI22_X1 port map( A1 => n30094, A2 => n36887, B1 => n30722, B2 => 
                           n36855, ZN => n36826);
   U2087 : INV_X1 port map( A => n36826, ZN => n2649);
   U2088 : OAI22_X1 port map( A1 => n30095, A2 => n36880, B1 => n30749, B2 => 
                           n36807, ZN => n36827);
   U2089 : INV_X1 port map( A => n36827, ZN => n2588);
   U2090 : OAI22_X1 port map( A1 => n30094, A2 => n36880, B1 => n30748, B2 => 
                           n36855, ZN => n36828);
   U2091 : INV_X1 port map( A => n36828, ZN => n2587);
   U2092 : OAI22_X1 port map( A1 => n30104, A2 => n36875, B1 => n30747, B2 => 
                           n36811, ZN => n36829);
   U2093 : INV_X1 port map( A => n36829, ZN => n2749);
   U2094 : OAI22_X1 port map( A1 => n30104, A2 => n36880, B1 => n30745, B2 => 
                           n36811, ZN => n36830);
   U2095 : INV_X1 port map( A => n36830, ZN => n2585);
   U2096 : OAI22_X1 port map( A1 => n30094, A2 => n36872, B1 => n30743, B2 => 
                           n36855, ZN => n36831);
   U2097 : INV_X1 port map( A => n36831, ZN => n2688);
   U2098 : OAI22_X1 port map( A1 => n30091, A2 => n36884, B1 => n30795, B2 => 
                           n36803, ZN => n36832);
   U2099 : INV_X1 port map( A => n36832, ZN => n2563);
   U2100 : CLKBUF_X1 port map( A => n36833, Z => n36891);
   U2101 : OAI22_X1 port map( A1 => n30098, A2 => n36889, B1 => n30896, B2 => 
                           n36891, ZN => n36834);
   U2102 : INV_X1 port map( A => n36834, ZN => n2766);
   U2103 : OAI22_X1 port map( A1 => n30102, A2 => n36880, B1 => n30779, B2 => 
                           n36835, ZN => n36836);
   U2104 : INV_X1 port map( A => n36836, ZN => n2593);
   U2105 : OAI22_X1 port map( A1 => n30102, A2 => n36892, B1 => n30780, B2 => 
                           n36835, ZN => n36837);
   U2106 : INV_X1 port map( A => n36837, ZN => n2601);
   U2107 : OAI22_X1 port map( A1 => n30115, A2 => n36884, B1 => n30133, B2 => 
                           n36799, ZN => n36838);
   U2108 : INV_X1 port map( A => n36838, ZN => n2543);
   U2109 : OAI22_X1 port map( A1 => n30102, A2 => n36887, B1 => n30781, B2 => 
                           n36835, ZN => n36839);
   U2110 : INV_X1 port map( A => n36839, ZN => n2657);
   U2111 : OAI22_X1 port map( A1 => n30104, A2 => n36863, B1 => n30700, B2 => 
                           n36811, ZN => n36840);
   U2112 : INV_X1 port map( A => n36840, ZN => n2720);
   U2113 : OAI22_X1 port map( A1 => n30102, A2 => n36872, B1 => n30782, B2 => 
                           n36835, ZN => n36841);
   U2114 : INV_X1 port map( A => n36841, ZN => n2689);
   U2115 : OAI22_X1 port map( A1 => n30102, A2 => n36857, B1 => n30783, B2 => 
                           n36835, ZN => n36842);
   U2116 : INV_X1 port map( A => n36842, ZN => n2700);
   U2117 : OAI22_X1 port map( A1 => n30104, A2 => n36892, B1 => n30891, B2 => 
                           n36811, ZN => n36843);
   U2118 : INV_X1 port map( A => n36843, ZN => n2598);
   U2119 : OAI22_X1 port map( A1 => n30098, A2 => n36863, B1 => n30874, B2 => 
                           n36891, ZN => n36844);
   U2120 : INV_X1 port map( A => n36844, ZN => n2702);
   U2121 : OAI22_X1 port map( A1 => n30095, A2 => n36875, B1 => n30692, B2 => 
                           n36807, ZN => n36845);
   U2122 : INV_X1 port map( A => n36845, ZN => n2748);
   U2123 : OAI22_X1 port map( A1 => n30094, A2 => n36875, B1 => n30691, B2 => 
                           n36855, ZN => n36846);
   U2124 : INV_X1 port map( A => n36846, ZN => n2747);
   U2125 : OAI22_X1 port map( A1 => n30100, A2 => n36870, B1 => n30888, B2 => 
                           n36805, ZN => n36847);
   U2126 : INV_X1 port map( A => n36847, ZN => n2764);
   U2127 : OAI22_X1 port map( A1 => n30102, A2 => n36884, B1 => n30790, B2 => 
                           n36835, ZN => n36848);
   U2128 : INV_X1 port map( A => n36848, ZN => n2560);
   U2129 : OAI22_X1 port map( A1 => n30104, A2 => n36884, B1 => n30792, B2 => 
                           n36811, ZN => n36849);
   U2130 : INV_X1 port map( A => n36849, ZN => n2562);
   U2131 : OAI22_X1 port map( A1 => n30091, A2 => n36875, B1 => n30689, B2 => 
                           n36803, ZN => n36850);
   U2132 : INV_X1 port map( A => n36850, ZN => n2745);
   U2133 : OAI22_X1 port map( A1 => n30115, A2 => n36851, B1 => n30257, B2 => 
                           n36799, ZN => n36852);
   U2134 : INV_X1 port map( A => n36852, ZN => n2616);
   U2135 : OAI22_X1 port map( A1 => n30094, A2 => n36889, B1 => n30868, B2 => 
                           n36855, ZN => n36853);
   U2136 : INV_X1 port map( A => n36853, ZN => n2787);
   U2137 : OAI22_X1 port map( A1 => n30092, A2 => n36884, B1 => n30796, B2 => 
                           n36801, ZN => n36854);
   U2138 : INV_X1 port map( A => n36854, ZN => n2564);
   U2139 : OAI22_X1 port map( A1 => n30094, A2 => n36882, B1 => n30798, B2 => 
                           n36855, ZN => n36856);
   U2140 : INV_X1 port map( A => n36856, ZN => n2535);
   U2141 : OAI22_X1 port map( A1 => n30100, A2 => n36857, B1 => n30719, B2 => 
                           n36805, ZN => n36858);
   U2142 : INV_X1 port map( A => n36858, ZN => n2698);
   U2143 : OAI22_X1 port map( A1 => n30095, A2 => n36882, B1 => n30799, B2 => 
                           n36807, ZN => n36859);
   U2144 : INV_X1 port map( A => n36859, ZN => n2536);
   U2145 : OAI22_X1 port map( A1 => n30102, A2 => n36875, B1 => n30894, B2 => 
                           n36835, ZN => n36860);
   U2146 : INV_X1 port map( A => n36860, ZN => n2755);
   U2147 : OAI22_X1 port map( A1 => n30092, A2 => n36872, B1 => n30984, B2 => 
                           n36801, ZN => n36861);
   U2148 : INV_X1 port map( A => n36861, ZN => n2693);
   U2149 : OAI22_X1 port map( A1 => n30102, A2 => n36870, B1 => n30885, B2 => 
                           n36835, ZN => n36862);
   U2150 : INV_X1 port map( A => n36862, ZN => n2762);
   U2151 : OAI22_X1 port map( A1 => n30115, A2 => n36863, B1 => n30276, B2 => 
                           n36799, ZN => n36864);
   U2152 : INV_X1 port map( A => n36864, ZN => n2714);
   U2153 : OAI22_X1 port map( A1 => n30092, A2 => n36880, B1 => n30966, B2 => 
                           n36801, ZN => n36865);
   U2154 : INV_X1 port map( A => n36865, ZN => n2597);
   U2155 : OAI22_X1 port map( A1 => n30115, A2 => n36866, B1 => n30969, B2 => 
                           n36799, ZN => n36867);
   U2156 : INV_X1 port map( A => n36867, ZN => n2568);
   U2157 : OAI22_X1 port map( A1 => n30104, A2 => n36870, B1 => n30876, B2 => 
                           n36811, ZN => n36868);
   U2158 : INV_X1 port map( A => n36868, ZN => n2760);
   U2159 : OAI22_X1 port map( A1 => n30115, A2 => n36878, B1 => n30975, B2 => 
                           n36799, ZN => n36869);
   U2160 : INV_X1 port map( A => n36869, ZN => n2630);
   U2161 : OAI22_X1 port map( A1 => n30091, A2 => n36870, B1 => n30871, B2 => 
                           n36803, ZN => n36871);
   U2162 : INV_X1 port map( A => n36871, ZN => n2759);
   U2163 : OAI22_X1 port map( A1 => n30098, A2 => n36872, B1 => n30873, B2 => 
                           n36891, ZN => n36873);
   U2164 : INV_X1 port map( A => n36873, ZN => n2691);
   U2165 : OAI22_X1 port map( A1 => n30098, A2 => n36875, B1 => n30875, B2 => 
                           n36891, ZN => n36874);
   U2166 : INV_X1 port map( A => n36874, ZN => n2754);
   U2167 : OAI22_X1 port map( A1 => n30100, A2 => n36875, B1 => n30820, B2 => 
                           n36805, ZN => n36876);
   U2168 : INV_X1 port map( A => n36876, ZN => n2751);
   U2169 : OAI22_X1 port map( A1 => n30092, A2 => n36896, B1 => n31002, B2 => 
                           n36801, ZN => n36877);
   U2170 : INV_X1 port map( A => n36877, ZN => n2732);
   U2171 : OAI22_X1 port map( A1 => n30092, A2 => n36878, B1 => n30989, B2 => 
                           n36801, ZN => n36879);
   U2172 : INV_X1 port map( A => n36879, ZN => n2637);
   U2173 : OAI22_X1 port map( A1 => n30098, A2 => n36880, B1 => n30864, B2 => 
                           n36891, ZN => n36881);
   U2174 : INV_X1 port map( A => n36881, ZN => n2595);
   U2175 : OAI22_X1 port map( A1 => n30100, A2 => n36882, B1 => n30803, B2 => 
                           n36805, ZN => n36883);
   U2176 : INV_X1 port map( A => n36883, ZN => n2540);
   U2177 : OAI22_X1 port map( A1 => n30098, A2 => n36884, B1 => n30863, B2 => 
                           n36891, ZN => n36885);
   U2178 : INV_X1 port map( A => n36885, ZN => n2542);
   U2179 : OAI22_X1 port map( A1 => n30095, A2 => n36889, B1 => n30867, B2 => 
                           n36807, ZN => n36886);
   U2180 : INV_X1 port map( A => n36886, ZN => n2786);
   U2181 : OAI22_X1 port map( A1 => n30098, A2 => n36887, B1 => n30872, B2 => 
                           n36891, ZN => n36888);
   U2182 : INV_X1 port map( A => n36888, ZN => n2659);
   U2183 : OAI22_X1 port map( A1 => n30092, A2 => n36889, B1 => n30870, B2 => 
                           n36801, ZN => n36890);
   U2184 : INV_X1 port map( A => n36890, ZN => n2789);
   U2185 : OAI22_X1 port map( A1 => n30098, A2 => n36892, B1 => n30865, B2 => 
                           n36891, ZN => n36893);
   U2186 : INV_X1 port map( A => n36893, ZN => n2599);
   U2187 : OAI22_X1 port map( A1 => n30115, A2 => n36894, B1 => n30994, B2 => 
                           n36799, ZN => n36895);
   U2188 : INV_X1 port map( A => n36895, ZN => n2666);
   U2189 : OAI22_X1 port map( A1 => n30115, A2 => n36896, B1 => n30998, B2 => 
                           n36799, ZN => n36897);
   U2190 : INV_X1 port map( A => n36897, ZN => n2729);
   U2191 : INV_X1 port map( A => ADD_WR(3), ZN => n3559);
   U2192 : INV_X1 port map( A => ADD_WR(4), ZN => n3558);
   U2193 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1),
                           ZN => n18284);
   U2194 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n31231, ZN => 
                           n36904);
   U2195 : NOR2_X1 port map( A1 => n30129, A2 => n36904, ZN => n36902);
   U2196 : NAND2_X1 port map( A1 => n30048, A2 => n36902, ZN => n18360);
   U2197 : INV_X1 port map( A => ADD_WR(0), ZN => n36898);
   U2198 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n36898, ZN
                           => n18283);
   U2199 : NAND2_X1 port map( A1 => n36902, A2 => n30046, ZN => n18359);
   U2200 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n36898, ZN => n36899);
   U2201 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n36899, ZN => n18358);
   U2202 : NAND2_X1 port map( A1 => n36902, A2 => n30121, ZN => n18357);
   U2203 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n36900);
   U2204 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n36900, ZN => n18356);
   U2205 : NAND2_X1 port map( A1 => n36902, A2 => n30118, ZN => n18355);
   U2206 : INV_X1 port map( A => ADD_WR(2), ZN => n36901);
   U2207 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n36901, ZN
                           => n18282);
   U2208 : NAND2_X1 port map( A1 => n36902, A2 => n30044, ZN => n18354);
   U2209 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n36898, A3 => n36901, ZN =>
                           n18281);
   U2210 : NAND2_X1 port map( A1 => n36902, A2 => n30042, ZN => n18353);
   U2211 : NOR2_X1 port map( A1 => n36901, A2 => n36899, ZN => n18352);
   U2212 : NAND2_X1 port map( A1 => n36902, A2 => n30113, ZN => n18351);
   U2213 : NOR2_X1 port map( A1 => n36901, A2 => n36900, ZN => n18350);
   U2214 : NAND2_X1 port map( A1 => n36902, A2 => n30110, ZN => n18349);
   U2215 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n30130, ZN => 
                           n36906);
   U2216 : NOR2_X1 port map( A1 => n30129, A2 => n36906, ZN => n36903);
   U2217 : NAND2_X1 port map( A1 => n30048, A2 => n36903, ZN => n18348);
   U2218 : NAND2_X1 port map( A1 => n30046, A2 => n36903, ZN => n18347);
   U2219 : NAND2_X1 port map( A1 => n30121, A2 => n36903, ZN => n18346);
   U2220 : NAND2_X1 port map( A1 => n30118, A2 => n36903, ZN => n18345);
   U2221 : NAND2_X1 port map( A1 => n30044, A2 => n36903, ZN => n18344);
   U2222 : NAND2_X1 port map( A1 => n30042, A2 => n36903, ZN => n18343);
   U2223 : NAND2_X1 port map( A1 => n30113, A2 => n36903, ZN => n18342);
   U2224 : NAND2_X1 port map( A1 => n30110, A2 => n36903, ZN => n18341);
   U2225 : NOR2_X1 port map( A1 => n31229, A2 => n36904, ZN => n36905);
   U2226 : NAND2_X1 port map( A1 => n30048, A2 => n36905, ZN => n18340);
   U2227 : NAND2_X1 port map( A1 => n30046, A2 => n36905, ZN => n18339);
   U2228 : NAND2_X1 port map( A1 => n30121, A2 => n36905, ZN => n18338);
   U2229 : NAND2_X1 port map( A1 => n30118, A2 => n36905, ZN => n18337);
   U2230 : NAND2_X1 port map( A1 => n30044, A2 => n36905, ZN => n18336);
   U2231 : NAND2_X1 port map( A1 => n30042, A2 => n36905, ZN => n18335);
   U2232 : NAND2_X1 port map( A1 => n30113, A2 => n36905, ZN => n18334);
   U2233 : NAND2_X1 port map( A1 => n30110, A2 => n36905, ZN => n18333);
   U2234 : NOR2_X1 port map( A1 => n31229, A2 => n36906, ZN => n36907);
   U2235 : NAND2_X1 port map( A1 => n30048, A2 => n36907, ZN => n18332);
   U2236 : NAND2_X1 port map( A1 => n30046, A2 => n36907, ZN => n18331);
   U2237 : NAND2_X1 port map( A1 => n30121, A2 => n36907, ZN => n18330);
   U2238 : NAND2_X1 port map( A1 => n30118, A2 => n36907, ZN => n18329);
   U2239 : NAND2_X1 port map( A1 => n30044, A2 => n36907, ZN => n18328);
   U2240 : NAND2_X1 port map( A1 => n30042, A2 => n36907, ZN => n18327);
   U2241 : NAND2_X1 port map( A1 => n30113, A2 => n36907, ZN => n18326);
   U2242 : NAND2_X1 port map( A1 => n30110, A2 => n36907, ZN => n18325);
   U2243 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n3569, ZN => n36916);
   U2244 : INV_X1 port map( A => n3573, ZN => n36909);
   U2245 : NOR2_X1 port map( A1 => n36916, A2 => n36909, ZN => n18324);
   U2246 : INV_X1 port map( A => n3574, ZN => n36914);
   U2247 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n36911)
                           ;
   U2248 : NOR2_X1 port map( A1 => n36914, A2 => n36911, ZN => n18323);
   U2249 : NOR2_X1 port map( A1 => n36911, A2 => n3572, ZN => n18322);
   U2250 : INV_X1 port map( A => n3575, ZN => n36908);
   U2251 : NOR2_X1 port map( A1 => n36911, A2 => n36908, ZN => n18321);
   U2252 : NOR2_X1 port map( A1 => n36916, A2 => n3572, ZN => n18320);
   U2253 : INV_X1 port map( A => n3576, ZN => n36913);
   U2254 : NOR2_X1 port map( A1 => n36911, A2 => n36913, ZN => n18319);
   U2255 : INV_X1 port map( A => n3571, ZN => n36915);
   U2256 : NOR2_X1 port map( A1 => n36911, A2 => n36915, ZN => n18318);
   U2257 : NOR2_X1 port map( A1 => n36916, A2 => n36908, ZN => n18317);
   U2258 : INV_X1 port map( A => n3570, ZN => n36910);
   U2259 : NOR2_X1 port map( A1 => n36916, A2 => n36910, ZN => n18316);
   U2260 : NOR2_X1 port map( A1 => n36909, A2 => n36911, ZN => n18315);
   U2261 : NOR2_X1 port map( A1 => n36911, A2 => n36910, ZN => n18314);
   U2262 : INV_X1 port map( A => n3577, ZN => n36912);
   U2263 : NOR2_X1 port map( A1 => n36911, A2 => n36912, ZN => n18313);
   U2264 : NOR2_X1 port map( A1 => n36916, A2 => n36912, ZN => n18312);
   U2265 : NOR2_X1 port map( A1 => n36916, A2 => n36913, ZN => n18311);
   U2266 : NOR2_X1 port map( A1 => n36916, A2 => n36914, ZN => n18310);
   U2267 : NOR2_X1 port map( A1 => n36916, A2 => n36915, ZN => n18309);
   U2268 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n31273, A3 => n31270, ZN 
                           => n37627);
   U2269 : AOI22_X1 port map( A1 => n29373, A2 => n30072, B1 => n29374, B2 => 
                           n31223, ZN => n36920);
   U2270 : AOI22_X1 port map( A1 => n29895, A2 => n30079, B1 => n29900, B2 => 
                           n31222, ZN => n36919);
   U2271 : AOI22_X1 port map( A1 => n29914, A2 => n30083, B1 => n29377, B2 => 
                           n30078, ZN => n36918);
   U2272 : AOI22_X1 port map( A1 => n29872, A2 => n30082, B1 => n29880, B2 => 
                           n31224, ZN => n36917);
   U2273 : NAND4_X1 port map( A1 => n36920, A2 => n36919, A3 => n36918, A4 => 
                           n36917, ZN => n36926);
   U2274 : AOI22_X1 port map( A1 => n29375, A2 => n31227, B1 => n29309, B2 => 
                           n31226, ZN => n36924);
   U2275 : AOI22_X1 port map( A1 => n29369, A2 => n31225, B1 => n29376, B2 => 
                           n31228, ZN => n36923);
   U2276 : AOI22_X1 port map( A1 => n29891, A2 => n30073, B1 => n29371, B2 => 
                           n30071, ZN => n36922);
   U2277 : AOI22_X1 port map( A1 => n29370, A2 => n30069, B1 => n29372, B2 => 
                           n30084, ZN => n36921);
   U2278 : NAND4_X1 port map( A1 => n36924, A2 => n36923, A3 => n36922, A4 => 
                           n36921, ZN => n36925);
   U2279 : NOR2_X1 port map( A1 => n36926, A2 => n36925, ZN => n36938);
   U2280 : NOR3_X1 port map( A1 => n31266, A2 => n31267, A3 => n37448, ZN => 
                           n37378);
   U2281 : CLKBUF_X1 port map( A => n37378, Z => n37423);
   U2282 : AOI22_X1 port map( A1 => n30028, A2 => n31219, B1 => n30034, B2 => 
                           n31168, ZN => n36930);
   U2283 : AOI22_X1 port map( A1 => n30033, A2 => n31218, B1 => n30031, B2 => 
                           n31155, ZN => n36929);
   U2284 : AOI22_X1 port map( A1 => n30032, A2 => n31220, B1 => n30041, B2 => 
                           n31158, ZN => n36928);
   U2285 : AOI22_X1 port map( A1 => n30040, A2 => n31221, B1 => n30039, B2 => 
                           n31156, ZN => n36927);
   U2286 : NAND4_X1 port map( A1 => n36930, A2 => n36929, A3 => n36928, A4 => 
                           n36927, ZN => n36936);
   U2287 : NOR3_X1 port map( A1 => n31267, A2 => n30132, A3 => n37448, ZN => 
                           n37156);
   U2288 : CLKBUF_X1 port map( A => n37156, Z => n37622);
   U2289 : AOI22_X1 port map( A1 => n29713, A2 => n31233, B1 => n29675, B2 => 
                           n30050, ZN => n36934);
   U2290 : AOI22_X1 port map( A1 => n31158, A2 => n29381, B1 => n29382, B2 => 
                           n31214, ZN => n36933);
   U2291 : AOI22_X1 port map( A1 => n29380, A2 => n31162, B1 => n29694, B2 => 
                           n31157, ZN => n36932);
   U2292 : AOI22_X1 port map( A1 => n29579, A2 => n31216, B1 => n29364, B2 => 
                           n31215, ZN => n36931);
   U2293 : NAND4_X1 port map( A1 => n36934, A2 => n36933, A3 => n36932, A4 => 
                           n36931, ZN => n36935);
   U2294 : AOI22_X1 port map( A1 => n37423, A2 => n36936, B1 => n37622, B2 => 
                           n36935, ZN => n36937);
   U2295 : OAI21_X1 port map( B1 => n37448, B2 => n36938, A => n36937, ZN => 
                           OUT2(31));
   U2296 : AOI22_X1 port map( A1 => n30078, A2 => n29419, B1 => n29611, B2 => 
                           n30075, ZN => n36942);
   U2297 : AOI22_X1 port map( A1 => n31227, A2 => n29426, B1 => n30083, B2 => 
                           n29604, ZN => n36941);
   U2298 : AOI22_X1 port map( A1 => n31224, A2 => n29599, B1 => n29418, B2 => 
                           n30076, ZN => n36940);
   U2299 : AOI22_X1 port map( A1 => n30069, A2 => n29421, B1 => n29194, B2 => 
                           n31211, ZN => n36939);
   U2300 : NAND4_X1 port map( A1 => n36942, A2 => n36941, A3 => n36940, A4 => 
                           n36939, ZN => n36948);
   U2301 : AOI22_X1 port map( A1 => n30071, A2 => n29422, B1 => n29640, B2 => 
                           n31213, ZN => n36946);
   U2302 : AOI22_X1 port map( A1 => n31226, A2 => n29308, B1 => n30082, B2 => 
                           n29209, ZN => n36945);
   U2303 : AOI22_X1 port map( A1 => n30079, A2 => n29627, B1 => n29424, B2 => 
                           n30070, ZN => n36944);
   U2304 : AOI22_X1 port map( A1 => n29423, A2 => n31212, B1 => n29206, B2 => 
                           n30074, ZN => n36943);
   U2305 : NAND4_X1 port map( A1 => n36946, A2 => n36945, A3 => n36944, A4 => 
                           n36943, ZN => n36947);
   U2306 : NOR2_X1 port map( A1 => n36948, A2 => n36947, ZN => n36960);
   U2307 : AOI22_X1 port map( A1 => n31162, A2 => n29204, B1 => n31216, B2 => 
                           n29205, ZN => n36952);
   U2308 : AOI22_X1 port map( A1 => n29202, A2 => n31161, B1 => n29615, B2 => 
                           n31210, ZN => n36951);
   U2309 : AOI22_X1 port map( A1 => n31219, A2 => n29636, B1 => n30050, B2 => 
                           n29179, ZN => n36950);
   U2310 : AOI22_X1 port map( A1 => n31158, A2 => n29203, B1 => n31156, B2 => 
                           n29199, ZN => n36949);
   U2311 : NAND4_X1 port map( A1 => n36952, A2 => n36951, A3 => n36950, A4 => 
                           n36949, ZN => n36958);
   U2312 : AOI22_X1 port map( A1 => n31162, A2 => n29427, B1 => n29648, B2 => 
                           n31209, ZN => n36956);
   U2313 : AOI22_X1 port map( A1 => n31233, A2 => n29662, B1 => n29189, B2 => 
                           n31208, ZN => n36955);
   U2314 : AOI22_X1 port map( A1 => n31161, A2 => n29393, B1 => n31210, B2 => 
                           n29655, ZN => n36954);
   U2315 : AOI22_X1 port map( A1 => n31156, A2 => n29365, B1 => n31216, B2 => 
                           n29598, ZN => n36953);
   U2316 : NAND4_X1 port map( A1 => n36956, A2 => n36955, A3 => n36954, A4 => 
                           n36953, ZN => n36957);
   U2317 : AOI22_X1 port map( A1 => n37423, A2 => n36958, B1 => n37622, B2 => 
                           n36957, ZN => n36959);
   U2318 : OAI21_X1 port map( B1 => n37448, B2 => n36960, A => n36959, ZN => 
                           OUT2(30));
   U2319 : AOI22_X1 port map( A1 => n30076, A2 => n29407, B1 => n29957, B2 => 
                           n31205, ZN => n36964);
   U2320 : AOI22_X1 port map( A1 => n30071, A2 => n29410, B1 => n30079, B2 => 
                           n30022, ZN => n36963);
   U2321 : AOI22_X1 port map( A1 => n30072, A2 => n29412, B1 => n30078, B2 => 
                           n29401, ZN => n36962);
   U2322 : AOI22_X1 port map( A1 => n31223, A2 => n29413, B1 => n31224, B2 => 
                           n30010, ZN => n36961);
   U2323 : NAND4_X1 port map( A1 => n36964, A2 => n36963, A3 => n36962, A4 => 
                           n36961, ZN => n36970);
   U2324 : AOI22_X1 port map( A1 => n31228, A2 => n29400, B1 => n29307, B2 => 
                           n30080, ZN => n36968);
   U2325 : AOI22_X1 port map( A1 => n30084, A2 => n29411, B1 => n31222, B2 => 
                           n29984, ZN => n36967);
   U2326 : AOI22_X1 port map( A1 => n30073, A2 => n29944, B1 => n29409, B2 => 
                           n31206, ZN => n36966);
   U2327 : AOI22_X1 port map( A1 => n29889, A2 => n31207, B1 => n29414, B2 => 
                           n30077, ZN => n36965);
   U2328 : NAND4_X1 port map( A1 => n36968, A2 => n36967, A3 => n36966, A4 => 
                           n36965, ZN => n36969);
   U2329 : NOR2_X1 port map( A1 => n36970, A2 => n36969, ZN => n36982);
   U2330 : AOI22_X1 port map( A1 => n31216, A2 => n29912, B1 => n30035, B2 => 
                           n31165, ZN => n36974);
   U2331 : AOI22_X1 port map( A1 => n30050, A2 => n29911, B1 => n29913, B2 => 
                           n31204, ZN => n36973);
   U2332 : AOI22_X1 port map( A1 => n31218, A2 => n30036, B1 => n31208, B2 => 
                           n29915, ZN => n36972);
   U2333 : AOI22_X1 port map( A1 => n31220, A2 => n29916, B1 => n31156, B2 => 
                           n29917, ZN => n36971);
   U2334 : NAND4_X1 port map( A1 => n36974, A2 => n36973, A3 => n36972, A4 => 
                           n36971, ZN => n36980);
   U2335 : AOI22_X1 port map( A1 => n31168, A2 => n29706, B1 => n31233, B2 => 
                           n29707, ZN => n36978);
   U2336 : AOI22_X1 port map( A1 => n31218, A2 => n29696, B1 => n31220, B2 => 
                           n29392, ZN => n36977);
   U2337 : AOI22_X1 port map( A1 => n31156, A2 => n29366, B1 => n31208, B2 => 
                           n29406, ZN => n36976);
   U2338 : AOI22_X1 port map( A1 => n31155, A2 => n29595, B1 => n31162, B2 => 
                           n29281, ZN => n36975);
   U2339 : NAND4_X1 port map( A1 => n36978, A2 => n36977, A3 => n36976, A4 => 
                           n36975, ZN => n36979);
   U2340 : AOI22_X1 port map( A1 => n37423, A2 => n36980, B1 => n37622, B2 => 
                           n36979, ZN => n36981);
   U2341 : OAI21_X1 port map( B1 => n37448, B2 => n36982, A => n36981, ZN => 
                           OUT2(29));
   U2342 : AOI22_X1 port map( A1 => n30082, A2 => n29184, B1 => n29608, B2 => 
                           n30081, ZN => n36986);
   U2343 : AOI22_X1 port map( A1 => n30078, A2 => n29439, B1 => n29626, B2 => 
                           n31203, ZN => n36985);
   U2344 : AOI22_X1 port map( A1 => n31228, A2 => n29183, B1 => n30072, B2 => 
                           n29449, ZN => n36984);
   U2345 : AOI22_X1 port map( A1 => n31222, A2 => n29618, B1 => n30076, B2 => 
                           n29420, ZN => n36983);
   U2346 : NAND4_X1 port map( A1 => n36986, A2 => n36985, A3 => n36984, A4 => 
                           n36983, ZN => n36992);
   U2347 : AOI22_X1 port map( A1 => n30071, A2 => n29444, B1 => n31213, B2 => 
                           n29639, ZN => n36990);
   U2348 : AOI22_X1 port map( A1 => n31223, A2 => n29450, B1 => n31211, B2 => 
                           n29186, ZN => n36989);
   U2349 : AOI22_X1 port map( A1 => n30069, A2 => n29443, B1 => n30080, B2 => 
                           n29300, ZN => n36988);
   U2350 : AOI22_X1 port map( A1 => n30083, A2 => n29619, B1 => n30077, B2 => 
                           n29437, ZN => n36987);
   U2351 : NAND4_X1 port map( A1 => n36990, A2 => n36989, A3 => n36988, A4 => 
                           n36987, ZN => n36991);
   U2352 : NOR2_X1 port map( A1 => n36992, A2 => n36991, ZN => n37004);
   U2353 : AOI22_X1 port map( A1 => n31158, A2 => n29197, B1 => n31221, B2 => 
                           n29196, ZN => n36996);
   U2354 : AOI22_X1 port map( A1 => n31156, A2 => n29200, B1 => n31165, B2 => 
                           n29635, ZN => n36995);
   U2355 : AOI22_X1 port map( A1 => n31168, A2 => n29190, B1 => n31214, B2 => 
                           n29198, ZN => n36994);
   U2356 : AOI22_X1 port map( A1 => n31157, A2 => n29614, B1 => n29191, B2 => 
                           n31217, ZN => n36993);
   U2357 : NAND4_X1 port map( A1 => n36996, A2 => n36995, A3 => n36994, A4 => 
                           n36993, ZN => n37002);
   U2358 : AOI22_X1 port map( A1 => n31214, A2 => n29391, B1 => n31157, B2 => 
                           n29654, ZN => n37000);
   U2359 : AOI22_X1 port map( A1 => n31155, A2 => n29583, B1 => n31233, B2 => 
                           n29632, ZN => n36999);
   U2360 : AOI22_X1 port map( A1 => n31162, A2 => n29441, B1 => n29367, B2 => 
                           n31202, ZN => n36998);
   U2361 : AOI22_X1 port map( A1 => n30050, A2 => n29647, B1 => n29185, B2 => 
                           n31201, ZN => n36997);
   U2362 : NAND4_X1 port map( A1 => n37000, A2 => n36999, A3 => n36998, A4 => 
                           n36997, ZN => n37001);
   U2363 : AOI22_X1 port map( A1 => n37423, A2 => n37002, B1 => n37622, B2 => 
                           n37001, ZN => n37003);
   U2364 : OAI21_X1 port map( B1 => n37448, B2 => n37004, A => n37003, ZN => 
                           OUT2(28));
   U2365 : AOI22_X1 port map( A1 => n30083, A2 => n29623, B1 => n29435, B2 => 
                           n31200, ZN => n37008);
   U2366 : AOI22_X1 port map( A1 => n30084, A2 => n29193, B1 => n30080, B2 => 
                           n29299, ZN => n37007);
   U2367 : AOI22_X1 port map( A1 => n30072, A2 => n29436, B1 => n30077, B2 => 
                           n29430, ZN => n37006);
   U2368 : AOI22_X1 port map( A1 => n31203, A2 => n29625, B1 => n30081, B2 => 
                           n29617, ZN => n37005);
   U2369 : NAND4_X1 port map( A1 => n37008, A2 => n37007, A3 => n37006, A4 => 
                           n37005, ZN => n37014);
   U2370 : AOI22_X1 port map( A1 => n30073, A2 => n29638, B1 => n30078, B2 => 
                           n29431, ZN => n37012);
   U2371 : AOI22_X1 port map( A1 => n30069, A2 => n29434, B1 => n30070, B2 => 
                           n29429, ZN => n37011);
   U2372 : AOI22_X1 port map( A1 => n30082, A2 => n29187, B1 => n30075, B2 => 
                           n29606, ZN => n37010);
   U2373 : AOI22_X1 port map( A1 => n31228, A2 => n29188, B1 => n30076, B2 => 
                           n29433, ZN => n37009);
   U2374 : NAND4_X1 port map( A1 => n37012, A2 => n37011, A3 => n37010, A4 => 
                           n37009, ZN => n37013);
   U2375 : NOR2_X1 port map( A1 => n37014, A2 => n37013, ZN => n37026);
   U2376 : AOI22_X1 port map( A1 => n31210, A2 => n29631, B1 => n31201, B2 => 
                           n29178, ZN => n37018);
   U2377 : AOI22_X1 port map( A1 => n31219, A2 => n29634, B1 => n30050, B2 => 
                           n29175, ZN => n37017);
   U2378 : AOI22_X1 port map( A1 => n31162, A2 => n29177, B1 => n31161, B2 => 
                           n29180, ZN => n37016);
   U2379 : AOI22_X1 port map( A1 => n31216, A2 => n29167, B1 => n31202, B2 => 
                           n29182, ZN => n37015);
   U2380 : NAND4_X1 port map( A1 => n37018, A2 => n37017, A3 => n37016, A4 => 
                           n37015, ZN => n37024);
   U2381 : AOI22_X1 port map( A1 => n31209, A2 => n29646, B1 => n31201, B2 => 
                           n29181, ZN => n37022);
   U2382 : AOI22_X1 port map( A1 => n31233, A2 => n29661, B1 => n31215, B2 => 
                           n29368, ZN => n37021);
   U2383 : AOI22_X1 port map( A1 => n31214, A2 => n29390, B1 => n31217, B2 => 
                           n29597, ZN => n37020);
   U2384 : AOI22_X1 port map( A1 => n31162, A2 => n29432, B1 => n31157, B2 => 
                           n29653, ZN => n37019);
   U2385 : NAND4_X1 port map( A1 => n37022, A2 => n37021, A3 => n37020, A4 => 
                           n37019, ZN => n37023);
   U2386 : AOI22_X1 port map( A1 => n37423, A2 => n37024, B1 => n37156, B2 => 
                           n37023, ZN => n37025);
   U2387 : OAI21_X1 port map( B1 => n37448, B2 => n37026, A => n37025, ZN => 
                           OUT2(27));
   U2388 : AOI22_X1 port map( A1 => n30083, A2 => n29945, B1 => n30081, B2 => 
                           n30017, ZN => n37030);
   U2389 : AOI22_X1 port map( A1 => n31227, A2 => n29467, B1 => n30070, B2 => 
                           n29466, ZN => n37029);
   U2390 : AOI22_X1 port map( A1 => n30073, A2 => n29964, B1 => n30078, B2 => 
                           n29469, ZN => n37028);
   U2391 : AOI22_X1 port map( A1 => n31226, A2 => n29298, B1 => n30074, B2 => 
                           n29468, ZN => n37027);
   U2392 : NAND4_X1 port map( A1 => n37030, A2 => n37029, A3 => n37028, A4 => 
                           n37027, ZN => n37036);
   U2393 : AOI22_X1 port map( A1 => n30079, A2 => n30023, B1 => n30075, B2 => 
                           n29983, ZN => n37034);
   U2394 : AOI22_X1 port map( A1 => n30076, A2 => n29453, B1 => n31207, B2 => 
                           n29890, ZN => n37033);
   U2395 : AOI22_X1 port map( A1 => n31212, A2 => n29465, B1 => n31200, B2 => 
                           n29463, ZN => n37032);
   U2396 : AOI22_X1 port map( A1 => n30069, A2 => n29461, B1 => n30084, B2 => 
                           n29464, ZN => n37031);
   U2397 : NAND4_X1 port map( A1 => n37034, A2 => n37033, A3 => n37032, A4 => 
                           n37031, ZN => n37035);
   U2398 : NOR2_X1 port map( A1 => n37036, A2 => n37035, ZN => n37048);
   U2399 : AOI22_X1 port map( A1 => n31155, A2 => n29898, B1 => n31215, B2 => 
                           n29909, ZN => n37040);
   U2400 : AOI22_X1 port map( A1 => n31168, A2 => n29899, B1 => n31208, B2 => 
                           n29896, ZN => n37039);
   U2401 : AOI22_X1 port map( A1 => n31219, A2 => n30037, B1 => n31161, B2 => 
                           n29910, ZN => n37038);
   U2402 : AOI22_X1 port map( A1 => n31162, A2 => n29897, B1 => n31157, B2 => 
                           n30029, ZN => n37037);
   U2403 : NAND4_X1 port map( A1 => n37040, A2 => n37039, A3 => n37038, A4 => 
                           n37037, ZN => n37046);
   U2404 : AOI22_X1 port map( A1 => n31218, A2 => n29681, B1 => n30050, B2 => 
                           n29682, ZN => n37044);
   U2405 : AOI22_X1 port map( A1 => n31155, A2 => n29587, B1 => n31161, B2 => 
                           n29389, ZN => n37043);
   U2406 : AOI22_X1 port map( A1 => n31219, A2 => n29704, B1 => n31158, B2 => 
                           n29428, ZN => n37042);
   U2407 : AOI22_X1 port map( A1 => n31162, A2 => n29472, B1 => n31215, B2 => 
                           n29378, ZN => n37041);
   U2408 : NAND4_X1 port map( A1 => n37044, A2 => n37043, A3 => n37042, A4 => 
                           n37041, ZN => n37045);
   U2409 : AOI22_X1 port map( A1 => n37423, A2 => n37046, B1 => n37156, B2 => 
                           n37045, ZN => n37047);
   U2410 : OAI21_X1 port map( B1 => n37448, B2 => n37048, A => n37047, ZN => 
                           OUT2(26));
   U2411 : AOI22_X1 port map( A1 => n30074, A2 => n29170, B1 => n30070, B2 => 
                           n29481, ZN => n37052);
   U2412 : AOI22_X1 port map( A1 => n30084, A2 => n29169, B1 => n30072, B2 => 
                           n29480, ZN => n37051);
   U2413 : AOI22_X1 port map( A1 => n31207, A2 => n29171, B1 => n30077, B2 => 
                           n29482, ZN => n37050);
   U2414 : AOI22_X1 port map( A1 => n31225, A2 => n29352, B1 => n30078, B2 => 
                           n29483, ZN => n37049);
   U2415 : NAND4_X1 port map( A1 => n37052, A2 => n37051, A3 => n37050, A4 => 
                           n37049, ZN => n37058);
   U2416 : AOI22_X1 port map( A1 => n30075, A2 => n29605, B1 => n31205, B2 => 
                           n29622, ZN => n37056);
   U2417 : AOI22_X1 port map( A1 => n31213, A2 => n29637, B1 => n31206, B2 => 
                           n29353, ZN => n37055);
   U2418 : AOI22_X1 port map( A1 => n31224, A2 => n29600, B1 => n31200, B2 => 
                           n29351, ZN => n37054);
   U2419 : AOI22_X1 port map( A1 => n30079, A2 => n29624, B1 => n30080, B2 => 
                           n29297, ZN => n37053);
   U2420 : NAND4_X1 port map( A1 => n37056, A2 => n37055, A3 => n37054, A4 => 
                           n37053, ZN => n37057);
   U2421 : NOR2_X1 port map( A1 => n37058, A2 => n37057, ZN => n37070);
   U2422 : AOI22_X1 port map( A1 => n31161, A2 => n29168, B1 => n31204, B2 => 
                           n29176, ZN => n37062);
   U2423 : AOI22_X1 port map( A1 => n31233, A2 => n29633, B1 => n31215, B2 => 
                           n29173, ZN => n37061);
   U2424 : AOI22_X1 port map( A1 => n30050, A2 => n29223, B1 => n31210, B2 => 
                           n29612, ZN => n37060);
   U2425 : AOI22_X1 port map( A1 => n31216, A2 => n29213, B1 => n31201, B2 => 
                           n29174, ZN => n37059);
   U2426 : NAND4_X1 port map( A1 => n37062, A2 => n37061, A3 => n37060, A4 => 
                           n37059, ZN => n37068);
   U2427 : AOI22_X1 port map( A1 => n31218, A2 => n29652, B1 => n31202, B2 => 
                           n29330, ZN => n37066);
   U2428 : AOI22_X1 port map( A1 => n31233, A2 => n29659, B1 => n31161, B2 => 
                           n29278, ZN => n37065);
   U2429 : AOI22_X1 port map( A1 => n31221, A2 => n29425, B1 => n31209, B2 => 
                           n29645, ZN => n37064);
   U2430 : AOI22_X1 port map( A1 => n31155, A2 => n29594, B1 => n31201, B2 => 
                           n29192, ZN => n37063);
   U2431 : NAND4_X1 port map( A1 => n37066, A2 => n37065, A3 => n37064, A4 => 
                           n37063, ZN => n37067);
   U2432 : AOI22_X1 port map( A1 => n37423, A2 => n37068, B1 => n37156, B2 => 
                           n37067, ZN => n37069);
   U2433 : OAI21_X1 port map( B1 => n37448, B2 => n37070, A => n37069, ZN => 
                           OUT2(25));
   U2434 : AOI22_X1 port map( A1 => n30075, A2 => n29982, B1 => n31207, B2 => 
                           n29930, ZN => n37074);
   U2435 : AOI22_X1 port map( A1 => n31227, A2 => n29303, B1 => n30071, B2 => 
                           n29306, ZN => n37073);
   U2436 : AOI22_X1 port map( A1 => n31203, A2 => n30025, B1 => n29301, B2 => 
                           n31199, ZN => n37072);
   U2437 : AOI22_X1 port map( A1 => n31205, A2 => n29960, B1 => n30081, B2 => 
                           n30018, ZN => n37071);
   U2438 : NAND4_X1 port map( A1 => n37074, A2 => n37073, A3 => n37072, A4 => 
                           n37071, ZN => n37080);
   U2439 : AOI22_X1 port map( A1 => n30074, A2 => n29302, B1 => n30080, B2 => 
                           n29276, ZN => n37078);
   U2440 : AOI22_X1 port map( A1 => n31225, A2 => n29284, B1 => n30073, B2 => 
                           n29952, ZN => n37077);
   U2441 : AOI22_X1 port map( A1 => n31223, A2 => n29304, B1 => n31211, B2 => 
                           n29554, ZN => n37076);
   U2442 : AOI22_X1 port map( A1 => n30072, A2 => n29305, B1 => n31206, B2 => 
                           n29283, ZN => n37075);
   U2443 : NAND4_X1 port map( A1 => n37078, A2 => n37077, A3 => n37076, A4 => 
                           n37075, ZN => n37079);
   U2444 : NOR2_X1 port map( A1 => n37080, A2 => n37079, ZN => n37092);
   U2445 : AOI22_X1 port map( A1 => n31156, A2 => n29927, B1 => n31216, B2 => 
                           n29929, ZN => n37084);
   U2446 : AOI22_X1 port map( A1 => n31168, A2 => n29928, B1 => n31208, B2 => 
                           n29931, ZN => n37083);
   U2447 : AOI22_X1 port map( A1 => n31221, A2 => n29926, B1 => n31165, B2 => 
                           n30030, ZN => n37082);
   U2448 : AOI22_X1 port map( A1 => n31214, A2 => n29932, B1 => n31157, B2 => 
                           n30038, ZN => n37081);
   U2449 : NAND4_X1 port map( A1 => n37084, A2 => n37083, A3 => n37082, A4 => 
                           n37081, ZN => n37090);
   U2450 : AOI22_X1 port map( A1 => n31214, A2 => n29287, B1 => n31208, B2 => 
                           n29288, ZN => n37088);
   U2451 : AOI22_X1 port map( A1 => n31157, A2 => n29712, B1 => n31217, B2 => 
                           n29588, ZN => n37087);
   U2452 : AOI22_X1 port map( A1 => n31221, A2 => n29296, B1 => n31233, B2 => 
                           n29692, ZN => n37086);
   U2453 : AOI22_X1 port map( A1 => n31168, A2 => n29684, B1 => n31215, B2 => 
                           n29286, ZN => n37085);
   U2454 : NAND4_X1 port map( A1 => n37088, A2 => n37087, A3 => n37086, A4 => 
                           n37085, ZN => n37089);
   U2455 : AOI22_X1 port map( A1 => n37423, A2 => n37090, B1 => n37156, B2 => 
                           n37089, ZN => n37091);
   U2456 : OAI21_X1 port map( B1 => n37448, B2 => n37092, A => n37091, ZN => 
                           OUT2(24));
   U2457 : AOI22_X1 port map( A1 => n30075, A2 => n29610, B1 => n31203, B2 => 
                           n29660, ZN => n37096);
   U2458 : AOI22_X1 port map( A1 => n31200, A2 => n29567, B1 => n31199, B2 => 
                           n29555, ZN => n37095);
   U2459 : AOI22_X1 port map( A1 => n31223, A2 => n29514, B1 => n30081, B2 => 
                           n29609, ZN => n37094);
   U2460 : AOI22_X1 port map( A1 => n31213, A2 => n29607, B1 => n30074, B2 => 
                           n29548, ZN => n37093);
   U2461 : NAND4_X1 port map( A1 => n37096, A2 => n37095, A3 => n37094, A4 => 
                           n37093, ZN => n37102);
   U2462 : AOI22_X1 port map( A1 => n30072, A2 => n29569, B1 => n30083, B2 => 
                           n29621, ZN => n37100);
   U2463 : AOI22_X1 port map( A1 => n30069, A2 => n29344, B1 => n30082, B2 => 
                           n29649, ZN => n37099);
   U2464 : AOI22_X1 port map( A1 => n31211, A2 => n29568, B1 => n30077, B2 => 
                           n29536, ZN => n37098);
   U2465 : AOI22_X1 port map( A1 => n31225, A2 => n29457, B1 => n30080, B2 => 
                           n29275, ZN => n37097);
   U2466 : NAND4_X1 port map( A1 => n37100, A2 => n37099, A3 => n37098, A4 => 
                           n37097, ZN => n37101);
   U2467 : NOR2_X1 port map( A1 => n37102, A2 => n37101, ZN => n37114);
   U2468 : AOI22_X1 port map( A1 => n30050, A2 => n29207, B1 => n31216, B2 => 
                           n29195, ZN => n37106);
   U2469 : AOI22_X1 port map( A1 => n31221, A2 => n29225, B1 => n31165, B2 => 
                           n29212, ZN => n37105);
   U2470 : AOI22_X1 port map( A1 => n31156, A2 => n29231, B1 => n31201, B2 => 
                           n29226, ZN => n37104);
   U2471 : AOI22_X1 port map( A1 => n31214, A2 => n29228, B1 => n31210, B2 => 
                           n29208, ZN => n37103);
   U2472 : NAND4_X1 port map( A1 => n37106, A2 => n37105, A3 => n37104, A4 => 
                           n37103, ZN => n37112);
   U2473 : AOI22_X1 port map( A1 => n31155, A2 => n29581, B1 => n31201, B2 => 
                           n29230, ZN => n37110);
   U2474 : AOI22_X1 port map( A1 => n31221, A2 => n29462, B1 => n31157, B2 => 
                           n29651, ZN => n37109);
   U2475 : AOI22_X1 port map( A1 => n30050, A2 => n29644, B1 => n31215, B2 => 
                           n29379, ZN => n37108);
   U2476 : AOI22_X1 port map( A1 => n31219, A2 => n29657, B1 => n31161, B2 => 
                           n29221, ZN => n37107);
   U2477 : NAND4_X1 port map( A1 => n37110, A2 => n37109, A3 => n37108, A4 => 
                           n37107, ZN => n37111);
   U2478 : AOI22_X1 port map( A1 => n37423, A2 => n37112, B1 => n37156, B2 => 
                           n37111, ZN => n37113);
   U2479 : OAI21_X1 port map( B1 => n37627, B2 => n37114, A => n37113, ZN => 
                           OUT2(23));
   U2480 : AOI22_X1 port map( A1 => n31223, A2 => n29507, B1 => n30074, B2 => 
                           n29549, ZN => n37118);
   U2481 : AOI22_X1 port map( A1 => n30077, A2 => n29537, B1 => n31199, B2 => 
                           n29556, ZN => n37117);
   U2482 : AOI22_X1 port map( A1 => n30073, A2 => n29629, B1 => n30079, B2 => 
                           n29658, ZN => n37116);
   U2483 : AOI22_X1 port map( A1 => n31205, A2 => n29620, B1 => n30081, B2 => 
                           n29613, ZN => n37115);
   U2484 : NAND4_X1 port map( A1 => n37118, A2 => n37117, A3 => n37116, A4 => 
                           n37115, ZN => n37124);
   U2485 : AOI22_X1 port map( A1 => n31211, A2 => n29566, B1 => n31207, B2 => 
                           n29630, ZN => n37122);
   U2486 : AOI22_X1 port map( A1 => n31226, A2 => n29274, B1 => n30069, B2 => 
                           n29343, ZN => n37121);
   U2487 : AOI22_X1 port map( A1 => n30071, A2 => n29565, B1 => n31222, B2 => 
                           n29642, ZN => n37120);
   U2488 : AOI22_X1 port map( A1 => n31212, A2 => n29564, B1 => n30076, B2 => 
                           n29458, ZN => n37119);
   U2489 : NAND4_X1 port map( A1 => n37122, A2 => n37121, A3 => n37120, A4 => 
                           n37119, ZN => n37123);
   U2490 : NOR2_X1 port map( A1 => n37124, A2 => n37123, ZN => n37136);
   U2491 : AOI22_X1 port map( A1 => n31221, A2 => n29222, B1 => n31157, B2 => 
                           n29218, ZN => n37128);
   U2492 : AOI22_X1 port map( A1 => n31233, A2 => n29217, B1 => n31201, B2 => 
                           n29224, ZN => n37127);
   U2493 : AOI22_X1 port map( A1 => n30050, A2 => n29219, B1 => n31217, B2 => 
                           n29220, ZN => n37126);
   U2494 : AOI22_X1 port map( A1 => n31156, A2 => n29229, B1 => n31214, B2 => 
                           n29227, ZN => n37125);
   U2495 : NAND4_X1 port map( A1 => n37128, A2 => n37127, A3 => n37126, A4 => 
                           n37125, ZN => n37134);
   U2496 : AOI22_X1 port map( A1 => n31208, A2 => n29214, B1 => n31217, B2 => 
                           n29589, ZN => n37132);
   U2497 : AOI22_X1 port map( A1 => n31221, A2 => n29456, B1 => n31209, B2 => 
                           n29643, ZN => n37131);
   U2498 : AOI22_X1 port map( A1 => n31156, A2 => n29383, B1 => n31214, B2 => 
                           n29216, ZN => n37130);
   U2499 : AOI22_X1 port map( A1 => n31233, A2 => n29656, B1 => n31157, B2 => 
                           n29650, ZN => n37129);
   U2500 : NAND4_X1 port map( A1 => n37132, A2 => n37131, A3 => n37130, A4 => 
                           n37129, ZN => n37133);
   U2501 : AOI22_X1 port map( A1 => n37423, A2 => n37134, B1 => n37156, B2 => 
                           n37133, ZN => n37135);
   U2502 : OAI21_X1 port map( B1 => n37627, B2 => n37136, A => n37135, ZN => 
                           OUT2(22));
   U2503 : AOI22_X1 port map( A1 => n30079, A2 => n29988, B1 => n31212, B2 => 
                           n29349, ZN => n37140);
   U2504 : AOI22_X1 port map( A1 => n31226, A2 => n29273, B1 => n30083, B2 => 
                           n29966, ZN => n37139);
   U2505 : AOI22_X1 port map( A1 => n31206, A2 => n29335, B1 => n30081, B2 => 
                           n30019, ZN => n37138);
   U2506 : AOI22_X1 port map( A1 => n30073, A2 => n29946, B1 => n30078, B2 => 
                           n29345, ZN => n37137);
   U2507 : NAND4_X1 port map( A1 => n37140, A2 => n37139, A3 => n37138, A4 => 
                           n37137, ZN => n37146);
   U2508 : AOI22_X1 port map( A1 => n30071, A2 => n29334, B1 => n30070, B2 => 
                           n29348, ZN => n37144);
   U2509 : AOI22_X1 port map( A1 => n30076, A2 => n29336, B1 => n30077, B2 => 
                           n29347, ZN => n37143);
   U2510 : AOI22_X1 port map( A1 => n30084, A2 => n29350, B1 => n30075, B2 => 
                           n29981, ZN => n37142);
   U2511 : AOI22_X1 port map( A1 => n30074, A2 => n29346, B1 => n31207, B2 => 
                           n29999, ZN => n37141);
   U2512 : NAND4_X1 port map( A1 => n37144, A2 => n37143, A3 => n37142, A4 => 
                           n37141, ZN => n37145);
   U2513 : NOR2_X1 port map( A1 => n37146, A2 => n37145, ZN => n37159);
   U2514 : AOI22_X1 port map( A1 => n31155, A2 => n29850, B1 => n31221, B2 => 
                           n29849, ZN => n37150);
   U2515 : AOI22_X1 port map( A1 => n31168, A2 => n29852, B1 => n31165, B2 => 
                           n29855, ZN => n37149);
   U2516 : AOI22_X1 port map( A1 => n31210, A2 => n29853, B1 => n31201, B2 => 
                           n29848, ZN => n37148);
   U2517 : AOI22_X1 port map( A1 => n31214, A2 => n29847, B1 => n31202, B2 => 
                           n29846, ZN => n37147);
   U2518 : NAND4_X1 port map( A1 => n37150, A2 => n37149, A3 => n37148, A4 => 
                           n37147, ZN => n37157);
   U2519 : AOI22_X1 port map( A1 => n31158, A2 => n29339, B1 => n31156, B2 => 
                           n29337, ZN => n37154);
   U2520 : AOI22_X1 port map( A1 => n31220, A2 => n29338, B1 => n31221, B2 => 
                           n29340, ZN => n37153);
   U2521 : AOI22_X1 port map( A1 => n31157, A2 => n29671, B1 => n31217, B2 => 
                           n29591, ZN => n37152);
   U2522 : AOI22_X1 port map( A1 => n31233, A2 => n29698, B1 => n30050, B2 => 
                           n29687, ZN => n37151);
   U2523 : NAND4_X1 port map( A1 => n37154, A2 => n37153, A3 => n37152, A4 => 
                           n37151, ZN => n37155);
   U2524 : AOI22_X1 port map( A1 => n37423, A2 => n37157, B1 => n37156, B2 => 
                           n37155, ZN => n37158);
   U2525 : OAI21_X1 port map( B1 => n37627, B2 => n37159, A => n37158, ZN => 
                           OUT2(21));
   U2526 : AOI22_X1 port map( A1 => n30073, A2 => n29601, B1 => n30070, B2 => 
                           n29506, ZN => n37163);
   U2527 : AOI22_X1 port map( A1 => n30080, A2 => n29272, B1 => n31205, B2 => 
                           n29602, ZN => n37162);
   U2528 : AOI22_X1 port map( A1 => n30071, A2 => n29570, B1 => n30077, B2 => 
                           n29538, ZN => n37161);
   U2529 : AOI22_X1 port map( A1 => n31228, A2 => n29550, B1 => n30082, B2 => 
                           n29628, ZN => n37160);
   U2530 : NAND4_X1 port map( A1 => n37163, A2 => n37162, A3 => n37161, A4 => 
                           n37160, ZN => n37169);
   U2531 : AOI22_X1 port map( A1 => n30079, A2 => n29616, B1 => n30072, B2 => 
                           n29576, ZN => n37167);
   U2532 : AOI22_X1 port map( A1 => n30078, A2 => n29557, B1 => n30076, B2 => 
                           n29459, ZN => n37166);
   U2533 : AOI22_X1 port map( A1 => n30069, A2 => n29342, B1 => n30075, B2 => 
                           n29641, ZN => n37165);
   U2534 : AOI22_X1 port map( A1 => n30084, A2 => n29575, B1 => n31224, B2 => 
                           n29603, ZN => n37164);
   U2535 : NAND4_X1 port map( A1 => n37167, A2 => n37166, A3 => n37165, A4 => 
                           n37164, ZN => n37168);
   U2536 : NOR2_X1 port map( A1 => n37169, A2 => n37168, ZN => n37181);
   U2537 : AOI22_X1 port map( A1 => n31210, A2 => n29240, B1 => n31208, B2 => 
                           n29238, ZN => n37173);
   U2538 : AOI22_X1 port map( A1 => n31219, A2 => n29234, B1 => n30050, B2 => 
                           n29232, ZN => n37172);
   U2539 : AOI22_X1 port map( A1 => n31155, A2 => n29235, B1 => n31221, B2 => 
                           n29243, ZN => n37171);
   U2540 : AOI22_X1 port map( A1 => n31156, A2 => n29241, B1 => n31161, B2 => 
                           n29242, ZN => n37170);
   U2541 : NAND4_X1 port map( A1 => n37173, A2 => n37172, A3 => n37171, A4 => 
                           n37170, ZN => n37179);
   U2542 : AOI22_X1 port map( A1 => n31233, A2 => n29157, B1 => n31209, B2 => 
                           n29161, ZN => n37177);
   U2543 : AOI22_X1 port map( A1 => n31157, A2 => n29164, B1 => n31201, B2 => 
                           n29211, ZN => n37176);
   U2544 : AOI22_X1 port map( A1 => n31221, A2 => n29455, B1 => n31156, B2 => 
                           n29384, ZN => n37175);
   U2545 : AOI22_X1 port map( A1 => n31214, A2 => n29172, B1 => n31217, B2 => 
                           n29119, ZN => n37174);
   U2546 : NAND4_X1 port map( A1 => n37177, A2 => n37176, A3 => n37175, A4 => 
                           n37174, ZN => n37178);
   U2547 : AOI22_X1 port map( A1 => n37423, A2 => n37179, B1 => n37622, B2 => 
                           n37178, ZN => n37180);
   U2548 : OAI21_X1 port map( B1 => n37627, B2 => n37181, A => n37180, ZN => 
                           OUT2(20));
   U2549 : AOI22_X1 port map( A1 => n30082, A2 => n30003, B1 => n31200, B2 => 
                           n29571, ZN => n37185);
   U2550 : AOI22_X1 port map( A1 => n30083, A2 => n29972, B1 => n31203, B2 => 
                           n29991, ZN => n37184);
   U2551 : AOI22_X1 port map( A1 => n30070, A2 => n29505, B1 => n30080, B2 => 
                           n29271, ZN => n37183);
   U2552 : AOI22_X1 port map( A1 => n31225, A2 => n29460, B1 => n31227, B2 => 
                           n29539, ZN => n37182);
   U2553 : NAND4_X1 port map( A1 => n37185, A2 => n37184, A3 => n37183, A4 => 
                           n37182, ZN => n37191);
   U2554 : AOI22_X1 port map( A1 => n30074, A2 => n29551, B1 => n31206, B2 => 
                           n29341, ZN => n37189);
   U2555 : AOI22_X1 port map( A1 => n31213, A2 => n29953, B1 => n30081, B2 => 
                           n30021, ZN => n37188);
   U2556 : AOI22_X1 port map( A1 => n30084, A2 => n29572, B1 => n30078, B2 => 
                           n29558, ZN => n37187);
   U2557 : AOI22_X1 port map( A1 => n31222, A2 => n29980, B1 => n30072, B2 => 
                           n29573, ZN => n37186);
   U2558 : NAND4_X1 port map( A1 => n37189, A2 => n37188, A3 => n37187, A4 => 
                           n37186, ZN => n37190);
   U2559 : NOR2_X1 port map( A1 => n37191, A2 => n37190, ZN => n37203);
   U2560 : AOI22_X1 port map( A1 => n31216, A2 => n29837, B1 => n31201, B2 => 
                           n29835, ZN => n37195);
   U2561 : AOI22_X1 port map( A1 => n31214, A2 => n29834, B1 => n31162, B2 => 
                           n29851, ZN => n37194);
   U2562 : AOI22_X1 port map( A1 => n31168, A2 => n29838, B1 => n31215, B2 => 
                           n29836, ZN => n37193);
   U2563 : AOI22_X1 port map( A1 => n31219, A2 => n29866, B1 => n31157, B2 => 
                           n29854, ZN => n37192);
   U2564 : NAND4_X1 port map( A1 => n37195, A2 => n37194, A3 => n37193, A4 => 
                           n37192, ZN => n37201);
   U2565 : AOI22_X1 port map( A1 => n31216, A2 => n29596, B1 => n31209, B2 => 
                           n29688, ZN => n37199);
   U2566 : AOI22_X1 port map( A1 => n31156, A2 => n29385, B1 => n31157, B2 => 
                           n29685, ZN => n37198);
   U2567 : AOI22_X1 port map( A1 => n31214, A2 => n29363, B1 => n31201, B2 => 
                           n29417, ZN => n37197);
   U2568 : AOI22_X1 port map( A1 => n31162, A2 => n29454, B1 => n31165, B2 => 
                           n29690, ZN => n37196);
   U2569 : NAND4_X1 port map( A1 => n37199, A2 => n37198, A3 => n37197, A4 => 
                           n37196, ZN => n37200);
   U2570 : AOI22_X1 port map( A1 => n37423, A2 => n37201, B1 => n37622, B2 => 
                           n37200, ZN => n37202);
   U2571 : OAI21_X1 port map( B1 => n37627, B2 => n37203, A => n37202, ZN => 
                           OUT2(19));
   U2572 : AOI22_X1 port map( A1 => n30076, A2 => n29470, B1 => n30077, B2 => 
                           n29540, ZN => n37207);
   U2573 : AOI22_X1 port map( A1 => n31228, A2 => n29552, B1 => n30075, B2 => 
                           n29979, ZN => n37206);
   U2574 : AOI22_X1 port map( A1 => n30069, A2 => n29333, B1 => n31203, B2 => 
                           n29995, ZN => n37205);
   U2575 : AOI22_X1 port map( A1 => n30072, A2 => n29561, B1 => n31205, B2 => 
                           n29974, ZN => n37204);
   U2576 : NAND4_X1 port map( A1 => n37207, A2 => n37206, A3 => n37205, A4 => 
                           n37204, ZN => n37213);
   U2577 : AOI22_X1 port map( A1 => n30082, A2 => n30004, B1 => n30078, B2 => 
                           n29559, ZN => n37211);
   U2578 : AOI22_X1 port map( A1 => n30071, A2 => n29562, B1 => n31223, B2 => 
                           n29504, ZN => n37210);
   U2579 : AOI22_X1 port map( A1 => n31226, A2 => n29270, B1 => n31213, B2 => 
                           n29956, ZN => n37209);
   U2580 : AOI22_X1 port map( A1 => n30084, A2 => n29563, B1 => n30081, B2 => 
                           n30024, ZN => n37208);
   U2581 : NAND4_X1 port map( A1 => n37211, A2 => n37210, A3 => n37209, A4 => 
                           n37208, ZN => n37212);
   U2582 : NOR2_X1 port map( A1 => n37213, A2 => n37212, ZN => n37225);
   U2583 : CLKBUF_X1 port map( A => n37378, Z => n37624);
   U2584 : AOI22_X1 port map( A1 => n31208, A2 => n29841, B1 => n31202, B2 => 
                           n29839, ZN => n37217);
   U2585 : AOI22_X1 port map( A1 => n31214, A2 => n29840, B1 => n31209, B2 => 
                           n29844, ZN => n37216);
   U2586 : AOI22_X1 port map( A1 => n31219, A2 => n29881, B1 => n31155, B2 => 
                           n29843, ZN => n37215);
   U2587 : AOI22_X1 port map( A1 => n31162, A2 => n29842, B1 => n31157, B2 => 
                           n29845, ZN => n37214);
   U2588 : NAND4_X1 port map( A1 => n37217, A2 => n37216, A3 => n37215, A4 => 
                           n37214, ZN => n37223);
   U2589 : AOI22_X1 port map( A1 => n31233, A2 => n29709, B1 => n31208, B2 => 
                           n29416, ZN => n37221);
   U2590 : AOI22_X1 port map( A1 => n31218, A2 => n29679, B1 => n31220, B2 => 
                           n29362, ZN => n37220);
   U2591 : AOI22_X1 port map( A1 => n31155, A2 => n29584, B1 => n31156, B2 => 
                           n29386, ZN => n37219);
   U2592 : AOI22_X1 port map( A1 => n31168, A2 => n29689, B1 => n31162, B2 => 
                           n29452, ZN => n37218);
   U2593 : NAND4_X1 port map( A1 => n37221, A2 => n37220, A3 => n37219, A4 => 
                           n37218, ZN => n37222);
   U2594 : AOI22_X1 port map( A1 => n37624, A2 => n37223, B1 => n37622, B2 => 
                           n37222, ZN => n37224);
   U2595 : OAI21_X1 port map( B1 => n37627, B2 => n37225, A => n37224, ZN => 
                           OUT2(18));
   U2596 : AOI22_X1 port map( A1 => n30081, A2 => n30026, B1 => n31199, B2 => 
                           n29318, ZN => n37229);
   U2597 : AOI22_X1 port map( A1 => n31222, A2 => n29969, B1 => n30074, B2 => 
                           n29319, ZN => n37228);
   U2598 : AOI22_X1 port map( A1 => n30083, A2 => n29976, B1 => n31212, B2 => 
                           n29322, ZN => n37227);
   U2599 : AOI22_X1 port map( A1 => n30073, A2 => n30008, B1 => n30079, B2 => 
                           n30001, ZN => n37226);
   U2600 : NAND4_X1 port map( A1 => n37229, A2 => n37228, A3 => n37227, A4 => 
                           n37226, ZN => n37235);
   U2601 : AOI22_X1 port map( A1 => n31226, A2 => n29282, B1 => n30070, B2 => 
                           n29321, ZN => n37233);
   U2602 : AOI22_X1 port map( A1 => n30069, A2 => n29310, B1 => n30071, B2 => 
                           n29325, ZN => n37232);
   U2603 : AOI22_X1 port map( A1 => n31227, A2 => n29320, B1 => n30082, B2 => 
                           n30005, ZN => n37231);
   U2604 : AOI22_X1 port map( A1 => n30084, A2 => n29323, B1 => n30076, B2 => 
                           n29311, ZN => n37230);
   U2605 : NAND4_X1 port map( A1 => n37233, A2 => n37232, A3 => n37231, A4 => 
                           n37230, ZN => n37234);
   U2606 : NOR2_X1 port map( A1 => n37235, A2 => n37234, ZN => n37247);
   U2607 : AOI22_X1 port map( A1 => n31168, A2 => n29765, B1 => n31208, B2 => 
                           n29764, ZN => n37239);
   U2608 : AOI22_X1 port map( A1 => n31215, A2 => n29768, B1 => n31210, B2 => 
                           n29766, ZN => n37238);
   U2609 : AOI22_X1 port map( A1 => n31219, A2 => n29873, B1 => n31216, B2 => 
                           n29774, ZN => n37237);
   U2610 : AOI22_X1 port map( A1 => n31220, A2 => n29770, B1 => n31162, B2 => 
                           n29772, ZN => n37236);
   U2611 : NAND4_X1 port map( A1 => n37239, A2 => n37238, A3 => n37237, A4 => 
                           n37236, ZN => n37245);
   U2612 : AOI22_X1 port map( A1 => n31156, A2 => n29312, B1 => n31214, B2 => 
                           n29313, ZN => n37243);
   U2613 : AOI22_X1 port map( A1 => n31162, A2 => n29315, B1 => n31208, B2 => 
                           n29314, ZN => n37242);
   U2614 : AOI22_X1 port map( A1 => n31219, A2 => n29145, B1 => n31155, B2 => 
                           n29118, ZN => n37241);
   U2615 : AOI22_X1 port map( A1 => n31157, A2 => n29163, B1 => n31209, B2 => 
                           n29160, ZN => n37240);
   U2616 : NAND4_X1 port map( A1 => n37243, A2 => n37242, A3 => n37241, A4 => 
                           n37240, ZN => n37244);
   U2617 : AOI22_X1 port map( A1 => n37624, A2 => n37245, B1 => n37622, B2 => 
                           n37244, ZN => n37246);
   U2618 : OAI21_X1 port map( B1 => n37627, B2 => n37247, A => n37246, ZN => 
                           OUT2(17));
   U2619 : AOI22_X1 port map( A1 => n30072, A2 => n29285, B1 => n30080, B2 => 
                           n29268, ZN => n37251);
   U2620 : AOI22_X1 port map( A1 => n31228, A2 => n29279, B1 => n31227, B2 => 
                           n29280, ZN => n37250);
   U2621 : AOI22_X1 port map( A1 => n30084, A2 => n29265, B1 => n30078, B2 => 
                           n29277, ZN => n37249);
   U2622 : AOI22_X1 port map( A1 => n30083, A2 => n29977, B1 => n30076, B2 => 
                           n29290, ZN => n37248);
   U2623 : NAND4_X1 port map( A1 => n37251, A2 => n37250, A3 => n37249, A4 => 
                           n37248, ZN => n37257);
   U2624 : AOI22_X1 port map( A1 => n30069, A2 => n29289, B1 => n30082, B2 => 
                           n30006, ZN => n37255);
   U2625 : AOI22_X1 port map( A1 => n31224, A2 => n29975, B1 => n31213, B2 => 
                           n29949, ZN => n37254);
   U2626 : AOI22_X1 port map( A1 => n30079, A2 => n30009, B1 => n30075, B2 => 
                           n29967, ZN => n37253);
   U2627 : AOI22_X1 port map( A1 => n30071, A2 => n29264, B1 => n31223, B2 => 
                           n29291, ZN => n37252);
   U2628 : NAND4_X1 port map( A1 => n37255, A2 => n37254, A3 => n37253, A4 => 
                           n37252, ZN => n37256);
   U2629 : NOR2_X1 port map( A1 => n37257, A2 => n37256, ZN => n37269);
   U2630 : AOI22_X1 port map( A1 => n31218, A2 => n29863, B1 => n31208, B2 => 
                           n29859, ZN => n37261);
   U2631 : AOI22_X1 port map( A1 => n31156, A2 => n29856, B1 => n31214, B2 => 
                           n29858, ZN => n37260);
   U2632 : AOI22_X1 port map( A1 => n31155, A2 => n29861, B1 => n31162, B2 => 
                           n29860, ZN => n37259);
   U2633 : AOI22_X1 port map( A1 => n30050, A2 => n29862, B1 => n31165, B2 => 
                           n29769, ZN => n37258);
   U2634 : NAND4_X1 port map( A1 => n37261, A2 => n37260, A3 => n37259, A4 => 
                           n37258, ZN => n37267);
   U2635 : AOI22_X1 port map( A1 => n31156, A2 => n29292, B1 => n31233, B2 => 
                           n29697, ZN => n37265);
   U2636 : AOI22_X1 port map( A1 => n31155, A2 => n29586, B1 => n31158, B2 => 
                           n29294, ZN => n37264);
   U2637 : AOI22_X1 port map( A1 => n31168, A2 => n29693, B1 => n31214, B2 => 
                           n29293, ZN => n37263);
   U2638 : AOI22_X1 port map( A1 => n31218, A2 => n29680, B1 => n31162, B2 => 
                           n29295, ZN => n37262);
   U2639 : NAND4_X1 port map( A1 => n37265, A2 => n37264, A3 => n37263, A4 => 
                           n37262, ZN => n37266);
   U2640 : AOI22_X1 port map( A1 => n37423, A2 => n37267, B1 => n37622, B2 => 
                           n37266, ZN => n37268);
   U2641 : OAI21_X1 port map( B1 => n37627, B2 => n37269, A => n37268, ZN => 
                           OUT2(16));
   U2642 : AOI22_X1 port map( A1 => n31227, A2 => n29527, B1 => n30072, B2 => 
                           n29524, ZN => n37273);
   U2643 : AOI22_X1 port map( A1 => n30069, A2 => n29332, B1 => n30078, B2 => 
                           n29525, ZN => n37272);
   U2644 : AOI22_X1 port map( A1 => n30073, A2 => n29954, B1 => n31205, B2 => 
                           n29978, ZN => n37271);
   U2645 : AOI22_X1 port map( A1 => n30080, A2 => n29269, B1 => n31207, B2 => 
                           n30007, ZN => n37270);
   U2646 : NAND4_X1 port map( A1 => n37273, A2 => n37272, A3 => n37271, A4 => 
                           n37270, ZN => n37279);
   U2647 : AOI22_X1 port map( A1 => n30070, A2 => n29503, B1 => n30081, B2 => 
                           n30027, ZN => n37277);
   U2648 : AOI22_X1 port map( A1 => n30084, A2 => n29528, B1 => n30071, B2 => 
                           n29529, ZN => n37276);
   U2649 : AOI22_X1 port map( A1 => n31225, A2 => n29471, B1 => n31203, B2 => 
                           n30002, ZN => n37275);
   U2650 : AOI22_X1 port map( A1 => n30074, A2 => n29526, B1 => n30075, B2 => 
                           n29965, ZN => n37274);
   U2651 : NAND4_X1 port map( A1 => n37277, A2 => n37276, A3 => n37275, A4 => 
                           n37274, ZN => n37278);
   U2652 : NOR2_X1 port map( A1 => n37279, A2 => n37278, ZN => n37291);
   U2653 : AOI22_X1 port map( A1 => n31208, A2 => n29812, B1 => n31217, B2 => 
                           n29821, ZN => n37283);
   U2654 : AOI22_X1 port map( A1 => n31156, A2 => n29816, B1 => n31214, B2 => 
                           n29815, ZN => n37282);
   U2655 : AOI22_X1 port map( A1 => n31162, A2 => n29811, B1 => n31210, B2 => 
                           n29799, ZN => n37281);
   U2656 : AOI22_X1 port map( A1 => n31209, A2 => n29810, B1 => n31165, B2 => 
                           n29904, ZN => n37280);
   U2657 : NAND4_X1 port map( A1 => n37283, A2 => n37282, A3 => n37281, A4 => 
                           n37280, ZN => n37289);
   U2658 : AOI22_X1 port map( A1 => n31155, A2 => n29122, B1 => n31208, B2 => 
                           n29415, ZN => n37287);
   U2659 : AOI22_X1 port map( A1 => n31214, A2 => n29361, B1 => n31209, B2 => 
                           n29146, ZN => n37286);
   U2660 : AOI22_X1 port map( A1 => n31157, A2 => n29162, B1 => n31165, B2 => 
                           n29148, ZN => n37285);
   U2661 : AOI22_X1 port map( A1 => n31162, A2 => n29451, B1 => n31202, B2 => 
                           n29387, ZN => n37284);
   U2662 : NAND4_X1 port map( A1 => n37287, A2 => n37286, A3 => n37285, A4 => 
                           n37284, ZN => n37288);
   U2663 : AOI22_X1 port map( A1 => n37423, A2 => n37289, B1 => n37622, B2 => 
                           n37288, ZN => n37290);
   U2664 : OAI21_X1 port map( B1 => n37627, B2 => n37291, A => n37290, ZN => 
                           OUT2(15));
   U2665 : AOI22_X1 port map( A1 => n31228, A2 => n29553, B1 => n31224, B2 => 
                           n30020, ZN => n37295);
   U2666 : AOI22_X1 port map( A1 => n30073, A2 => n29942, B1 => n30070, B2 => 
                           n29502, ZN => n37294);
   U2667 : AOI22_X1 port map( A1 => n30080, A2 => n29266, B1 => n31199, B2 => 
                           n29560, ZN => n37293);
   U2668 : AOI22_X1 port map( A1 => n31225, A2 => n29473, B1 => n30072, B2 => 
                           n29523, ZN => n37292);
   U2669 : NAND4_X1 port map( A1 => n37295, A2 => n37294, A3 => n37293, A4 => 
                           n37292, ZN => n37301);
   U2670 : AOI22_X1 port map( A1 => n30082, A2 => n30011, B1 => n31203, B2 => 
                           n30000, ZN => n37299);
   U2671 : AOI22_X1 port map( A1 => n31222, A2 => n29963, B1 => n31211, B2 => 
                           n29577, ZN => n37298);
   U2672 : AOI22_X1 port map( A1 => n31227, A2 => n29544, B1 => n30083, B2 => 
                           n29986, ZN => n37297);
   U2673 : AOI22_X1 port map( A1 => n30069, A2 => n29331, B1 => n30071, B2 => 
                           n29574, ZN => n37296);
   U2674 : NAND4_X1 port map( A1 => n37299, A2 => n37298, A3 => n37297, A4 => 
                           n37296, ZN => n37300);
   U2675 : NOR2_X1 port map( A1 => n37301, A2 => n37300, ZN => n37313);
   U2676 : AOI22_X1 port map( A1 => n31209, A2 => n29908, B1 => n31165, B2 => 
                           n29778, ZN => n37305);
   U2677 : AOI22_X1 port map( A1 => n31155, A2 => n29901, B1 => n31201, B2 => 
                           n29903, ZN => n37304);
   U2678 : AOI22_X1 port map( A1 => n31161, A2 => n29905, B1 => n31210, B2 => 
                           n29907, ZN => n37303);
   U2679 : AOI22_X1 port map( A1 => n31162, A2 => n29902, B1 => n31202, B2 => 
                           n29906, ZN => n37302);
   U2680 : NAND4_X1 port map( A1 => n37305, A2 => n37304, A3 => n37303, A4 => 
                           n37302, ZN => n37311);
   U2681 : AOI22_X1 port map( A1 => n31155, A2 => n29578, B1 => n31158, B2 => 
                           n29408, ZN => n37309);
   U2682 : AOI22_X1 port map( A1 => n31162, A2 => n29448, B1 => n31157, B2 => 
                           n29672, ZN => n37308);
   U2683 : AOI22_X1 port map( A1 => n31168, A2 => n29695, B1 => n31202, B2 => 
                           n29388, ZN => n37307);
   U2684 : AOI22_X1 port map( A1 => n31233, A2 => n29674, B1 => n31214, B2 => 
                           n29360, ZN => n37306);
   U2685 : NAND4_X1 port map( A1 => n37309, A2 => n37308, A3 => n37307, A4 => 
                           n37306, ZN => n37310);
   U2686 : AOI22_X1 port map( A1 => n37423, A2 => n37311, B1 => n37622, B2 => 
                           n37310, ZN => n37312);
   U2687 : OAI21_X1 port map( B1 => n37627, B2 => n37313, A => n37312, ZN => 
                           OUT2(14));
   U2688 : AOI22_X1 port map( A1 => n31225, A2 => n29474, B1 => n30070, B2 => 
                           n29501, ZN => n37317);
   U2689 : AOI22_X1 port map( A1 => n31213, A2 => n29941, B1 => n31200, B2 => 
                           n29520, ZN => n37316);
   U2690 : AOI22_X1 port map( A1 => n31222, A2 => n29961, B1 => n30074, B2 => 
                           n29516, ZN => n37315);
   U2691 : AOI22_X1 port map( A1 => n30079, A2 => n29998, B1 => n31205, B2 => 
                           n29987, ZN => n37314);
   U2692 : NAND4_X1 port map( A1 => n37317, A2 => n37316, A3 => n37315, A4 => 
                           n37314, ZN => n37323);
   U2693 : AOI22_X1 port map( A1 => n30084, A2 => n29519, B1 => n31212, B2 => 
                           n29518, ZN => n37321);
   U2694 : AOI22_X1 port map( A1 => n31207, A2 => n30012, B1 => n31199, B2 => 
                           n29515, ZN => n37320);
   U2695 : AOI22_X1 port map( A1 => n31226, A2 => n29267, B1 => n31224, B2 => 
                           n29958, ZN => n37319);
   U2696 : AOI22_X1 port map( A1 => n30077, A2 => n29517, B1 => n31206, B2 => 
                           n29329, ZN => n37318);
   U2697 : NAND4_X1 port map( A1 => n37321, A2 => n37320, A3 => n37319, A4 => 
                           n37318, ZN => n37322);
   U2698 : NOR2_X1 port map( A1 => n37323, A2 => n37322, ZN => n37335);
   U2699 : AOI22_X1 port map( A1 => n31217, A2 => n29885, B1 => n31202, B2 => 
                           n29892, ZN => n37327);
   U2700 : AOI22_X1 port map( A1 => n31157, A2 => n29887, B1 => n31165, B2 => 
                           n29888, ZN => n37326);
   U2701 : AOI22_X1 port map( A1 => n31158, A2 => n29894, B1 => n31161, B2 => 
                           n29893, ZN => n37325);
   U2702 : AOI22_X1 port map( A1 => n31168, A2 => n29886, B1 => n31221, B2 => 
                           n29884, ZN => n37324);
   U2703 : NAND4_X1 port map( A1 => n37327, A2 => n37326, A3 => n37325, A4 => 
                           n37324, ZN => n37333);
   U2704 : AOI22_X1 port map( A1 => n31157, A2 => n29701, B1 => n31209, B2 => 
                           n29708, ZN => n37331);
   U2705 : AOI22_X1 port map( A1 => n31214, A2 => n29359, B1 => n31216, B2 => 
                           n29585, ZN => n37330);
   U2706 : AOI22_X1 port map( A1 => n31158, A2 => n29405, B1 => n31202, B2 => 
                           n29394, ZN => n37329);
   U2707 : AOI22_X1 port map( A1 => n31221, A2 => n29447, B1 => n31165, B2 => 
                           n29691, ZN => n37328);
   U2708 : NAND4_X1 port map( A1 => n37331, A2 => n37330, A3 => n37329, A4 => 
                           n37328, ZN => n37332);
   U2709 : AOI22_X1 port map( A1 => n37423, A2 => n37333, B1 => n37622, B2 => 
                           n37332, ZN => n37334);
   U2710 : OAI21_X1 port map( B1 => n37627, B2 => n37335, A => n37334, ZN => 
                           OUT2(13));
   U2711 : AOI22_X1 port map( A1 => n30080, A2 => n29263, B1 => n31200, B2 => 
                           n29513, ZN => n37339);
   U2712 : AOI22_X1 port map( A1 => n30079, A2 => n29997, B1 => n31199, B2 => 
                           n29508, ZN => n37338);
   U2713 : AOI22_X1 port map( A1 => n30073, A2 => n29959, B1 => n30077, B2 => 
                           n29510, ZN => n37337);
   U2714 : AOI22_X1 port map( A1 => n30083, A2 => n29989, B1 => n30075, B2 => 
                           n29947, ZN => n37336);
   U2715 : NAND4_X1 port map( A1 => n37339, A2 => n37338, A3 => n37337, A4 => 
                           n37336, ZN => n37345);
   U2716 : AOI22_X1 port map( A1 => n31224, A2 => n29955, B1 => n31211, B2 => 
                           n29512, ZN => n37343);
   U2717 : AOI22_X1 port map( A1 => n31223, A2 => n29500, B1 => n30076, B2 => 
                           n29475, ZN => n37342);
   U2718 : AOI22_X1 port map( A1 => n30082, A2 => n30013, B1 => n31212, B2 => 
                           n29511, ZN => n37341);
   U2719 : AOI22_X1 port map( A1 => n30069, A2 => n29328, B1 => n30074, B2 => 
                           n29509, ZN => n37340);
   U2720 : NAND4_X1 port map( A1 => n37343, A2 => n37342, A3 => n37341, A4 => 
                           n37340, ZN => n37344);
   U2721 : NOR2_X1 port map( A1 => n37345, A2 => n37344, ZN => n37357);
   U2722 : AOI22_X1 port map( A1 => n31161, A2 => n29883, B1 => n31202, B2 => 
                           n29882, ZN => n37349);
   U2723 : AOI22_X1 port map( A1 => n31168, A2 => n29877, B1 => n31210, B2 => 
                           n29878, ZN => n37348);
   U2724 : AOI22_X1 port map( A1 => n31219, A2 => n29879, B1 => n31155, B2 => 
                           n29876, ZN => n37347);
   U2725 : AOI22_X1 port map( A1 => n31158, A2 => n29874, B1 => n31221, B2 => 
                           n29875, ZN => n37346);
   U2726 : NAND4_X1 port map( A1 => n37349, A2 => n37348, A3 => n37347, A4 => 
                           n37346, ZN => n37355);
   U2727 : AOI22_X1 port map( A1 => n31157, A2 => n29669, B1 => n31217, B2 => 
                           n29593, ZN => n37353);
   U2728 : AOI22_X1 port map( A1 => n31214, A2 => n29358, B1 => n31215, B2 => 
                           n29395, ZN => n37352);
   U2729 : AOI22_X1 port map( A1 => n31158, A2 => n29404, B1 => n31165, B2 => 
                           n29670, ZN => n37351);
   U2730 : AOI22_X1 port map( A1 => n31168, A2 => n29699, B1 => n31221, B2 => 
                           n29446, ZN => n37350);
   U2731 : NAND4_X1 port map( A1 => n37353, A2 => n37352, A3 => n37351, A4 => 
                           n37350, ZN => n37354);
   U2732 : AOI22_X1 port map( A1 => n37423, A2 => n37355, B1 => n37622, B2 => 
                           n37354, ZN => n37356);
   U2733 : OAI21_X1 port map( B1 => n37627, B2 => n37357, A => n37356, ZN => 
                           OUT2(12));
   U2734 : AOI22_X1 port map( A1 => n30073, A2 => n29943, B1 => n31211, B2 => 
                           n29498, ZN => n37361);
   U2735 : AOI22_X1 port map( A1 => n30079, A2 => n29996, B1 => n30074, B2 => 
                           n29494, ZN => n37360);
   U2736 : AOI22_X1 port map( A1 => n30077, A2 => n29495, B1 => n31205, B2 => 
                           n29990, ZN => n37359);
   U2737 : AOI22_X1 port map( A1 => n31223, A2 => n29496, B1 => n30076, B2 => 
                           n29476, ZN => n37358);
   U2738 : NAND4_X1 port map( A1 => n37361, A2 => n37360, A3 => n37359, A4 => 
                           n37358, ZN => n37367);
   U2739 : AOI22_X1 port map( A1 => n31207, A2 => n30014, B1 => n31206, B2 => 
                           n29327, ZN => n37365);
   U2740 : AOI22_X1 port map( A1 => n30080, A2 => n29324, B1 => n30081, B2 => 
                           n29951, ZN => n37364);
   U2741 : AOI22_X1 port map( A1 => n30071, A2 => n29499, B1 => n30075, B2 => 
                           n29971, ZN => n37363);
   U2742 : AOI22_X1 port map( A1 => n30072, A2 => n29497, B1 => n30078, B2 => 
                           n29493, ZN => n37362);
   U2743 : NAND4_X1 port map( A1 => n37365, A2 => n37364, A3 => n37363, A4 => 
                           n37362, ZN => n37366);
   U2744 : NOR2_X1 port map( A1 => n37367, A2 => n37366, ZN => n37380);
   U2745 : AOI22_X1 port map( A1 => n31168, A2 => n29868, B1 => n31233, B2 => 
                           n29870, ZN => n37371);
   U2746 : AOI22_X1 port map( A1 => n31221, A2 => n29865, B1 => n31156, B2 => 
                           n29871, ZN => n37370);
   U2747 : AOI22_X1 port map( A1 => n31216, A2 => n29867, B1 => n31161, B2 => 
                           n29857, ZN => n37369);
   U2748 : AOI22_X1 port map( A1 => n31158, A2 => n29864, B1 => n31157, B2 => 
                           n29869, ZN => n37368);
   U2749 : NAND4_X1 port map( A1 => n37371, A2 => n37370, A3 => n37369, A4 => 
                           n37368, ZN => n37377);
   U2750 : AOI22_X1 port map( A1 => n31219, A2 => n29683, B1 => n31161, B2 => 
                           n29357, ZN => n37375);
   U2751 : AOI22_X1 port map( A1 => n31155, A2 => n29592, B1 => n31210, B2 => 
                           n29703, ZN => n37374);
   U2752 : AOI22_X1 port map( A1 => n31168, A2 => n29700, B1 => n31158, B2 => 
                           n29399, ZN => n37373);
   U2753 : AOI22_X1 port map( A1 => n31221, A2 => n29445, B1 => n31215, B2 => 
                           n29396, ZN => n37372);
   U2754 : NAND4_X1 port map( A1 => n37375, A2 => n37374, A3 => n37373, A4 => 
                           n37372, ZN => n37376);
   U2755 : AOI22_X1 port map( A1 => n37378, A2 => n37377, B1 => n37622, B2 => 
                           n37376, ZN => n37379);
   U2756 : OAI21_X1 port map( B1 => n37448, B2 => n37380, A => n37379, ZN => 
                           OUT2(11));
   U2757 : AOI22_X1 port map( A1 => n30069, A2 => n29326, B1 => n31222, B2 => 
                           n29714, ZN => n37384);
   U2758 : AOI22_X1 port map( A1 => n30074, A2 => n29486, B1 => n31207, B2 => 
                           n29719, ZN => n37383);
   U2759 : AOI22_X1 port map( A1 => n31224, A2 => n29717, B1 => n30077, B2 => 
                           n29487, ZN => n37382);
   U2760 : AOI22_X1 port map( A1 => n31212, A2 => n29489, B1 => n31200, B2 => 
                           n29490, ZN => n37381);
   U2761 : NAND4_X1 port map( A1 => n37384, A2 => n37383, A3 => n37382, A4 => 
                           n37381, ZN => n37390);
   U2762 : AOI22_X1 port map( A1 => n30078, A2 => n29485, B1 => n30070, B2 => 
                           n29488, ZN => n37388);
   U2763 : AOI22_X1 port map( A1 => n30073, A2 => n29715, B1 => n30076, B2 => 
                           n29477, ZN => n37387);
   U2764 : AOI22_X1 port map( A1 => n30084, A2 => n29251, B1 => n30079, B2 => 
                           n29716, ZN => n37386);
   U2765 : AOI22_X1 port map( A1 => n30083, A2 => n29718, B1 => n30080, B2 => 
                           n29530, ZN => n37385);
   U2766 : NAND4_X1 port map( A1 => n37388, A2 => n37387, A3 => n37386, A4 => 
                           n37385, ZN => n37389);
   U2767 : NOR2_X1 port map( A1 => n37390, A2 => n37389, ZN => n37402);
   U2768 : AOI22_X1 port map( A1 => n31221, A2 => n29253, B1 => n31216, B2 => 
                           n29256, ZN => n37394);
   U2769 : AOI22_X1 port map( A1 => n31158, A2 => n29259, B1 => n31202, B2 => 
                           n29257, ZN => n37393);
   U2770 : AOI22_X1 port map( A1 => n31161, A2 => n29254, B1 => n31209, B2 => 
                           n29252, ZN => n37392);
   U2771 : AOI22_X1 port map( A1 => n31233, A2 => n29250, B1 => n31157, B2 => 
                           n29249, ZN => n37391);
   U2772 : NAND4_X1 port map( A1 => n37394, A2 => n37393, A3 => n37392, A4 => 
                           n37391, ZN => n37400);
   U2773 : AOI22_X1 port map( A1 => n31210, A2 => n29676, B1 => n31209, B2 => 
                           n29710, ZN => n37398);
   U2774 : AOI22_X1 port map( A1 => n31155, A2 => n29590, B1 => n31158, B2 => 
                           n29258, ZN => n37397);
   U2775 : AOI22_X1 port map( A1 => n31221, A2 => n29442, B1 => n31202, B2 => 
                           n29255, ZN => n37396);
   U2776 : AOI22_X1 port map( A1 => n31219, A2 => n29686, B1 => n31161, B2 => 
                           n29354, ZN => n37395);
   U2777 : NAND4_X1 port map( A1 => n37398, A2 => n37397, A3 => n37396, A4 => 
                           n37395, ZN => n37399);
   U2778 : AOI22_X1 port map( A1 => n37423, A2 => n37400, B1 => n37622, B2 => 
                           n37399, ZN => n37401);
   U2779 : OAI21_X1 port map( B1 => n37448, B2 => n37402, A => n37401, ZN => 
                           OUT2(10));
   U2780 : AOI22_X1 port map( A1 => n30071, A2 => n29535, B1 => n30074, B2 => 
                           n29533, ZN => n37406);
   U2781 : AOI22_X1 port map( A1 => n30072, A2 => n29522, B1 => n30083, B2 => 
                           n29992, ZN => n37405);
   U2782 : AOI22_X1 port map( A1 => n31211, A2 => n29531, B1 => n31203, B2 => 
                           n29994, ZN => n37404);
   U2783 : AOI22_X1 port map( A1 => n30082, A2 => n30015, B1 => n30075, B2 => 
                           n29970, ZN => n37403);
   U2784 : NAND4_X1 port map( A1 => n37406, A2 => n37405, A3 => n37404, A4 => 
                           n37403, ZN => n37412);
   U2785 : AOI22_X1 port map( A1 => n31225, A2 => n29478, B1 => n30081, B2 => 
                           n29950, ZN => n37410);
   U2786 : AOI22_X1 port map( A1 => n31226, A2 => n29534, B1 => n31206, B2 => 
                           n29317, ZN => n37409);
   U2787 : AOI22_X1 port map( A1 => n31227, A2 => n29532, B1 => n30078, B2 => 
                           n29484, ZN => n37408);
   U2788 : AOI22_X1 port map( A1 => n30073, A2 => n29962, B1 => n30070, B2 => 
                           n29492, ZN => n37407);
   U2789 : NAND4_X1 port map( A1 => n37410, A2 => n37409, A3 => n37408, A4 => 
                           n37407, ZN => n37411);
   U2790 : NOR2_X1 port map( A1 => n37412, A2 => n37411, ZN => n37425);
   U2791 : AOI22_X1 port map( A1 => n31221, A2 => n29937, B1 => n31215, B2 => 
                           n29934, ZN => n37416);
   U2792 : AOI22_X1 port map( A1 => n31158, A2 => n29935, B1 => n31233, B2 => 
                           n29940, ZN => n37415);
   U2793 : AOI22_X1 port map( A1 => n31210, A2 => n29936, B1 => n31217, B2 => 
                           n29939, ZN => n37414);
   U2794 : AOI22_X1 port map( A1 => n31168, A2 => n29938, B1 => n31161, B2 => 
                           n29933, ZN => n37413);
   U2795 : NAND4_X1 port map( A1 => n37416, A2 => n37415, A3 => n37414, A4 => 
                           n37413, ZN => n37422);
   U2796 : AOI22_X1 port map( A1 => n31165, A2 => n29711, B1 => n31202, B2 => 
                           n29402, ZN => n37420);
   U2797 : AOI22_X1 port map( A1 => n31218, A2 => n29677, B1 => n31220, B2 => 
                           n29355, ZN => n37419);
   U2798 : AOI22_X1 port map( A1 => n31158, A2 => n29398, B1 => n31209, B2 => 
                           n29702, ZN => n37418);
   U2799 : AOI22_X1 port map( A1 => n31155, A2 => n29580, B1 => n31221, B2 => 
                           n29440, ZN => n37417);
   U2800 : NAND4_X1 port map( A1 => n37420, A2 => n37419, A3 => n37418, A4 => 
                           n37417, ZN => n37421);
   U2801 : AOI22_X1 port map( A1 => n37423, A2 => n37422, B1 => n37622, B2 => 
                           n37421, ZN => n37424);
   U2802 : OAI21_X1 port map( B1 => n37448, B2 => n37425, A => n37424, ZN => 
                           OUT2(9));
   U2803 : AOI22_X1 port map( A1 => n31226, A2 => n29545, B1 => n30074, B2 => 
                           n29542, ZN => n37429);
   U2804 : AOI22_X1 port map( A1 => n30082, A2 => n30016, B1 => n30077, B2 => 
                           n29541, ZN => n37428);
   U2805 : AOI22_X1 port map( A1 => n30071, A2 => n29546, B1 => n30081, B2 => 
                           n29948, ZN => n37427);
   U2806 : AOI22_X1 port map( A1 => n30078, A2 => n29543, B1 => n30075, B2 => 
                           n29968, ZN => n37426);
   U2807 : NAND4_X1 port map( A1 => n37429, A2 => n37428, A3 => n37427, A4 => 
                           n37426, ZN => n37435);
   U2808 : AOI22_X1 port map( A1 => n30084, A2 => n29547, B1 => n31203, B2 => 
                           n29985, ZN => n37433);
   U2809 : AOI22_X1 port map( A1 => n30070, A2 => n29491, B1 => n30076, B2 => 
                           n29479, ZN => n37432);
   U2810 : AOI22_X1 port map( A1 => n30069, A2 => n29316, B1 => n31212, B2 => 
                           n29521, ZN => n37431);
   U2811 : AOI22_X1 port map( A1 => n30083, A2 => n29993, B1 => n31213, B2 => 
                           n29973, ZN => n37430);
   U2812 : NAND4_X1 port map( A1 => n37433, A2 => n37432, A3 => n37431, A4 => 
                           n37430, ZN => n37434);
   U2813 : NOR2_X1 port map( A1 => n37435, A2 => n37434, ZN => n37447);
   U2814 : AOI22_X1 port map( A1 => n31168, A2 => n29923, B1 => n31220, B2 => 
                           n29918, ZN => n37439);
   U2815 : AOI22_X1 port map( A1 => n31221, A2 => n29924, B1 => n31165, B2 => 
                           n29922, ZN => n37438);
   U2816 : AOI22_X1 port map( A1 => n31208, A2 => n29919, B1 => n31217, B2 => 
                           n29920, ZN => n37437);
   U2817 : AOI22_X1 port map( A1 => n31218, A2 => n29921, B1 => n31202, B2 => 
                           n29925, ZN => n37436);
   U2818 : NAND4_X1 port map( A1 => n37439, A2 => n37438, A3 => n37437, A4 => 
                           n37436, ZN => n37445);
   U2819 : AOI22_X1 port map( A1 => n31220, A2 => n29356, B1 => n31158, B2 => 
                           n29397, ZN => n37443);
   U2820 : AOI22_X1 port map( A1 => n31233, A2 => n29678, B1 => n31215, B2 => 
                           n29403, ZN => n37442);
   U2821 : AOI22_X1 port map( A1 => n31221, A2 => n29438, B1 => n31217, B2 => 
                           n29582, ZN => n37441);
   U2822 : AOI22_X1 port map( A1 => n31218, A2 => n29673, B1 => n30050, B2 => 
                           n29705, ZN => n37440);
   U2823 : NAND4_X1 port map( A1 => n37443, A2 => n37442, A3 => n37441, A4 => 
                           n37440, ZN => n37444);
   U2824 : AOI22_X1 port map( A1 => n37624, A2 => n37445, B1 => n37622, B2 => 
                           n37444, ZN => n37446);
   U2825 : OAI21_X1 port map( B1 => n37448, B2 => n37447, A => n37446, ZN => 
                           OUT2(8));
   U2826 : AOI22_X1 port map( A1 => n30084, A2 => n29018, B1 => n31199, B2 => 
                           n29023, ZN => n37452);
   U2827 : AOI22_X1 port map( A1 => n31228, A2 => n29024, B1 => n31224, B2 => 
                           n29665, ZN => n37451);
   U2828 : AOI22_X1 port map( A1 => n30082, A2 => n29667, B1 => n30083, B2 => 
                           n29666, ZN => n37450);
   U2829 : AOI22_X1 port map( A1 => n31223, A2 => n29035, B1 => n30080, B2 => 
                           n29020, ZN => n37449);
   U2830 : NAND4_X1 port map( A1 => n37452, A2 => n37451, A3 => n37450, A4 => 
                           n37449, ZN => n37458);
   U2831 : AOI22_X1 port map( A1 => n31222, A2 => n29668, B1 => n31200, B2 => 
                           n29028, ZN => n37456);
   U2832 : AOI22_X1 port map( A1 => n30072, A2 => n29019, B1 => n30077, B2 => 
                           n29033, ZN => n37455);
   U2833 : AOI22_X1 port map( A1 => n30069, A2 => n29038, B1 => n30076, B2 => 
                           n29047, ZN => n37454);
   U2834 : AOI22_X1 port map( A1 => n30073, A2 => n29664, B1 => n30079, B2 => 
                           n29663, ZN => n37453);
   U2835 : NAND4_X1 port map( A1 => n37456, A2 => n37455, A3 => n37454, A4 => 
                           n37453, ZN => n37457);
   U2836 : NOR2_X1 port map( A1 => n37458, A2 => n37457, ZN => n37470);
   U2837 : AOI22_X1 port map( A1 => n30050, A2 => n29237, B1 => n31208, B2 => 
                           n29239, ZN => n37462);
   U2838 : AOI22_X1 port map( A1 => n31215, A2 => n29245, B1 => n31161, B2 => 
                           n29246, ZN => n37461);
   U2839 : AOI22_X1 port map( A1 => n31204, A2 => n29247, B1 => n31217, B2 => 
                           n29236, ZN => n37460);
   U2840 : AOI22_X1 port map( A1 => n31219, A2 => n29233, B1 => n31218, B2 => 
                           n29244, ZN => n37459);
   U2841 : NAND4_X1 port map( A1 => n37462, A2 => n37461, A3 => n37460, A4 => 
                           n37459, ZN => n37468);
   U2842 : AOI22_X1 port map( A1 => n31168, A2 => n29150, B1 => n31208, B2 => 
                           n29111, ZN => n37466);
   U2843 : AOI22_X1 port map( A1 => n31156, A2 => n29086, B1 => n31217, B2 => 
                           n29124, ZN => n37465);
   U2844 : AOI22_X1 port map( A1 => n31165, A2 => n29155, B1 => n31204, B2 => 
                           n29021, ZN => n37464);
   U2845 : AOI22_X1 port map( A1 => n31218, A2 => n29152, B1 => n31220, B2 => 
                           n29114, ZN => n37463);
   U2846 : NAND4_X1 port map( A1 => n37466, A2 => n37465, A3 => n37464, A4 => 
                           n37463, ZN => n37467);
   U2847 : AOI22_X1 port map( A1 => n37624, A2 => n37468, B1 => n37622, B2 => 
                           n37467, ZN => n37469);
   U2848 : OAI21_X1 port map( B1 => n37627, B2 => n37470, A => n37469, ZN => 
                           OUT2(7));
   U2849 : AOI22_X1 port map( A1 => n30082, A2 => n29728, B1 => n30077, B2 => 
                           n29026, ZN => n37474);
   U2850 : AOI22_X1 port map( A1 => n30079, A2 => n29726, B1 => n30081, B2 => 
                           n29754, ZN => n37473);
   U2851 : AOI22_X1 port map( A1 => n31228, A2 => n29050, B1 => n30080, B2 => 
                           n29022, ZN => n37472);
   U2852 : AOI22_X1 port map( A1 => n30069, A2 => n29044, B1 => n31211, B2 => 
                           n29049, ZN => n37471);
   U2853 : NAND4_X1 port map( A1 => n37474, A2 => n37473, A3 => n37472, A4 => 
                           n37471, ZN => n37480);
   U2854 : AOI22_X1 port map( A1 => n30072, A2 => n29051, B1 => n31223, B2 => 
                           n29054, ZN => n37478);
   U2855 : AOI22_X1 port map( A1 => n30075, A2 => n29744, B1 => n31200, B2 => 
                           n29048, ZN => n37477);
   U2856 : AOI22_X1 port map( A1 => n31213, A2 => n29745, B1 => n30076, B2 => 
                           n29041, ZN => n37476);
   U2857 : AOI22_X1 port map( A1 => n31205, A2 => n29736, B1 => n31199, B2 => 
                           n29029, ZN => n37475);
   U2858 : NAND4_X1 port map( A1 => n37478, A2 => n37477, A3 => n37476, A4 => 
                           n37475, ZN => n37479);
   U2859 : NOR2_X1 port map( A1 => n37480, A2 => n37479, ZN => n37492);
   U2860 : AOI22_X1 port map( A1 => n31209, A2 => n29813, B1 => n31208, B2 => 
                           n29820, ZN => n37484);
   U2861 : AOI22_X1 port map( A1 => n31218, A2 => n29805, B1 => n31165, B2 => 
                           n29784, ZN => n37483);
   U2862 : AOI22_X1 port map( A1 => n31156, A2 => n29818, B1 => n31204, B2 => 
                           n29822, ZN => n37482);
   U2863 : AOI22_X1 port map( A1 => n31220, A2 => n29819, B1 => n31217, B2 => 
                           n29823, ZN => n37481);
   U2864 : NAND4_X1 port map( A1 => n37484, A2 => n37483, A3 => n37482, A4 => 
                           n37481, ZN => n37490);
   U2865 : AOI22_X1 port map( A1 => n31218, A2 => n29141, B1 => n31156, B2 => 
                           n29040, ZN => n37488);
   U2866 : AOI22_X1 port map( A1 => n31165, A2 => n29156, B1 => n31217, B2 => 
                           n29120, ZN => n37487);
   U2867 : AOI22_X1 port map( A1 => n31220, A2 => n29115, B1 => n31204, B2 => 
                           n29039, ZN => n37486);
   U2868 : AOI22_X1 port map( A1 => n30050, A2 => n29140, B1 => n31208, B2 => 
                           n29105, ZN => n37485);
   U2869 : NAND4_X1 port map( A1 => n37488, A2 => n37487, A3 => n37486, A4 => 
                           n37485, ZN => n37489);
   U2870 : AOI22_X1 port map( A1 => n37624, A2 => n37490, B1 => n37622, B2 => 
                           n37489, ZN => n37491);
   U2871 : OAI21_X1 port map( B1 => n37627, B2 => n37492, A => n37491, ZN => 
                           OUT2(6));
   U2872 : AOI22_X1 port map( A1 => n31222, A2 => n29734, B1 => n30082, B2 => 
                           n29752, ZN => n37496);
   U2873 : AOI22_X1 port map( A1 => n30084, A2 => n29071, B1 => n30078, B2 => 
                           n29060, ZN => n37495);
   U2874 : AOI22_X1 port map( A1 => n30070, A2 => n29073, B1 => n30077, B2 => 
                           n29057, ZN => n37494);
   U2875 : AOI22_X1 port map( A1 => n30079, A2 => n29723, B1 => n30072, B2 => 
                           n29052, ZN => n37493);
   U2876 : NAND4_X1 port map( A1 => n37496, A2 => n37495, A3 => n37494, A4 => 
                           n37493, ZN => n37502);
   U2877 : AOI22_X1 port map( A1 => n30073, A2 => n29732, B1 => n30080, B2 => 
                           n29061, ZN => n37500);
   U2878 : AOI22_X1 port map( A1 => n30083, A2 => n29737, B1 => n30076, B2 => 
                           n29046, ZN => n37499);
   U2879 : AOI22_X1 port map( A1 => n31228, A2 => n29058, B1 => n31206, B2 => 
                           n29068, ZN => n37498);
   U2880 : AOI22_X1 port map( A1 => n30081, A2 => n29751, B1 => n31200, B2 => 
                           n29069, ZN => n37497);
   U2881 : NAND4_X1 port map( A1 => n37500, A2 => n37499, A3 => n37498, A4 => 
                           n37497, ZN => n37501);
   U2882 : NOR2_X1 port map( A1 => n37502, A2 => n37501, ZN => n37514);
   U2883 : AOI22_X1 port map( A1 => n30050, A2 => n29814, B1 => n31208, B2 => 
                           n29827, ZN => n37506);
   U2884 : AOI22_X1 port map( A1 => n31219, A2 => n29809, B1 => n31218, B2 => 
                           n29806, ZN => n37505);
   U2885 : AOI22_X1 port map( A1 => n31204, A2 => n29826, B1 => n31202, B2 => 
                           n29817, ZN => n37504);
   U2886 : AOI22_X1 port map( A1 => n31220, A2 => n29825, B1 => n31217, B2 => 
                           n29824, ZN => n37503);
   U2887 : NAND4_X1 port map( A1 => n37506, A2 => n37505, A3 => n37504, A4 => 
                           n37503, ZN => n37512);
   U2888 : AOI22_X1 port map( A1 => n31219, A2 => n29138, B1 => n31216, B2 => 
                           n29121, ZN => n37510);
   U2889 : AOI22_X1 port map( A1 => n31218, A2 => n29151, B1 => n31208, B2 => 
                           n29109, ZN => n37509);
   U2890 : AOI22_X1 port map( A1 => n31220, A2 => n29110, B1 => n31209, B2 => 
                           n29137, ZN => n37508);
   U2891 : AOI22_X1 port map( A1 => n31156, A2 => n29063, B1 => n31204, B2 => 
                           n29065, ZN => n37507);
   U2892 : NAND4_X1 port map( A1 => n37510, A2 => n37509, A3 => n37508, A4 => 
                           n37507, ZN => n37511);
   U2893 : AOI22_X1 port map( A1 => n37624, A2 => n37512, B1 => n37622, B2 => 
                           n37511, ZN => n37513);
   U2894 : OAI21_X1 port map( B1 => n37627, B2 => n37514, A => n37513, ZN => 
                           OUT2(5));
   U2895 : AOI22_X1 port map( A1 => n31225, A2 => n29025, B1 => n31206, B2 => 
                           n29101, ZN => n37518);
   U2896 : AOI22_X1 port map( A1 => n30078, A2 => n29077, B1 => n30077, B2 => 
                           n29056, ZN => n37517);
   U2897 : AOI22_X1 port map( A1 => n31226, A2 => n29078, B1 => n31205, B2 => 
                           n29738, ZN => n37516);
   U2898 : AOI22_X1 port map( A1 => n30074, A2 => n29080, B1 => n30070, B2 => 
                           n29079, ZN => n37515);
   U2899 : NAND4_X1 port map( A1 => n37518, A2 => n37517, A3 => n37516, A4 => 
                           n37515, ZN => n37524);
   U2900 : AOI22_X1 port map( A1 => n31213, A2 => n29729, B1 => n30081, B2 => 
                           n29750, ZN => n37522);
   U2901 : AOI22_X1 port map( A1 => n30082, A2 => n29730, B1 => n30075, B2 => 
                           n29735, ZN => n37521);
   U2902 : AOI22_X1 port map( A1 => n30084, A2 => n29096, B1 => n31212, B2 => 
                           n29053, ZN => n37520);
   U2903 : AOI22_X1 port map( A1 => n30071, A2 => n29100, B1 => n31203, B2 => 
                           n29733, ZN => n37519);
   U2904 : NAND4_X1 port map( A1 => n37522, A2 => n37521, A3 => n37520, A4 => 
                           n37519, ZN => n37523);
   U2905 : NOR2_X1 port map( A1 => n37524, A2 => n37523, ZN => n37536);
   U2906 : AOI22_X1 port map( A1 => n31155, A2 => n29771, B1 => n31215, B2 => 
                           n29775, ZN => n37528);
   U2907 : AOI22_X1 port map( A1 => n31219, A2 => n29798, B1 => n31204, B2 => 
                           n29785, ZN => n37527);
   U2908 : AOI22_X1 port map( A1 => n31168, A2 => n29792, B1 => n31158, B2 => 
                           n29802, ZN => n37526);
   U2909 : AOI22_X1 port map( A1 => n31218, A2 => n29791, B1 => n31161, B2 => 
                           n29803, ZN => n37525);
   U2910 : NAND4_X1 port map( A1 => n37528, A2 => n37527, A3 => n37526, A4 => 
                           n37525, ZN => n37534);
   U2911 : AOI22_X1 port map( A1 => n31220, A2 => n29112, B1 => n31217, B2 => 
                           n29117, ZN => n37532);
   U2912 : AOI22_X1 port map( A1 => n31209, A2 => n29144, B1 => n31201, B2 => 
                           n29102, ZN => n37531);
   U2913 : AOI22_X1 port map( A1 => n31218, A2 => n29153, B1 => n31165, B2 => 
                           n29142, ZN => n37530);
   U2914 : AOI22_X1 port map( A1 => n31215, A2 => n29085, B1 => n31204, B2 => 
                           n29066, ZN => n37529);
   U2915 : NAND4_X1 port map( A1 => n37532, A2 => n37531, A3 => n37530, A4 => 
                           n37529, ZN => n37533);
   U2916 : AOI22_X1 port map( A1 => n37624, A2 => n37534, B1 => n37622, B2 => 
                           n37533, ZN => n37535);
   U2917 : OAI21_X1 port map( B1 => n37627, B2 => n37536, A => n37535, ZN => 
                           OUT2(4));
   U2918 : AOI22_X1 port map( A1 => n30079, A2 => n29727, B1 => n30081, B2 => 
                           n29749, ZN => n37540);
   U2919 : AOI22_X1 port map( A1 => n31225, A2 => n29027, B1 => n30074, B2 => 
                           n29082, ZN => n37539);
   U2920 : AOI22_X1 port map( A1 => n31227, A2 => n29055, B1 => n31200, B2 => 
                           n29092, ZN => n37538);
   U2921 : AOI22_X1 port map( A1 => n30073, A2 => n29755, B1 => n31212, B2 => 
                           n29059, ZN => n37537);
   U2922 : NAND4_X1 port map( A1 => n37540, A2 => n37539, A3 => n37538, A4 => 
                           n37537, ZN => n37546);
   U2923 : AOI22_X1 port map( A1 => n30069, A2 => n29094, B1 => n30083, B2 => 
                           n29740, ZN => n37544);
   U2924 : AOI22_X1 port map( A1 => n31226, A2 => n29089, B1 => n30070, B2 => 
                           n29081, ZN => n37543);
   U2925 : AOI22_X1 port map( A1 => n30084, A2 => n29091, B1 => n30078, B2 => 
                           n29088, ZN => n37542);
   U2926 : AOI22_X1 port map( A1 => n30082, A2 => n29724, B1 => n30075, B2 => 
                           n29721, ZN => n37541);
   U2927 : NAND4_X1 port map( A1 => n37544, A2 => n37543, A3 => n37542, A4 => 
                           n37541, ZN => n37545);
   U2928 : NOR2_X1 port map( A1 => n37546, A2 => n37545, ZN => n37558);
   U2929 : AOI22_X1 port map( A1 => n31208, A2 => n29794, B1 => n31217, B2 => 
                           n29808, ZN => n37550);
   U2930 : AOI22_X1 port map( A1 => n30050, A2 => n29807, B1 => n31204, B2 => 
                           n29793, ZN => n37549);
   U2931 : AOI22_X1 port map( A1 => n31165, A2 => n29787, B1 => n31202, B2 => 
                           n29796, ZN => n37548);
   U2932 : AOI22_X1 port map( A1 => n31218, A2 => n29804, B1 => n31220, B2 => 
                           n29795, ZN => n37547);
   U2933 : NAND4_X1 port map( A1 => n37550, A2 => n37549, A3 => n37548, A4 => 
                           n37547, ZN => n37556);
   U2934 : AOI22_X1 port map( A1 => n31158, A2 => n29106, B1 => n31165, B2 => 
                           n29154, ZN => n37554);
   U2935 : AOI22_X1 port map( A1 => n31209, A2 => n29147, B1 => n31204, B2 => 
                           n29067, ZN => n37553);
   U2936 : AOI22_X1 port map( A1 => n31155, A2 => n29125, B1 => n31215, B2 => 
                           n29076, ZN => n37552);
   U2937 : AOI22_X1 port map( A1 => n31220, A2 => n29104, B1 => n31157, B2 => 
                           n29158, ZN => n37551);
   U2938 : NAND4_X1 port map( A1 => n37554, A2 => n37553, A3 => n37552, A4 => 
                           n37551, ZN => n37555);
   U2939 : AOI22_X1 port map( A1 => n37624, A2 => n37556, B1 => n37622, B2 => 
                           n37555, ZN => n37557);
   U2940 : OAI21_X1 port map( B1 => n37627, B2 => n37558, A => n37557, ZN => 
                           OUT2(3));
   U2941 : AOI22_X1 port map( A1 => n30073, A2 => n29741, B1 => n31206, B2 => 
                           n29090, ZN => n37562);
   U2942 : AOI22_X1 port map( A1 => n31212, A2 => n29036, B1 => n30074, B2 => 
                           n29030, ZN => n37561);
   U2943 : AOI22_X1 port map( A1 => n30082, A2 => n29725, B1 => n30077, B2 => 
                           n29031, ZN => n37560);
   U2944 : AOI22_X1 port map( A1 => n31225, A2 => n29093, B1 => n30080, B2 => 
                           n29045, ZN => n37559);
   U2945 : NAND4_X1 port map( A1 => n37562, A2 => n37561, A3 => n37560, A4 => 
                           n37559, ZN => n37568);
   U2946 : AOI22_X1 port map( A1 => n30071, A2 => n29043, B1 => n31205, B2 => 
                           n29743, ZN => n37566);
   U2947 : AOI22_X1 port map( A1 => n30075, A2 => n29720, B1 => n31199, B2 => 
                           n29037, ZN => n37565);
   U2948 : AOI22_X1 port map( A1 => n30079, A2 => n29731, B1 => n30081, B2 => 
                           n29748, ZN => n37564);
   U2949 : AOI22_X1 port map( A1 => n30070, A2 => n29034, B1 => n31211, B2 => 
                           n29042, ZN => n37563);
   U2950 : NAND4_X1 port map( A1 => n37566, A2 => n37565, A3 => n37564, A4 => 
                           n37563, ZN => n37567);
   U2951 : NOR2_X1 port map( A1 => n37568, A2 => n37567, ZN => n37580);
   U2952 : AOI22_X1 port map( A1 => n31218, A2 => n29797, B1 => n31155, B2 => 
                           n29779, ZN => n37572);
   U2953 : AOI22_X1 port map( A1 => n31215, A2 => n29800, B1 => n31161, B2 => 
                           n29801, ZN => n37571);
   U2954 : AOI22_X1 port map( A1 => n31165, A2 => n29788, B1 => n31204, B2 => 
                           n29777, ZN => n37570);
   U2955 : AOI22_X1 port map( A1 => n30050, A2 => n29789, B1 => n31208, B2 => 
                           n29776, ZN => n37569);
   U2956 : NAND4_X1 port map( A1 => n37572, A2 => n37571, A3 => n37570, A4 => 
                           n37569, ZN => n37578);
   U2957 : AOI22_X1 port map( A1 => n31218, A2 => n29165, B1 => n31208, B2 => 
                           n29113, ZN => n37576);
   U2958 : AOI22_X1 port map( A1 => n31204, A2 => n29070, B1 => n31202, B2 => 
                           n29075, ZN => n37575);
   U2959 : AOI22_X1 port map( A1 => n31219, A2 => n29159, B1 => n31217, B2 => 
                           n29123, ZN => n37574);
   U2960 : AOI22_X1 port map( A1 => n31168, A2 => n29166, B1 => n31220, B2 => 
                           n29107, ZN => n37573);
   U2961 : NAND4_X1 port map( A1 => n37576, A2 => n37575, A3 => n37574, A4 => 
                           n37573, ZN => n37577);
   U2962 : AOI22_X1 port map( A1 => n37624, A2 => n37578, B1 => n37622, B2 => 
                           n37577, ZN => n37579);
   U2963 : OAI21_X1 port map( B1 => n37627, B2 => n37580, A => n37579, ZN => 
                           OUT2(2));
   U2964 : AOI22_X1 port map( A1 => n30080, A2 => n29062, B1 => n30081, B2 => 
                           n29746, ZN => n37584);
   U2965 : AOI22_X1 port map( A1 => n31222, A2 => n29739, B1 => n30070, B2 => 
                           n29083, ZN => n37583);
   U2966 : AOI22_X1 port map( A1 => n30069, A2 => n29098, B1 => n31207, B2 => 
                           n29747, ZN => n37582);
   U2967 : AOI22_X1 port map( A1 => n30073, A2 => n29742, B1 => n30071, B2 => 
                           n29097, ZN => n37581);
   U2968 : NAND4_X1 port map( A1 => n37584, A2 => n37583, A3 => n37582, A4 => 
                           n37581, ZN => n37590);
   U2969 : AOI22_X1 port map( A1 => n31227, A2 => n29032, B1 => n30076, B2 => 
                           n29099, ZN => n37588);
   U2970 : AOI22_X1 port map( A1 => n30079, A2 => n29722, B1 => n30074, B2 => 
                           n29084, ZN => n37587);
   U2971 : AOI22_X1 port map( A1 => n30072, A2 => n29064, B1 => n31199, B2 => 
                           n29087, ZN => n37586);
   U2972 : AOI22_X1 port map( A1 => n30084, A2 => n29095, B1 => n30083, B2 => 
                           n29753, ZN => n37585);
   U2973 : NAND4_X1 port map( A1 => n37588, A2 => n37587, A3 => n37586, A4 => 
                           n37585, ZN => n37589);
   U2974 : NOR2_X1 port map( A1 => n37590, A2 => n37589, ZN => n37602);
   U2975 : AOI22_X1 port map( A1 => n31162, A2 => n29783, B1 => n31161, B2 => 
                           n29790, ZN => n37594);
   U2976 : AOI22_X1 port map( A1 => n31219, A2 => n29767, B1 => n31218, B2 => 
                           n29780, ZN => n37593);
   U2977 : AOI22_X1 port map( A1 => n30050, A2 => n29781, B1 => n31215, B2 => 
                           n29773, ZN => n37592);
   U2978 : AOI22_X1 port map( A1 => n31158, A2 => n29786, B1 => n31217, B2 => 
                           n29782, ZN => n37591);
   U2979 : NAND4_X1 port map( A1 => n37594, A2 => n37593, A3 => n37592, A4 => 
                           n37591, ZN => n37600);
   U2980 : AOI22_X1 port map( A1 => n31220, A2 => n29108, B1 => n31202, B2 => 
                           n29074, ZN => n37598);
   U2981 : AOI22_X1 port map( A1 => n31158, A2 => n29103, B1 => n31162, B2 => 
                           n29072, ZN => n37597);
   U2982 : AOI22_X1 port map( A1 => n31218, A2 => n29143, B1 => n31217, B2 => 
                           n29116, ZN => n37596);
   U2983 : AOI22_X1 port map( A1 => n31168, A2 => n29139, B1 => n31165, B2 => 
                           n29149, ZN => n37595);
   U2984 : NAND4_X1 port map( A1 => n37598, A2 => n37597, A3 => n37596, A4 => 
                           n37595, ZN => n37599);
   U2985 : AOI22_X1 port map( A1 => n37624, A2 => n37600, B1 => n37622, B2 => 
                           n37599, ZN => n37601);
   U2986 : OAI21_X1 port map( B1 => n37627, B2 => n37602, A => n37601, ZN => 
                           OUT2(1));
   U2987 : AOI22_X1 port map( A1 => n30070, A2 => n29126, B1 => n30075, B2 => 
                           n29828, ZN => n37606);
   U2988 : AOI22_X1 port map( A1 => n31228, A2 => n29127, B1 => n30083, B2 => 
                           n29832, ZN => n37605);
   U2989 : AOI22_X1 port map( A1 => n31213, A2 => n29831, B1 => n30077, B2 => 
                           n29135, ZN => n37604);
   U2990 : AOI22_X1 port map( A1 => n30080, A2 => n29130, B1 => n31206, B2 => 
                           n29215, ZN => n37603);
   U2991 : NAND4_X1 port map( A1 => n37606, A2 => n37605, A3 => n37604, A4 => 
                           n37603, ZN => n37612);
   U2992 : AOI22_X1 port map( A1 => n30072, A2 => n29132, B1 => n31211, B2 => 
                           n29201, ZN => n37610);
   U2993 : AOI22_X1 port map( A1 => n31224, A2 => n29829, B1 => n31207, B2 => 
                           n29833, ZN => n37609);
   U2994 : AOI22_X1 port map( A1 => n30076, A2 => n29131, B1 => n31199, B2 => 
                           n29128, ZN => n37608);
   U2995 : AOI22_X1 port map( A1 => n30071, A2 => n29136, B1 => n31203, B2 => 
                           n29830, ZN => n37607);
   U2996 : NAND4_X1 port map( A1 => n37610, A2 => n37609, A3 => n37608, A4 => 
                           n37607, ZN => n37611);
   U2997 : NOR2_X1 port map( A1 => n37612, A2 => n37611, ZN => n37626);
   U2998 : AOI22_X1 port map( A1 => n31162, A2 => n29757, B1 => n31217, B2 => 
                           n29759, ZN => n37616);
   U2999 : AOI22_X1 port map( A1 => n31220, A2 => n29762, B1 => n31165, B2 => 
                           n29761, ZN => n37615);
   U3000 : AOI22_X1 port map( A1 => n31158, A2 => n29758, B1 => n31215, B2 => 
                           n29756, ZN => n37614);
   U3001 : AOI22_X1 port map( A1 => n31168, A2 => n29763, B1 => n31218, B2 => 
                           n29760, ZN => n37613);
   U3002 : NAND4_X1 port map( A1 => n37616, A2 => n37615, A3 => n37614, A4 => 
                           n37613, ZN => n37623);
   U3003 : AOI22_X1 port map( A1 => n31155, A2 => n29248, B1 => n31158, B2 => 
                           n29134, ZN => n37620);
   U3004 : AOI22_X1 port map( A1 => n31162, A2 => n29133, B1 => n31157, B2 => 
                           n29262, ZN => n37619);
   U3005 : AOI22_X1 port map( A1 => n31209, A2 => n29261, B1 => n31202, B2 => 
                           n29210, ZN => n37618);
   U3006 : AOI22_X1 port map( A1 => n31233, A2 => n29260, B1 => n31161, B2 => 
                           n29129, ZN => n37617);
   U3007 : NAND4_X1 port map( A1 => n37620, A2 => n37619, A3 => n37618, A4 => 
                           n37617, ZN => n37621);
   U3008 : AOI22_X1 port map( A1 => n37624, A2 => n37623, B1 => n37622, B2 => 
                           n37621, ZN => n37625);
   U3009 : OAI21_X1 port map( B1 => n37627, B2 => n37626, A => n37625, ZN => 
                           OUT2(0));
   U3010 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n37631)
                           ;
   U3011 : NOR2_X1 port map( A1 => n3566, A2 => n37631, ZN => n18308);
   U3012 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n3560, ZN => n37630);
   U3013 : INV_X1 port map( A => n3568, ZN => n37628);
   U3014 : NOR2_X1 port map( A1 => n37630, A2 => n37628, ZN => n18307);
   U3015 : NOR2_X1 port map( A1 => n3566, A2 => n37630, ZN => n18306);
   U3016 : NOR2_X1 port map( A1 => n37631, A2 => n3564, ZN => n18305);
   U3017 : NOR2_X1 port map( A1 => n37630, A2 => n3561, ZN => n18304);
   U3018 : NOR2_X1 port map( A1 => n37630, A2 => n3562, ZN => n18303);
   U3019 : NOR2_X1 port map( A1 => n37630, A2 => n3565, ZN => n18302);
   U3020 : NOR2_X1 port map( A1 => n37630, A2 => n3564, ZN => n18301);
   U3021 : NOR2_X1 port map( A1 => n37631, A2 => n37628, ZN => n18300);
   U3022 : NOR2_X1 port map( A1 => n37631, A2 => n3562, ZN => n18299);
   U3023 : INV_X1 port map( A => n3563, ZN => n37629);
   U3024 : NOR2_X1 port map( A1 => n37630, A2 => n37629, ZN => n18298);
   U3025 : NOR2_X1 port map( A1 => n37631, A2 => n37629, ZN => n18297);
   U3026 : NOR2_X1 port map( A1 => n37630, A2 => n3567, ZN => n18296);
   U3027 : NOR2_X1 port map( A1 => n37631, A2 => n3565, ZN => n18295);
   U3028 : NOR2_X1 port map( A1 => n37631, A2 => n3561, ZN => n18294);
   U3029 : NOR2_X1 port map( A1 => n37631, A2 => n3567, ZN => n18293);
   U3030 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n31273, A3 => n31271, ZN 
                           => n38342);
   U3031 : AOI22_X1 port map( A1 => n29372, A2 => n30067, B1 => n29880, B2 => 
                           n31198, ZN => n37635);
   U3032 : AOI22_X1 port map( A1 => n29369, A2 => n30066, B1 => n29900, B2 => 
                           n30060, ZN => n37634);
   U3033 : AOI22_X1 port map( A1 => n29375, A2 => n30063, B1 => n29370, B2 => 
                           n30056, ZN => n37633);
   U3034 : AOI22_X1 port map( A1 => n29309, A2 => n30061, B1 => n29914, B2 => 
                           n30057, ZN => n37632);
   U3035 : NAND4_X1 port map( A1 => n37635, A2 => n37634, A3 => n37633, A4 => 
                           n37632, ZN => n37641);
   U3036 : AOI22_X1 port map( A1 => n29891, A2 => n31197, B1 => n29377, B2 => 
                           n30053, ZN => n37639);
   U3037 : AOI22_X1 port map( A1 => n29376, A2 => n30068, B1 => n29373, B2 => 
                           n31195, ZN => n37638);
   U3038 : AOI22_X1 port map( A1 => n29371, A2 => n31196, B1 => n29895, B2 => 
                           n30055, ZN => n37637);
   U3039 : AOI22_X1 port map( A1 => n29374, A2 => n30058, B1 => n29872, B2 => 
                           n30065, ZN => n37636);
   U3040 : NAND4_X1 port map( A1 => n37639, A2 => n37638, A3 => n37637, A4 => 
                           n37636, ZN => n37640);
   U3041 : NOR2_X1 port map( A1 => n37641, A2 => n37640, ZN => n37653);
   U3042 : NOR3_X1 port map( A1 => n31268, A2 => n31269, A3 => n38295, ZN => 
                           n38172);
   U3043 : CLKBUF_X1 port map( A => n38172, Z => n38159);
   U3044 : AOI22_X1 port map( A1 => n30033, A2 => n31192, B1 => n30039, B2 => 
                           n31169, ZN => n37645);
   U3045 : AOI22_X1 port map( A1 => n30028, A2 => n30051, B1 => n30034, B2 => 
                           n30052, ZN => n37644);
   U3046 : AOI22_X1 port map( A1 => n30031, A2 => n31194, B1 => n30032, B2 => 
                           n31191, ZN => n37643);
   U3047 : AOI22_X1 port map( A1 => n30041, A2 => n31164, B1 => n30040, B2 => 
                           n31193, ZN => n37642);
   U3048 : NAND4_X1 port map( A1 => n37645, A2 => n37644, A3 => n37643, A4 => 
                           n37642, ZN => n37651);
   U3049 : NOR3_X1 port map( A1 => n31269, A2 => n30131, A3 => n38295, ZN => 
                           n37871);
   U3050 : AOI22_X1 port map( A1 => n29380, A2 => n31190, B1 => n29364, B2 => 
                           n30128, ZN => n37649);
   U3051 : AOI22_X1 port map( A1 => n29694, A2 => n31167, B1 => n29579, B2 => 
                           n30127, ZN => n37648);
   U3052 : AOI22_X1 port map( A1 => n29713, A2 => n31166, B1 => n29381, B2 => 
                           n31164, ZN => n37647);
   U3053 : AOI22_X1 port map( A1 => n29675, A2 => n31170, B1 => n29382, B2 => 
                           n31160, ZN => n37646);
   U3054 : NAND4_X1 port map( A1 => n37649, A2 => n37648, A3 => n37647, A4 => 
                           n37646, ZN => n37650);
   U3055 : AOI22_X1 port map( A1 => n38159, A2 => n37651, B1 => n37871, B2 => 
                           n37650, ZN => n37652);
   U3056 : OAI21_X1 port map( B1 => n38295, B2 => n37653, A => n37652, ZN => 
                           OUT1(31));
   U3057 : AOI22_X1 port map( A1 => n29206, A2 => n30068, B1 => n29424, B2 => 
                           n30058, ZN => n37657);
   U3058 : AOI22_X1 port map( A1 => n29422, A2 => n30062, B1 => n29421, B2 => 
                           n30056, ZN => n37656);
   U3059 : AOI22_X1 port map( A1 => n29423, A2 => n31195, B1 => n29194, B2 => 
                           n31189, ZN => n37655);
   U3060 : AOI22_X1 port map( A1 => n29599, A2 => n30059, B1 => n29418, B2 => 
                           n30066, ZN => n37654);
   U3061 : NAND4_X1 port map( A1 => n37657, A2 => n37656, A3 => n37655, A4 => 
                           n37654, ZN => n37663);
   U3062 : AOI22_X1 port map( A1 => n29426, A2 => n31188, B1 => n29611, B2 => 
                           n30060, ZN => n37661);
   U3063 : AOI22_X1 port map( A1 => n29627, A2 => n30055, B1 => n29419, B2 => 
                           n30053, ZN => n37660);
   U3064 : AOI22_X1 port map( A1 => n29209, A2 => n30065, B1 => n29640, B2 => 
                           n30054, ZN => n37659);
   U3065 : AOI22_X1 port map( A1 => n29308, A2 => n30061, B1 => n29604, B2 => 
                           n30057, ZN => n37658);
   U3066 : NAND4_X1 port map( A1 => n37661, A2 => n37660, A3 => n37659, A4 => 
                           n37658, ZN => n37662);
   U3067 : NOR2_X1 port map( A1 => n37663, A2 => n37662, ZN => n37675);
   U3068 : AOI22_X1 port map( A1 => n29205, A2 => n31171, B1 => n29636, B2 => 
                           n31186, ZN => n37667);
   U3069 : AOI22_X1 port map( A1 => n29202, A2 => n31191, B1 => n29203, B2 => 
                           n31187, ZN => n37666);
   U3070 : AOI22_X1 port map( A1 => n29204, A2 => n31159, B1 => n29615, B2 => 
                           n30126, ZN => n37665);
   U3071 : AOI22_X1 port map( A1 => n29179, A2 => n30052, B1 => n29199, B2 => 
                           n31169, ZN => n37664);
   U3072 : NAND4_X1 port map( A1 => n37667, A2 => n37666, A3 => n37665, A4 => 
                           n37664, ZN => n37673);
   U3073 : CLKBUF_X1 port map( A => n37871, Z => n38337);
   U3074 : AOI22_X1 port map( A1 => n29427, A2 => n31193, B1 => n29189, B2 => 
                           n31187, ZN => n37671);
   U3075 : AOI22_X1 port map( A1 => n29648, A2 => n31170, B1 => n29365, B2 => 
                           n31169, ZN => n37670);
   U3076 : AOI22_X1 port map( A1 => n29655, A2 => n31192, B1 => n29598, B2 => 
                           n31194, ZN => n37669);
   U3077 : AOI22_X1 port map( A1 => n29662, A2 => n31166, B1 => n29393, B2 => 
                           n31191, ZN => n37668);
   U3078 : NAND4_X1 port map( A1 => n37671, A2 => n37670, A3 => n37669, A4 => 
                           n37668, ZN => n37672);
   U3079 : AOI22_X1 port map( A1 => n38159, A2 => n37673, B1 => n38337, B2 => 
                           n37672, ZN => n37674);
   U3080 : OAI21_X1 port map( B1 => n38295, B2 => n37675, A => n37674, ZN => 
                           OUT1(30));
   U3081 : AOI22_X1 port map( A1 => n29400, A2 => n31184, B1 => n29412, B2 => 
                           n30064, ZN => n37679);
   U3082 : AOI22_X1 port map( A1 => n29414, A2 => n30063, B1 => n29409, B2 => 
                           n30056, ZN => n37678);
   U3083 : AOI22_X1 port map( A1 => n29984, A2 => n30060, B1 => n29413, B2 => 
                           n30058, ZN => n37677);
   U3084 : AOI22_X1 port map( A1 => n29957, A2 => n30057, B1 => n30010, B2 => 
                           n30059, ZN => n37676);
   U3085 : NAND4_X1 port map( A1 => n37679, A2 => n37678, A3 => n37677, A4 => 
                           n37676, ZN => n37685);
   U3086 : AOI22_X1 port map( A1 => n29410, A2 => n31196, B1 => n29401, B2 => 
                           n30053, ZN => n37683);
   U3087 : AOI22_X1 port map( A1 => n29411, A2 => n30067, B1 => n29944, B2 => 
                           n30054, ZN => n37682);
   U3088 : AOI22_X1 port map( A1 => n29307, A2 => n30061, B1 => n29407, B2 => 
                           n31183, ZN => n37681);
   U3089 : AOI22_X1 port map( A1 => n29889, A2 => n31185, B1 => n30022, B2 => 
                           n30055, ZN => n37680);
   U3090 : NAND4_X1 port map( A1 => n37683, A2 => n37682, A3 => n37681, A4 => 
                           n37680, ZN => n37684);
   U3091 : NOR2_X1 port map( A1 => n37685, A2 => n37684, ZN => n37697);
   U3092 : AOI22_X1 port map( A1 => n29911, A2 => n30052, B1 => n30036, B2 => 
                           n31167, ZN => n37689);
   U3093 : AOI22_X1 port map( A1 => n29912, A2 => n31171, B1 => n29915, B2 => 
                           n31164, ZN => n37688);
   U3094 : AOI22_X1 port map( A1 => n29913, A2 => n31193, B1 => n29916, B2 => 
                           n31160, ZN => n37687);
   U3095 : AOI22_X1 port map( A1 => n30035, A2 => n30051, B1 => n29917, B2 => 
                           n30128, ZN => n37686);
   U3096 : NAND4_X1 port map( A1 => n37689, A2 => n37688, A3 => n37687, A4 => 
                           n37686, ZN => n37695);
   U3097 : AOI22_X1 port map( A1 => n29707, A2 => n31166, B1 => n29595, B2 => 
                           n30127, ZN => n37693);
   U3098 : AOI22_X1 port map( A1 => n29392, A2 => n31160, B1 => n29406, B2 => 
                           n31187, ZN => n37692);
   U3099 : AOI22_X1 port map( A1 => n29696, A2 => n31192, B1 => n29281, B2 => 
                           n31159, ZN => n37691);
   U3100 : AOI22_X1 port map( A1 => n29706, A2 => n31182, B1 => n29366, B2 => 
                           n31169, ZN => n37690);
   U3101 : NAND4_X1 port map( A1 => n37693, A2 => n37692, A3 => n37691, A4 => 
                           n37690, ZN => n37694);
   U3102 : AOI22_X1 port map( A1 => n38159, A2 => n37695, B1 => n37871, B2 => 
                           n37694, ZN => n37696);
   U3103 : OAI21_X1 port map( B1 => n38295, B2 => n37697, A => n37696, ZN => 
                           OUT1(29));
   U3104 : AOI22_X1 port map( A1 => n29619, A2 => n31181, B1 => n29618, B2 => 
                           n30060, ZN => n37701);
   U3105 : AOI22_X1 port map( A1 => n29443, A2 => n30056, B1 => n29420, B2 => 
                           n30066, ZN => n37700);
   U3106 : AOI22_X1 port map( A1 => n29444, A2 => n30062, B1 => n29183, B2 => 
                           n30068, ZN => n37699);
   U3107 : AOI22_X1 port map( A1 => n29450, A2 => n30058, B1 => n29300, B2 => 
                           n30061, ZN => n37698);
   U3108 : NAND4_X1 port map( A1 => n37701, A2 => n37700, A3 => n37699, A4 => 
                           n37698, ZN => n37707);
   U3109 : AOI22_X1 port map( A1 => n29639, A2 => n31197, B1 => n29439, B2 => 
                           n30053, ZN => n37705);
   U3110 : AOI22_X1 port map( A1 => n29437, A2 => n30063, B1 => n29626, B2 => 
                           n30055, ZN => n37704);
   U3111 : AOI22_X1 port map( A1 => n29608, A2 => n31198, B1 => n29449, B2 => 
                           n31195, ZN => n37703);
   U3112 : AOI22_X1 port map( A1 => n29186, A2 => n30067, B1 => n29184, B2 => 
                           n30065, ZN => n37702);
   U3113 : NAND4_X1 port map( A1 => n37705, A2 => n37704, A3 => n37703, A4 => 
                           n37702, ZN => n37706);
   U3114 : NOR2_X1 port map( A1 => n37707, A2 => n37706, ZN => n37719);
   U3115 : AOI22_X1 port map( A1 => n29200, A2 => n30128, B1 => n29190, B2 => 
                           n30052, ZN => n37711);
   U3116 : AOI22_X1 port map( A1 => n29196, A2 => n31159, B1 => n29614, B2 => 
                           n31192, ZN => n37710);
   U3117 : AOI22_X1 port map( A1 => n29197, A2 => n30125, B1 => n29198, B2 => 
                           n31160, ZN => n37709);
   U3118 : AOI22_X1 port map( A1 => n29635, A2 => n31186, B1 => n29191, B2 => 
                           n31171, ZN => n37708);
   U3119 : NAND4_X1 port map( A1 => n37711, A2 => n37710, A3 => n37709, A4 => 
                           n37708, ZN => n37717);
   U3120 : AOI22_X1 port map( A1 => n29632, A2 => n31186, B1 => n29647, B2 => 
                           n31182, ZN => n37715);
   U3121 : AOI22_X1 port map( A1 => n29391, A2 => n31179, B1 => n29441, B2 => 
                           n31159, ZN => n37714);
   U3122 : AOI22_X1 port map( A1 => n29654, A2 => n30126, B1 => n29367, B2 => 
                           n31180, ZN => n37713);
   U3123 : AOI22_X1 port map( A1 => n29583, A2 => n31171, B1 => n29185, B2 => 
                           n31164, ZN => n37712);
   U3124 : NAND4_X1 port map( A1 => n37715, A2 => n37714, A3 => n37713, A4 => 
                           n37712, ZN => n37716);
   U3125 : AOI22_X1 port map( A1 => n38159, A2 => n37717, B1 => n38337, B2 => 
                           n37716, ZN => n37718);
   U3126 : OAI21_X1 port map( B1 => n38295, B2 => n37719, A => n37718, ZN => 
                           OUT1(28));
   U3127 : AOI22_X1 port map( A1 => n29431, A2 => n30053, B1 => n29188, B2 => 
                           n31184, ZN => n37723);
   U3128 : AOI22_X1 port map( A1 => n29433, A2 => n30066, B1 => n29193, B2 => 
                           n31189, ZN => n37722);
   U3129 : AOI22_X1 port map( A1 => n29435, A2 => n31196, B1 => n29625, B2 => 
                           n30055, ZN => n37721);
   U3130 : AOI22_X1 port map( A1 => n29429, A2 => n31177, B1 => n29434, B2 => 
                           n30056, ZN => n37720);
   U3131 : NAND4_X1 port map( A1 => n37723, A2 => n37722, A3 => n37721, A4 => 
                           n37720, ZN => n37729);
   U3132 : AOI22_X1 port map( A1 => n29187, A2 => n31185, B1 => n29430, B2 => 
                           n30063, ZN => n37727);
   U3133 : AOI22_X1 port map( A1 => n29606, A2 => n31176, B1 => n29617, B2 => 
                           n30059, ZN => n37726);
   U3134 : AOI22_X1 port map( A1 => n29299, A2 => n31178, B1 => n29436, B2 => 
                           n30064, ZN => n37725);
   U3135 : AOI22_X1 port map( A1 => n29638, A2 => n31197, B1 => n29623, B2 => 
                           n30057, ZN => n37724);
   U3136 : NAND4_X1 port map( A1 => n37727, A2 => n37726, A3 => n37725, A4 => 
                           n37724, ZN => n37728);
   U3137 : NOR2_X1 port map( A1 => n37729, A2 => n37728, ZN => n37741);
   U3138 : AOI22_X1 port map( A1 => n29180, A2 => n31191, B1 => n29182, B2 => 
                           n30128, ZN => n37733);
   U3139 : AOI22_X1 port map( A1 => n29631, A2 => n31167, B1 => n29175, B2 => 
                           n30052, ZN => n37732);
   U3140 : AOI22_X1 port map( A1 => n29177, A2 => n31159, B1 => n29167, B2 => 
                           n31194, ZN => n37731);
   U3141 : AOI22_X1 port map( A1 => n29178, A2 => n31187, B1 => n29634, B2 => 
                           n31166, ZN => n37730);
   U3142 : NAND4_X1 port map( A1 => n37733, A2 => n37732, A3 => n37731, A4 => 
                           n37730, ZN => n37739);
   U3143 : AOI22_X1 port map( A1 => n29646, A2 => n31170, B1 => n29432, B2 => 
                           n31190, ZN => n37737);
   U3144 : AOI22_X1 port map( A1 => n29368, A2 => n31180, B1 => n29661, B2 => 
                           n30051, ZN => n37736);
   U3145 : AOI22_X1 port map( A1 => n29597, A2 => n31194, B1 => n29390, B2 => 
                           n31160, ZN => n37735);
   U3146 : AOI22_X1 port map( A1 => n29181, A2 => n31164, B1 => n29653, B2 => 
                           n31167, ZN => n37734);
   U3147 : NAND4_X1 port map( A1 => n37737, A2 => n37736, A3 => n37735, A4 => 
                           n37734, ZN => n37738);
   U3148 : AOI22_X1 port map( A1 => n38159, A2 => n37739, B1 => n37871, B2 => 
                           n37738, ZN => n37740);
   U3149 : OAI21_X1 port map( B1 => n38295, B2 => n37741, A => n37740, ZN => 
                           OUT1(27));
   U3150 : AOI22_X1 port map( A1 => n29453, A2 => n30066, B1 => n29469, B2 => 
                           n31175, ZN => n37745);
   U3151 : AOI22_X1 port map( A1 => n29468, A2 => n30068, B1 => n29964, B2 => 
                           n30054, ZN => n37744);
   U3152 : AOI22_X1 port map( A1 => n29890, A2 => n31185, B1 => n29945, B2 => 
                           n31181, ZN => n37743);
   U3153 : AOI22_X1 port map( A1 => n30023, A2 => n31174, B1 => n29465, B2 => 
                           n30064, ZN => n37742);
   U3154 : NAND4_X1 port map( A1 => n37745, A2 => n37744, A3 => n37743, A4 => 
                           n37742, ZN => n37751);
   U3155 : AOI22_X1 port map( A1 => n29983, A2 => n30060, B1 => n29467, B2 => 
                           n30063, ZN => n37749);
   U3156 : AOI22_X1 port map( A1 => n30017, A2 => n31198, B1 => n29298, B2 => 
                           n30061, ZN => n37748);
   U3157 : AOI22_X1 port map( A1 => n29464, A2 => n30067, B1 => n29463, B2 => 
                           n30062, ZN => n37747);
   U3158 : AOI22_X1 port map( A1 => n29461, A2 => n30056, B1 => n29466, B2 => 
                           n30058, ZN => n37746);
   U3159 : NAND4_X1 port map( A1 => n37749, A2 => n37748, A3 => n37747, A4 => 
                           n37746, ZN => n37750);
   U3160 : NOR2_X1 port map( A1 => n37751, A2 => n37750, ZN => n37763);
   U3161 : AOI22_X1 port map( A1 => n29899, A2 => n31182, B1 => n29910, B2 => 
                           n31179, ZN => n37755);
   U3162 : AOI22_X1 port map( A1 => n29898, A2 => n31194, B1 => n29909, B2 => 
                           n31180, ZN => n37754);
   U3163 : AOI22_X1 port map( A1 => n30037, A2 => n31186, B1 => n30029, B2 => 
                           n31192, ZN => n37753);
   U3164 : AOI22_X1 port map( A1 => n29896, A2 => n31187, B1 => n29897, B2 => 
                           n31193, ZN => n37752);
   U3165 : NAND4_X1 port map( A1 => n37755, A2 => n37754, A3 => n37753, A4 => 
                           n37752, ZN => n37761);
   U3166 : AOI22_X1 port map( A1 => n29704, A2 => n31186, B1 => n29378, B2 => 
                           n31169, ZN => n37759);
   U3167 : AOI22_X1 port map( A1 => n29681, A2 => n31192, B1 => n29389, B2 => 
                           n31160, ZN => n37758);
   U3168 : AOI22_X1 port map( A1 => n29587, A2 => n30127, B1 => n29428, B2 => 
                           n30125, ZN => n37757);
   U3169 : AOI22_X1 port map( A1 => n29682, A2 => n30052, B1 => n29472, B2 => 
                           n31193, ZN => n37756);
   U3170 : NAND4_X1 port map( A1 => n37759, A2 => n37758, A3 => n37757, A4 => 
                           n37756, ZN => n37760);
   U3171 : AOI22_X1 port map( A1 => n38159, A2 => n37761, B1 => n38337, B2 => 
                           n37760, ZN => n37762);
   U3172 : OAI21_X1 port map( B1 => n38295, B2 => n37763, A => n37762, ZN => 
                           OUT1(26));
   U3173 : AOI22_X1 port map( A1 => n29169, A2 => n30067, B1 => n29481, B2 => 
                           n31177, ZN => n37767);
   U3174 : AOI22_X1 port map( A1 => n29353, A2 => n31173, B1 => n29600, B2 => 
                           n31198, ZN => n37766);
   U3175 : AOI22_X1 port map( A1 => n29297, A2 => n30061, B1 => n29480, B2 => 
                           n30064, ZN => n37765);
   U3176 : AOI22_X1 port map( A1 => n29170, A2 => n30068, B1 => n29171, B2 => 
                           n30065, ZN => n37764);
   U3177 : NAND4_X1 port map( A1 => n37767, A2 => n37766, A3 => n37765, A4 => 
                           n37764, ZN => n37773);
   U3178 : AOI22_X1 port map( A1 => n29624, A2 => n31174, B1 => n29482, B2 => 
                           n31188, ZN => n37771);
   U3179 : AOI22_X1 port map( A1 => n29605, A2 => n31176, B1 => n29351, B2 => 
                           n30062, ZN => n37770);
   U3180 : AOI22_X1 port map( A1 => n29637, A2 => n30054, B1 => n29622, B2 => 
                           n30057, ZN => n37769);
   U3181 : AOI22_X1 port map( A1 => n29352, A2 => n31183, B1 => n29483, B2 => 
                           n31175, ZN => n37768);
   U3182 : NAND4_X1 port map( A1 => n37771, A2 => n37770, A3 => n37769, A4 => 
                           n37768, ZN => n37772);
   U3183 : NOR2_X1 port map( A1 => n37773, A2 => n37772, ZN => n37785);
   U3184 : AOI22_X1 port map( A1 => n29633, A2 => n31166, B1 => n29213, B2 => 
                           n30127, ZN => n37777);
   U3185 : AOI22_X1 port map( A1 => n29168, A2 => n31160, B1 => n29612, B2 => 
                           n31167, ZN => n37776);
   U3186 : AOI22_X1 port map( A1 => n29176, A2 => n31190, B1 => n29174, B2 => 
                           n31164, ZN => n37775);
   U3187 : AOI22_X1 port map( A1 => n29173, A2 => n30128, B1 => n29223, B2 => 
                           n31182, ZN => n37774);
   U3188 : NAND4_X1 port map( A1 => n37777, A2 => n37776, A3 => n37775, A4 => 
                           n37774, ZN => n37783);
   U3189 : AOI22_X1 port map( A1 => n29659, A2 => n30051, B1 => n29425, B2 => 
                           n31190, ZN => n37781);
   U3190 : AOI22_X1 port map( A1 => n29652, A2 => n30126, B1 => n29278, B2 => 
                           n31179, ZN => n37780);
   U3191 : AOI22_X1 port map( A1 => n29192, A2 => n31187, B1 => n29594, B2 => 
                           n31194, ZN => n37779);
   U3192 : AOI22_X1 port map( A1 => n29330, A2 => n31169, B1 => n29645, B2 => 
                           n30052, ZN => n37778);
   U3193 : NAND4_X1 port map( A1 => n37781, A2 => n37780, A3 => n37779, A4 => 
                           n37778, ZN => n37782);
   U3194 : AOI22_X1 port map( A1 => n38159, A2 => n37783, B1 => n38337, B2 => 
                           n37782, ZN => n37784);
   U3195 : OAI21_X1 port map( B1 => n38295, B2 => n37785, A => n37784, ZN => 
                           OUT1(25));
   U3196 : AOI22_X1 port map( A1 => n29930, A2 => n31185, B1 => n29301, B2 => 
                           n30053, ZN => n37789);
   U3197 : AOI22_X1 port map( A1 => n29283, A2 => n31173, B1 => n29960, B2 => 
                           n31181, ZN => n37788);
   U3198 : AOI22_X1 port map( A1 => n29302, A2 => n30068, B1 => n30018, B2 => 
                           n31198, ZN => n37787);
   U3199 : AOI22_X1 port map( A1 => n29305, A2 => n31195, B1 => n29306, B2 => 
                           n30062, ZN => n37786);
   U3200 : NAND4_X1 port map( A1 => n37789, A2 => n37788, A3 => n37787, A4 => 
                           n37786, ZN => n37795);
   U3201 : AOI22_X1 port map( A1 => n29303, A2 => n30063, B1 => n29982, B2 => 
                           n30060, ZN => n37793);
   U3202 : AOI22_X1 port map( A1 => n29304, A2 => n31177, B1 => n30025, B2 => 
                           n30055, ZN => n37792);
   U3203 : AOI22_X1 port map( A1 => n29952, A2 => n30054, B1 => n29284, B2 => 
                           n30066, ZN => n37791);
   U3204 : AOI22_X1 port map( A1 => n29276, A2 => n31178, B1 => n29554, B2 => 
                           n31189, ZN => n37790);
   U3205 : NAND4_X1 port map( A1 => n37793, A2 => n37792, A3 => n37791, A4 => 
                           n37790, ZN => n37794);
   U3206 : NOR2_X1 port map( A1 => n37795, A2 => n37794, ZN => n37807);
   U3207 : AOI22_X1 port map( A1 => n29928, A2 => n31182, B1 => n29932, B2 => 
                           n31191, ZN => n37799);
   U3208 : AOI22_X1 port map( A1 => n29926, A2 => n31190, B1 => n30030, B2 => 
                           n31186, ZN => n37798);
   U3209 : AOI22_X1 port map( A1 => n29929, A2 => n31171, B1 => n30038, B2 => 
                           n30126, ZN => n37797);
   U3210 : AOI22_X1 port map( A1 => n29927, A2 => n31169, B1 => n29931, B2 => 
                           n31164, ZN => n37796);
   U3211 : NAND4_X1 port map( A1 => n37799, A2 => n37798, A3 => n37797, A4 => 
                           n37796, ZN => n37805);
   U3212 : AOI22_X1 port map( A1 => n29287, A2 => n31191, B1 => n29296, B2 => 
                           n31159, ZN => n37803);
   U3213 : AOI22_X1 port map( A1 => n29712, A2 => n31192, B1 => n29684, B2 => 
                           n31170, ZN => n37802);
   U3214 : AOI22_X1 port map( A1 => n29288, A2 => n31187, B1 => n29286, B2 => 
                           n31180, ZN => n37801);
   U3215 : AOI22_X1 port map( A1 => n29588, A2 => n30127, B1 => n29692, B2 => 
                           n31186, ZN => n37800);
   U3216 : NAND4_X1 port map( A1 => n37803, A2 => n37802, A3 => n37801, A4 => 
                           n37800, ZN => n37804);
   U3217 : AOI22_X1 port map( A1 => n38159, A2 => n37805, B1 => n37871, B2 => 
                           n37804, ZN => n37806);
   U3218 : OAI21_X1 port map( B1 => n38295, B2 => n37807, A => n37806, ZN => 
                           OUT1(24));
   U3219 : AOI22_X1 port map( A1 => n29569, A2 => n30064, B1 => n29555, B2 => 
                           n30053, ZN => n37811);
   U3220 : AOI22_X1 port map( A1 => n29548, A2 => n30068, B1 => n29609, B2 => 
                           n31198, ZN => n37810);
   U3221 : AOI22_X1 port map( A1 => n29621, A2 => n31181, B1 => n29660, B2 => 
                           n31174, ZN => n37809);
   U3222 : AOI22_X1 port map( A1 => n29275, A2 => n30061, B1 => n29514, B2 => 
                           n30058, ZN => n37808);
   U3223 : NAND4_X1 port map( A1 => n37811, A2 => n37810, A3 => n37809, A4 => 
                           n37808, ZN => n37817);
   U3224 : AOI22_X1 port map( A1 => n29536, A2 => n31188, B1 => n29607, B2 => 
                           n30054, ZN => n37815);
   U3225 : AOI22_X1 port map( A1 => n29344, A2 => n30056, B1 => n29567, B2 => 
                           n31196, ZN => n37814);
   U3226 : AOI22_X1 port map( A1 => n29649, A2 => n30065, B1 => n29610, B2 => 
                           n30060, ZN => n37813);
   U3227 : AOI22_X1 port map( A1 => n29457, A2 => n31183, B1 => n29568, B2 => 
                           n30067, ZN => n37812);
   U3228 : NAND4_X1 port map( A1 => n37815, A2 => n37814, A3 => n37813, A4 => 
                           n37812, ZN => n37816);
   U3229 : NOR2_X1 port map( A1 => n37817, A2 => n37816, ZN => n37829);
   U3230 : AOI22_X1 port map( A1 => n29195, A2 => n31194, B1 => n29225, B2 => 
                           n31190, ZN => n37821);
   U3231 : AOI22_X1 port map( A1 => n29212, A2 => n30051, B1 => n29231, B2 => 
                           n30128, ZN => n37820);
   U3232 : AOI22_X1 port map( A1 => n29226, A2 => n30125, B1 => n29208, B2 => 
                           n30126, ZN => n37819);
   U3233 : AOI22_X1 port map( A1 => n29207, A2 => n30052, B1 => n29228, B2 => 
                           n31160, ZN => n37818);
   U3234 : NAND4_X1 port map( A1 => n37821, A2 => n37820, A3 => n37819, A4 => 
                           n37818, ZN => n37827);
   U3235 : AOI22_X1 port map( A1 => n29581, A2 => n30127, B1 => n29221, B2 => 
                           n31160, ZN => n37825);
   U3236 : AOI22_X1 port map( A1 => n29230, A2 => n31164, B1 => n29379, B2 => 
                           n31180, ZN => n37824);
   U3237 : AOI22_X1 port map( A1 => n29462, A2 => n31159, B1 => n29657, B2 => 
                           n30051, ZN => n37823);
   U3238 : AOI22_X1 port map( A1 => n29651, A2 => n30126, B1 => n29644, B2 => 
                           n31182, ZN => n37822);
   U3239 : NAND4_X1 port map( A1 => n37825, A2 => n37824, A3 => n37823, A4 => 
                           n37822, ZN => n37826);
   U3240 : AOI22_X1 port map( A1 => n38159, A2 => n37827, B1 => n37871, B2 => 
                           n37826, ZN => n37828);
   U3241 : OAI21_X1 port map( B1 => n38342, B2 => n37829, A => n37828, ZN => 
                           OUT1(23));
   U3242 : AOI22_X1 port map( A1 => n29566, A2 => n30067, B1 => n29620, B2 => 
                           n30057, ZN => n37833);
   U3243 : AOI22_X1 port map( A1 => n29458, A2 => n31183, B1 => n29537, B2 => 
                           n31188, ZN => n37832);
   U3244 : AOI22_X1 port map( A1 => n29343, A2 => n30056, B1 => n29507, B2 => 
                           n30058, ZN => n37831);
   U3245 : AOI22_X1 port map( A1 => n29549, A2 => n31184, B1 => n29629, B2 => 
                           n31197, ZN => n37830);
   U3246 : NAND4_X1 port map( A1 => n37833, A2 => n37832, A3 => n37831, A4 => 
                           n37830, ZN => n37839);
   U3247 : AOI22_X1 port map( A1 => n29565, A2 => n31196, B1 => n29613, B2 => 
                           n31198, ZN => n37837);
   U3248 : AOI22_X1 port map( A1 => n29274, A2 => n31178, B1 => n29642, B2 => 
                           n30060, ZN => n37836);
   U3249 : AOI22_X1 port map( A1 => n29630, A2 => n30065, B1 => n29564, B2 => 
                           n31195, ZN => n37835);
   U3250 : AOI22_X1 port map( A1 => n29556, A2 => n30053, B1 => n29658, B2 => 
                           n30055, ZN => n37834);
   U3251 : NAND4_X1 port map( A1 => n37837, A2 => n37836, A3 => n37835, A4 => 
                           n37834, ZN => n37838);
   U3252 : NOR2_X1 port map( A1 => n37839, A2 => n37838, ZN => n37851);
   U3253 : AOI22_X1 port map( A1 => n29222, A2 => n31159, B1 => n29227, B2 => 
                           n31179, ZN => n37843);
   U3254 : AOI22_X1 port map( A1 => n29224, A2 => n31187, B1 => n29220, B2 => 
                           n31171, ZN => n37842);
   U3255 : AOI22_X1 port map( A1 => n29217, A2 => n31166, B1 => n29219, B2 => 
                           n30052, ZN => n37841);
   U3256 : AOI22_X1 port map( A1 => n29218, A2 => n31167, B1 => n29229, B2 => 
                           n31169, ZN => n37840);
   U3257 : NAND4_X1 port map( A1 => n37843, A2 => n37842, A3 => n37841, A4 => 
                           n37840, ZN => n37849);
   U3258 : AOI22_X1 port map( A1 => n29456, A2 => n31159, B1 => n29650, B2 => 
                           n30126, ZN => n37847);
   U3259 : AOI22_X1 port map( A1 => n29643, A2 => n30052, B1 => n29656, B2 => 
                           n30051, ZN => n37846);
   U3260 : AOI22_X1 port map( A1 => n29589, A2 => n31171, B1 => n29216, B2 => 
                           n31160, ZN => n37845);
   U3261 : AOI22_X1 port map( A1 => n29214, A2 => n31164, B1 => n29383, B2 => 
                           n31169, ZN => n37844);
   U3262 : NAND4_X1 port map( A1 => n37847, A2 => n37846, A3 => n37845, A4 => 
                           n37844, ZN => n37848);
   U3263 : AOI22_X1 port map( A1 => n38159, A2 => n37849, B1 => n37871, B2 => 
                           n37848, ZN => n37850);
   U3264 : OAI21_X1 port map( B1 => n38342, B2 => n37851, A => n37850, ZN => 
                           OUT1(22));
   U3265 : AOI22_X1 port map( A1 => n29348, A2 => n31177, B1 => n29346, B2 => 
                           n31184, ZN => n37855);
   U3266 : AOI22_X1 port map( A1 => n29336, A2 => n30066, B1 => n29334, B2 => 
                           n30062, ZN => n37854);
   U3267 : AOI22_X1 port map( A1 => n29350, A2 => n31189, B1 => n29345, B2 => 
                           n30053, ZN => n37853);
   U3268 : AOI22_X1 port map( A1 => n29347, A2 => n30063, B1 => n29981, B2 => 
                           n31176, ZN => n37852);
   U3269 : NAND4_X1 port map( A1 => n37855, A2 => n37854, A3 => n37853, A4 => 
                           n37852, ZN => n37861);
   U3270 : AOI22_X1 port map( A1 => n29999, A2 => n30065, B1 => n29335, B2 => 
                           n30056, ZN => n37859);
   U3271 : AOI22_X1 port map( A1 => n29966, A2 => n30057, B1 => n30019, B2 => 
                           n30059, ZN => n37858);
   U3272 : AOI22_X1 port map( A1 => n29349, A2 => n30064, B1 => n29946, B2 => 
                           n31197, ZN => n37857);
   U3273 : AOI22_X1 port map( A1 => n29273, A2 => n30061, B1 => n29988, B2 => 
                           n31174, ZN => n37856);
   U3274 : NAND4_X1 port map( A1 => n37859, A2 => n37858, A3 => n37857, A4 => 
                           n37856, ZN => n37860);
   U3275 : NOR2_X1 port map( A1 => n37861, A2 => n37860, ZN => n37874);
   U3276 : AOI22_X1 port map( A1 => n29850, A2 => n30127, B1 => n29847, B2 => 
                           n31160, ZN => n37865);
   U3277 : AOI22_X1 port map( A1 => n29852, A2 => n31170, B1 => n29853, B2 => 
                           n31167, ZN => n37864);
   U3278 : AOI22_X1 port map( A1 => n29855, A2 => n31186, B1 => n29848, B2 => 
                           n31164, ZN => n37863);
   U3279 : AOI22_X1 port map( A1 => n29849, A2 => n31190, B1 => n29846, B2 => 
                           n30128, ZN => n37862);
   U3280 : NAND4_X1 port map( A1 => n37865, A2 => n37864, A3 => n37863, A4 => 
                           n37862, ZN => n37872);
   U3281 : AOI22_X1 port map( A1 => n29338, A2 => n31160, B1 => n29687, B2 => 
                           n30052, ZN => n37869);
   U3282 : AOI22_X1 port map( A1 => n29340, A2 => n31190, B1 => n29591, B2 => 
                           n30127, ZN => n37868);
   U3283 : AOI22_X1 port map( A1 => n29671, A2 => n31192, B1 => n29698, B2 => 
                           n30051, ZN => n37867);
   U3284 : AOI22_X1 port map( A1 => n29337, A2 => n30128, B1 => n29339, B2 => 
                           n31164, ZN => n37866);
   U3285 : NAND4_X1 port map( A1 => n37869, A2 => n37868, A3 => n37867, A4 => 
                           n37866, ZN => n37870);
   U3286 : AOI22_X1 port map( A1 => n38159, A2 => n37872, B1 => n37871, B2 => 
                           n37870, ZN => n37873);
   U3287 : OAI21_X1 port map( B1 => n38342, B2 => n37874, A => n37873, ZN => 
                           OUT1(21));
   U3288 : AOI22_X1 port map( A1 => n29616, A2 => n30055, B1 => n29506, B2 => 
                           n31177, ZN => n37878);
   U3289 : AOI22_X1 port map( A1 => n29603, A2 => n30059, B1 => n29570, B2 => 
                           n31196, ZN => n37877);
   U3290 : AOI22_X1 port map( A1 => n29459, A2 => n31183, B1 => n29342, B2 => 
                           n31173, ZN => n37876);
   U3291 : AOI22_X1 port map( A1 => n29557, A2 => n30053, B1 => n29575, B2 => 
                           n30067, ZN => n37875);
   U3292 : NAND4_X1 port map( A1 => n37878, A2 => n37877, A3 => n37876, A4 => 
                           n37875, ZN => n37884);
   U3293 : AOI22_X1 port map( A1 => n29628, A2 => n31185, B1 => n29538, B2 => 
                           n30063, ZN => n37882);
   U3294 : AOI22_X1 port map( A1 => n29602, A2 => n31181, B1 => n29601, B2 => 
                           n30054, ZN => n37881);
   U3295 : AOI22_X1 port map( A1 => n29576, A2 => n30064, B1 => n29272, B2 => 
                           n30061, ZN => n37880);
   U3296 : AOI22_X1 port map( A1 => n29641, A2 => n31176, B1 => n29550, B2 => 
                           n31184, ZN => n37879);
   U3297 : NAND4_X1 port map( A1 => n37882, A2 => n37881, A3 => n37880, A4 => 
                           n37879, ZN => n37883);
   U3298 : NOR2_X1 port map( A1 => n37884, A2 => n37883, ZN => n37896);
   U3299 : AOI22_X1 port map( A1 => n29232, A2 => n31170, B1 => n29241, B2 => 
                           n31169, ZN => n37888);
   U3300 : AOI22_X1 port map( A1 => n29240, A2 => n31167, B1 => n29243, B2 => 
                           n31190, ZN => n37887);
   U3301 : AOI22_X1 port map( A1 => n29238, A2 => n31187, B1 => n29242, B2 => 
                           n31191, ZN => n37886);
   U3302 : AOI22_X1 port map( A1 => n29234, A2 => n31166, B1 => n29235, B2 => 
                           n31171, ZN => n37885);
   U3303 : NAND4_X1 port map( A1 => n37888, A2 => n37887, A3 => n37886, A4 => 
                           n37885, ZN => n37894);
   U3304 : AOI22_X1 port map( A1 => n29161, A2 => n31170, B1 => n29211, B2 => 
                           n31187, ZN => n37892);
   U3305 : AOI22_X1 port map( A1 => n29157, A2 => n31186, B1 => n29172, B2 => 
                           n31160, ZN => n37891);
   U3306 : AOI22_X1 port map( A1 => n29164, A2 => n31192, B1 => n29455, B2 => 
                           n31190, ZN => n37890);
   U3307 : AOI22_X1 port map( A1 => n29384, A2 => n31169, B1 => n29119, B2 => 
                           n31194, ZN => n37889);
   U3308 : NAND4_X1 port map( A1 => n37892, A2 => n37891, A3 => n37890, A4 => 
                           n37889, ZN => n37893);
   U3309 : AOI22_X1 port map( A1 => n38159, A2 => n37894, B1 => n38337, B2 => 
                           n37893, ZN => n37895);
   U3310 : OAI21_X1 port map( B1 => n38342, B2 => n37896, A => n37895, ZN => 
                           OUT1(20));
   U3311 : AOI22_X1 port map( A1 => n29953, A2 => n30054, B1 => n29505, B2 => 
                           n30058, ZN => n37900);
   U3312 : AOI22_X1 port map( A1 => n29558, A2 => n31175, B1 => n29539, B2 => 
                           n30063, ZN => n37899);
   U3313 : AOI22_X1 port map( A1 => n29972, A2 => n30057, B1 => n29571, B2 => 
                           n31196, ZN => n37898);
   U3314 : AOI22_X1 port map( A1 => n30021, A2 => n30059, B1 => n29341, B2 => 
                           n31173, ZN => n37897);
   U3315 : NAND4_X1 port map( A1 => n37900, A2 => n37899, A3 => n37898, A4 => 
                           n37897, ZN => n37906);
   U3316 : AOI22_X1 port map( A1 => n29551, A2 => n30068, B1 => n29980, B2 => 
                           n30060, ZN => n37904);
   U3317 : AOI22_X1 port map( A1 => n30003, A2 => n31185, B1 => n29271, B2 => 
                           n30061, ZN => n37903);
   U3318 : AOI22_X1 port map( A1 => n29573, A2 => n30064, B1 => n29991, B2 => 
                           n30055, ZN => n37902);
   U3319 : AOI22_X1 port map( A1 => n29572, A2 => n31189, B1 => n29460, B2 => 
                           n30066, ZN => n37901);
   U3320 : NAND4_X1 port map( A1 => n37904, A2 => n37903, A3 => n37902, A4 => 
                           n37901, ZN => n37905);
   U3321 : NOR2_X1 port map( A1 => n37906, A2 => n37905, ZN => n37918);
   U3322 : AOI22_X1 port map( A1 => n29834, A2 => n31160, B1 => n29854, B2 => 
                           n31192, ZN => n37910);
   U3323 : AOI22_X1 port map( A1 => n29835, A2 => n31187, B1 => n29837, B2 => 
                           n30127, ZN => n37909);
   U3324 : AOI22_X1 port map( A1 => n29838, A2 => n31182, B1 => n29836, B2 => 
                           n31180, ZN => n37908);
   U3325 : AOI22_X1 port map( A1 => n29851, A2 => n31190, B1 => n29866, B2 => 
                           n31166, ZN => n37907);
   U3326 : NAND4_X1 port map( A1 => n37910, A2 => n37909, A3 => n37908, A4 => 
                           n37907, ZN => n37916);
   U3327 : AOI22_X1 port map( A1 => n29688, A2 => n31170, B1 => n29454, B2 => 
                           n31193, ZN => n37914);
   U3328 : AOI22_X1 port map( A1 => n29596, A2 => n31171, B1 => n29690, B2 => 
                           n30051, ZN => n37913);
   U3329 : AOI22_X1 port map( A1 => n29685, A2 => n31167, B1 => n29417, B2 => 
                           n31164, ZN => n37912);
   U3330 : AOI22_X1 port map( A1 => n29385, A2 => n31169, B1 => n29363, B2 => 
                           n31191, ZN => n37911);
   U3331 : NAND4_X1 port map( A1 => n37914, A2 => n37913, A3 => n37912, A4 => 
                           n37911, ZN => n37915);
   U3332 : AOI22_X1 port map( A1 => n38159, A2 => n37916, B1 => n38337, B2 => 
                           n37915, ZN => n37917);
   U3333 : OAI21_X1 port map( B1 => n38342, B2 => n37918, A => n37917, ZN => 
                           OUT1(19));
   U3334 : AOI22_X1 port map( A1 => n29504, A2 => n30058, B1 => n29563, B2 => 
                           n30067, ZN => n37922);
   U3335 : AOI22_X1 port map( A1 => n29956, A2 => n30054, B1 => n29540, B2 => 
                           n30063, ZN => n37921);
   U3336 : AOI22_X1 port map( A1 => n29562, A2 => n30062, B1 => n29974, B2 => 
                           n30057, ZN => n37920);
   U3337 : AOI22_X1 port map( A1 => n30004, A2 => n30065, B1 => n29270, B2 => 
                           n31178, ZN => n37919);
   U3338 : NAND4_X1 port map( A1 => n37922, A2 => n37921, A3 => n37920, A4 => 
                           n37919, ZN => n37928);
   U3339 : AOI22_X1 port map( A1 => n29559, A2 => n31175, B1 => n29995, B2 => 
                           n31174, ZN => n37926);
   U3340 : AOI22_X1 port map( A1 => n30024, A2 => n31198, B1 => n29333, B2 => 
                           n31173, ZN => n37925);
   U3341 : AOI22_X1 port map( A1 => n29979, A2 => n30060, B1 => n29552, B2 => 
                           n31184, ZN => n37924);
   U3342 : AOI22_X1 port map( A1 => n29470, A2 => n30066, B1 => n29561, B2 => 
                           n31195, ZN => n37923);
   U3343 : NAND4_X1 port map( A1 => n37926, A2 => n37925, A3 => n37924, A4 => 
                           n37923, ZN => n37927);
   U3344 : NOR2_X1 port map( A1 => n37928, A2 => n37927, ZN => n37940);
   U3345 : AOI22_X1 port map( A1 => n29840, A2 => n31191, B1 => n29842, B2 => 
                           n31159, ZN => n37932);
   U3346 : AOI22_X1 port map( A1 => n29843, A2 => n30127, B1 => n29845, B2 => 
                           n30126, ZN => n37931);
   U3347 : AOI22_X1 port map( A1 => n29841, A2 => n30125, B1 => n29881, B2 => 
                           n31166, ZN => n37930);
   U3348 : AOI22_X1 port map( A1 => n29839, A2 => n31180, B1 => n29844, B2 => 
                           n31182, ZN => n37929);
   U3349 : NAND4_X1 port map( A1 => n37932, A2 => n37931, A3 => n37930, A4 => 
                           n37929, ZN => n37938);
   U3350 : AOI22_X1 port map( A1 => n29679, A2 => n31167, B1 => n29386, B2 => 
                           n30128, ZN => n37936);
   U3351 : AOI22_X1 port map( A1 => n29362, A2 => n31160, B1 => n29452, B2 => 
                           n31159, ZN => n37935);
   U3352 : AOI22_X1 port map( A1 => n29416, A2 => n31187, B1 => n29689, B2 => 
                           n30052, ZN => n37934);
   U3353 : AOI22_X1 port map( A1 => n29709, A2 => n31166, B1 => n29584, B2 => 
                           n31194, ZN => n37933);
   U3354 : NAND4_X1 port map( A1 => n37936, A2 => n37935, A3 => n37934, A4 => 
                           n37933, ZN => n37937);
   U3355 : AOI22_X1 port map( A1 => n38159, A2 => n37938, B1 => n38337, B2 => 
                           n37937, ZN => n37939);
   U3356 : OAI21_X1 port map( B1 => n38342, B2 => n37940, A => n37939, ZN => 
                           OUT1(18));
   U3357 : AOI22_X1 port map( A1 => n29318, A2 => n30053, B1 => n29322, B2 => 
                           n30064, ZN => n37944);
   U3358 : AOI22_X1 port map( A1 => n29310, A2 => n30056, B1 => n29323, B2 => 
                           n30067, ZN => n37943);
   U3359 : AOI22_X1 port map( A1 => n29321, A2 => n31177, B1 => n30026, B2 => 
                           n30059, ZN => n37942);
   U3360 : AOI22_X1 port map( A1 => n29282, A2 => n31178, B1 => n30001, B2 => 
                           n30055, ZN => n37941);
   U3361 : NAND4_X1 port map( A1 => n37944, A2 => n37943, A3 => n37942, A4 => 
                           n37941, ZN => n37950);
   U3362 : AOI22_X1 port map( A1 => n29325, A2 => n30062, B1 => n30005, B2 => 
                           n30065, ZN => n37948);
   U3363 : AOI22_X1 port map( A1 => n29320, A2 => n31188, B1 => n29969, B2 => 
                           n30060, ZN => n37947);
   U3364 : AOI22_X1 port map( A1 => n29319, A2 => n30068, B1 => n30008, B2 => 
                           n31197, ZN => n37946);
   U3365 : AOI22_X1 port map( A1 => n29311, A2 => n31183, B1 => n29976, B2 => 
                           n30057, ZN => n37945);
   U3366 : NAND4_X1 port map( A1 => n37948, A2 => n37947, A3 => n37946, A4 => 
                           n37945, ZN => n37949);
   U3367 : NOR2_X1 port map( A1 => n37950, A2 => n37949, ZN => n37962);
   U3368 : AOI22_X1 port map( A1 => n29766, A2 => n30126, B1 => n29772, B2 => 
                           n31190, ZN => n37954);
   U3369 : AOI22_X1 port map( A1 => n29764, A2 => n31164, B1 => n29873, B2 => 
                           n31166, ZN => n37953);
   U3370 : AOI22_X1 port map( A1 => n29765, A2 => n31170, B1 => n29770, B2 => 
                           n31191, ZN => n37952);
   U3371 : AOI22_X1 port map( A1 => n29768, A2 => n30128, B1 => n29774, B2 => 
                           n31171, ZN => n37951);
   U3372 : NAND4_X1 port map( A1 => n37954, A2 => n37953, A3 => n37952, A4 => 
                           n37951, ZN => n37960);
   U3373 : AOI22_X1 port map( A1 => n29315, A2 => n31190, B1 => n29163, B2 => 
                           n30126, ZN => n37958);
   U3374 : AOI22_X1 port map( A1 => n29312, A2 => n31169, B1 => n29145, B2 => 
                           n31166, ZN => n37957);
   U3375 : AOI22_X1 port map( A1 => n29313, A2 => n31160, B1 => n29314, B2 => 
                           n30125, ZN => n37956);
   U3376 : AOI22_X1 port map( A1 => n29118, A2 => n31171, B1 => n29160, B2 => 
                           n30052, ZN => n37955);
   U3377 : NAND4_X1 port map( A1 => n37958, A2 => n37957, A3 => n37956, A4 => 
                           n37955, ZN => n37959);
   U3378 : AOI22_X1 port map( A1 => n38159, A2 => n37960, B1 => n38337, B2 => 
                           n37959, ZN => n37961);
   U3379 : OAI21_X1 port map( B1 => n38342, B2 => n37962, A => n37961, ZN => 
                           OUT1(17));
   U3380 : AOI22_X1 port map( A1 => n30006, A2 => n31185, B1 => n30009, B2 => 
                           n31174, ZN => n37966);
   U3381 : AOI22_X1 port map( A1 => n29280, A2 => n30063, B1 => n29268, B2 => 
                           n31178, ZN => n37965);
   U3382 : AOI22_X1 port map( A1 => n29291, A2 => n30058, B1 => n29977, B2 => 
                           n31181, ZN => n37964);
   U3383 : AOI22_X1 port map( A1 => n29290, A2 => n30066, B1 => n29265, B2 => 
                           n31189, ZN => n37963);
   U3384 : NAND4_X1 port map( A1 => n37966, A2 => n37965, A3 => n37964, A4 => 
                           n37963, ZN => n37972);
   U3385 : AOI22_X1 port map( A1 => n29949, A2 => n30054, B1 => n29967, B2 => 
                           n31176, ZN => n37970);
   U3386 : AOI22_X1 port map( A1 => n29975, A2 => n30059, B1 => n29289, B2 => 
                           n31173, ZN => n37969);
   U3387 : AOI22_X1 port map( A1 => n29264, A2 => n30062, B1 => n29277, B2 => 
                           n30053, ZN => n37968);
   U3388 : AOI22_X1 port map( A1 => n29279, A2 => n30068, B1 => n29285, B2 => 
                           n30064, ZN => n37967);
   U3389 : NAND4_X1 port map( A1 => n37970, A2 => n37969, A3 => n37968, A4 => 
                           n37967, ZN => n37971);
   U3390 : NOR2_X1 port map( A1 => n37972, A2 => n37971, ZN => n37984);
   U3391 : AOI22_X1 port map( A1 => n29858, A2 => n31160, B1 => n29861, B2 => 
                           n30127, ZN => n37976);
   U3392 : AOI22_X1 port map( A1 => n29769, A2 => n30051, B1 => n29862, B2 => 
                           n30052, ZN => n37975);
   U3393 : AOI22_X1 port map( A1 => n29859, A2 => n30125, B1 => n29860, B2 => 
                           n31190, ZN => n37974);
   U3394 : AOI22_X1 port map( A1 => n29863, A2 => n31167, B1 => n29856, B2 => 
                           n31169, ZN => n37973);
   U3395 : NAND4_X1 port map( A1 => n37976, A2 => n37975, A3 => n37974, A4 => 
                           n37973, ZN => n37982);
   U3396 : AOI22_X1 port map( A1 => n29292, A2 => n31169, B1 => n29693, B2 => 
                           n31170, ZN => n37980);
   U3397 : AOI22_X1 port map( A1 => n29295, A2 => n31159, B1 => n29680, B2 => 
                           n30126, ZN => n37979);
   U3398 : AOI22_X1 port map( A1 => n29697, A2 => n31166, B1 => n29586, B2 => 
                           n31171, ZN => n37978);
   U3399 : AOI22_X1 port map( A1 => n29294, A2 => n31164, B1 => n29293, B2 => 
                           n31179, ZN => n37977);
   U3400 : NAND4_X1 port map( A1 => n37980, A2 => n37979, A3 => n37978, A4 => 
                           n37977, ZN => n37981);
   U3401 : AOI22_X1 port map( A1 => n38159, A2 => n37982, B1 => n38337, B2 => 
                           n37981, ZN => n37983);
   U3402 : OAI21_X1 port map( B1 => n38342, B2 => n37984, A => n37983, ZN => 
                           OUT1(16));
   U3403 : AOI22_X1 port map( A1 => n29529, A2 => n30062, B1 => n30027, B2 => 
                           n30059, ZN => n37988);
   U3404 : AOI22_X1 port map( A1 => n29528, A2 => n30067, B1 => n29525, B2 => 
                           n30053, ZN => n37987);
   U3405 : AOI22_X1 port map( A1 => n29526, A2 => n30068, B1 => n29332, B2 => 
                           n30056, ZN => n37986);
   U3406 : AOI22_X1 port map( A1 => n29503, A2 => n30058, B1 => n29965, B2 => 
                           n30060, ZN => n37985);
   U3407 : NAND4_X1 port map( A1 => n37988, A2 => n37987, A3 => n37986, A4 => 
                           n37985, ZN => n37994);
   U3408 : AOI22_X1 port map( A1 => n29471, A2 => n30066, B1 => n30007, B2 => 
                           n30065, ZN => n37992);
   U3409 : AOI22_X1 port map( A1 => n30002, A2 => n31174, B1 => n29527, B2 => 
                           n30063, ZN => n37991);
   U3410 : AOI22_X1 port map( A1 => n29524, A2 => n31195, B1 => n29269, B2 => 
                           n30061, ZN => n37990);
   U3411 : AOI22_X1 port map( A1 => n29978, A2 => n30057, B1 => n29954, B2 => 
                           n30054, ZN => n37989);
   U3412 : NAND4_X1 port map( A1 => n37992, A2 => n37991, A3 => n37990, A4 => 
                           n37989, ZN => n37993);
   U3413 : NOR2_X1 port map( A1 => n37994, A2 => n37993, ZN => n38006);
   U3414 : AOI22_X1 port map( A1 => n29821, A2 => n31194, B1 => n29811, B2 => 
                           n31193, ZN => n37998);
   U3415 : AOI22_X1 port map( A1 => n29812, A2 => n31164, B1 => n29815, B2 => 
                           n31179, ZN => n37997);
   U3416 : AOI22_X1 port map( A1 => n29816, A2 => n31180, B1 => n29810, B2 => 
                           n31182, ZN => n37996);
   U3417 : AOI22_X1 port map( A1 => n29799, A2 => n31192, B1 => n29904, B2 => 
                           n31186, ZN => n37995);
   U3418 : NAND4_X1 port map( A1 => n37998, A2 => n37997, A3 => n37996, A4 => 
                           n37995, ZN => n38004);
   U3419 : AOI22_X1 port map( A1 => n29361, A2 => n31160, B1 => n29451, B2 => 
                           n31193, ZN => n38002);
   U3420 : AOI22_X1 port map( A1 => n29162, A2 => n31192, B1 => n29387, B2 => 
                           n31169, ZN => n38001);
   U3421 : AOI22_X1 port map( A1 => n29122, A2 => n30127, B1 => n29146, B2 => 
                           n30052, ZN => n38000);
   U3422 : AOI22_X1 port map( A1 => n29415, A2 => n31164, B1 => n29148, B2 => 
                           n31166, ZN => n37999);
   U3423 : NAND4_X1 port map( A1 => n38002, A2 => n38001, A3 => n38000, A4 => 
                           n37999, ZN => n38003);
   U3424 : AOI22_X1 port map( A1 => n38159, A2 => n38004, B1 => n38337, B2 => 
                           n38003, ZN => n38005);
   U3425 : OAI21_X1 port map( B1 => n38342, B2 => n38006, A => n38005, ZN => 
                           OUT1(15));
   U3426 : AOI22_X1 port map( A1 => n29331, A2 => n31173, B1 => n29574, B2 => 
                           n31196, ZN => n38010);
   U3427 : AOI22_X1 port map( A1 => n30000, A2 => n31174, B1 => n29544, B2 => 
                           n31188, ZN => n38009);
   U3428 : AOI22_X1 port map( A1 => n29986, A2 => n30057, B1 => n29560, B2 => 
                           n30053, ZN => n38008);
   U3429 : AOI22_X1 port map( A1 => n29577, A2 => n30067, B1 => n29523, B2 => 
                           n31195, ZN => n38007);
   U3430 : NAND4_X1 port map( A1 => n38010, A2 => n38009, A3 => n38008, A4 => 
                           n38007, ZN => n38016);
   U3431 : AOI22_X1 port map( A1 => n30011, A2 => n30065, B1 => n29942, B2 => 
                           n31197, ZN => n38014);
   U3432 : AOI22_X1 port map( A1 => n30020, A2 => n30059, B1 => n29473, B2 => 
                           n30066, ZN => n38013);
   U3433 : AOI22_X1 port map( A1 => n29963, A2 => n31176, B1 => n29502, B2 => 
                           n31177, ZN => n38012);
   U3434 : AOI22_X1 port map( A1 => n29553, A2 => n31184, B1 => n29266, B2 => 
                           n30061, ZN => n38011);
   U3435 : NAND4_X1 port map( A1 => n38014, A2 => n38013, A3 => n38012, A4 => 
                           n38011, ZN => n38015);
   U3436 : NOR2_X1 port map( A1 => n38016, A2 => n38015, ZN => n38028);
   U3437 : AOI22_X1 port map( A1 => n29901, A2 => n31194, B1 => n29902, B2 => 
                           n31159, ZN => n38020);
   U3438 : AOI22_X1 port map( A1 => n29903, A2 => n31164, B1 => n29906, B2 => 
                           n31180, ZN => n38019);
   U3439 : AOI22_X1 port map( A1 => n29908, A2 => n31170, B1 => n29907, B2 => 
                           n31192, ZN => n38018);
   U3440 : AOI22_X1 port map( A1 => n29778, A2 => n31186, B1 => n29905, B2 => 
                           n31160, ZN => n38017);
   U3441 : NAND4_X1 port map( A1 => n38020, A2 => n38019, A3 => n38018, A4 => 
                           n38017, ZN => n38026);
   U3442 : AOI22_X1 port map( A1 => n29408, A2 => n31187, B1 => n29448, B2 => 
                           n31159, ZN => n38024);
   U3443 : AOI22_X1 port map( A1 => n29388, A2 => n31180, B1 => n29674, B2 => 
                           n31166, ZN => n38023);
   U3444 : AOI22_X1 port map( A1 => n29578, A2 => n31194, B1 => n29695, B2 => 
                           n31170, ZN => n38022);
   U3445 : AOI22_X1 port map( A1 => n29672, A2 => n31192, B1 => n29360, B2 => 
                           n31191, ZN => n38021);
   U3446 : NAND4_X1 port map( A1 => n38024, A2 => n38023, A3 => n38022, A4 => 
                           n38021, ZN => n38025);
   U3447 : AOI22_X1 port map( A1 => n38159, A2 => n38026, B1 => n38337, B2 => 
                           n38025, ZN => n38027);
   U3448 : OAI21_X1 port map( B1 => n38342, B2 => n38028, A => n38027, ZN => 
                           OUT1(14));
   U3449 : AOI22_X1 port map( A1 => n29515, A2 => n31175, B1 => n29501, B2 => 
                           n30058, ZN => n38032);
   U3450 : AOI22_X1 port map( A1 => n29519, A2 => n30067, B1 => n29987, B2 => 
                           n31181, ZN => n38031);
   U3451 : AOI22_X1 port map( A1 => n29517, A2 => n30063, B1 => n29958, B2 => 
                           n30059, ZN => n38030);
   U3452 : AOI22_X1 port map( A1 => n29518, A2 => n30064, B1 => n29520, B2 => 
                           n31196, ZN => n38029);
   U3453 : NAND4_X1 port map( A1 => n38032, A2 => n38031, A3 => n38030, A4 => 
                           n38029, ZN => n38038);
   U3454 : AOI22_X1 port map( A1 => n29474, A2 => n30066, B1 => n29516, B2 => 
                           n30068, ZN => n38036);
   U3455 : AOI22_X1 port map( A1 => n29941, A2 => n31197, B1 => n29961, B2 => 
                           n31176, ZN => n38035);
   U3456 : AOI22_X1 port map( A1 => n30012, A2 => n30065, B1 => n29998, B2 => 
                           n30055, ZN => n38034);
   U3457 : AOI22_X1 port map( A1 => n29329, A2 => n30056, B1 => n29267, B2 => 
                           n30061, ZN => n38033);
   U3458 : NAND4_X1 port map( A1 => n38036, A2 => n38035, A3 => n38034, A4 => 
                           n38033, ZN => n38037);
   U3459 : NOR2_X1 port map( A1 => n38038, A2 => n38037, ZN => n38050);
   U3460 : AOI22_X1 port map( A1 => n29887, A2 => n31167, B1 => n29893, B2 => 
                           n31160, ZN => n38042);
   U3461 : AOI22_X1 port map( A1 => n29885, A2 => n31171, B1 => n29886, B2 => 
                           n30052, ZN => n38041);
   U3462 : AOI22_X1 port map( A1 => n29894, A2 => n31187, B1 => n29884, B2 => 
                           n31190, ZN => n38040);
   U3463 : AOI22_X1 port map( A1 => n29892, A2 => n30128, B1 => n29888, B2 => 
                           n30051, ZN => n38039);
   U3464 : NAND4_X1 port map( A1 => n38042, A2 => n38041, A3 => n38040, A4 => 
                           n38039, ZN => n38048);
   U3465 : AOI22_X1 port map( A1 => n29359, A2 => n31160, B1 => n29691, B2 => 
                           n31186, ZN => n38046);
   U3466 : AOI22_X1 port map( A1 => n29708, A2 => n31170, B1 => n29447, B2 => 
                           n31159, ZN => n38045);
   U3467 : AOI22_X1 port map( A1 => n29701, A2 => n31192, B1 => n29405, B2 => 
                           n30125, ZN => n38044);
   U3468 : AOI22_X1 port map( A1 => n29585, A2 => n31194, B1 => n29394, B2 => 
                           n30128, ZN => n38043);
   U3469 : NAND4_X1 port map( A1 => n38046, A2 => n38045, A3 => n38044, A4 => 
                           n38043, ZN => n38047);
   U3470 : AOI22_X1 port map( A1 => n38159, A2 => n38048, B1 => n38337, B2 => 
                           n38047, ZN => n38049);
   U3471 : OAI21_X1 port map( B1 => n38342, B2 => n38050, A => n38049, ZN => 
                           OUT1(13));
   U3472 : AOI22_X1 port map( A1 => n29512, A2 => n31189, B1 => n29959, B2 => 
                           n30054, ZN => n38054);
   U3473 : AOI22_X1 port map( A1 => n29500, A2 => n30058, B1 => n29508, B2 => 
                           n30053, ZN => n38053);
   U3474 : AOI22_X1 port map( A1 => n29513, A2 => n30062, B1 => n29989, B2 => 
                           n30057, ZN => n38052);
   U3475 : AOI22_X1 port map( A1 => n29475, A2 => n30066, B1 => n29511, B2 => 
                           n30064, ZN => n38051);
   U3476 : NAND4_X1 port map( A1 => n38054, A2 => n38053, A3 => n38052, A4 => 
                           n38051, ZN => n38060);
   U3477 : AOI22_X1 port map( A1 => n29509, A2 => n30068, B1 => n29510, B2 => 
                           n30063, ZN => n38058);
   U3478 : AOI22_X1 port map( A1 => n29955, A2 => n31198, B1 => n29328, B2 => 
                           n30056, ZN => n38057);
   U3479 : AOI22_X1 port map( A1 => n29997, A2 => n30055, B1 => n29947, B2 => 
                           n30060, ZN => n38056);
   U3480 : AOI22_X1 port map( A1 => n30013, A2 => n31185, B1 => n29263, B2 => 
                           n30061, ZN => n38055);
   U3481 : NAND4_X1 port map( A1 => n38058, A2 => n38057, A3 => n38056, A4 => 
                           n38055, ZN => n38059);
   U3482 : NOR2_X1 port map( A1 => n38060, A2 => n38059, ZN => n38072);
   U3483 : AOI22_X1 port map( A1 => n29877, A2 => n31182, B1 => n29879, B2 => 
                           n31186, ZN => n38064);
   U3484 : AOI22_X1 port map( A1 => n29882, A2 => n31169, B1 => n29874, B2 => 
                           n31187, ZN => n38063);
   U3485 : AOI22_X1 port map( A1 => n29883, A2 => n31160, B1 => n29875, B2 => 
                           n31159, ZN => n38062);
   U3486 : AOI22_X1 port map( A1 => n29878, A2 => n31192, B1 => n29876, B2 => 
                           n30127, ZN => n38061);
   U3487 : NAND4_X1 port map( A1 => n38064, A2 => n38063, A3 => n38062, A4 => 
                           n38061, ZN => n38070);
   U3488 : AOI22_X1 port map( A1 => n29593, A2 => n31171, B1 => n29699, B2 => 
                           n31170, ZN => n38068);
   U3489 : AOI22_X1 port map( A1 => n29669, A2 => n31192, B1 => n29446, B2 => 
                           n31190, ZN => n38067);
   U3490 : AOI22_X1 port map( A1 => n29358, A2 => n31160, B1 => n29670, B2 => 
                           n30051, ZN => n38066);
   U3491 : AOI22_X1 port map( A1 => n29395, A2 => n30128, B1 => n29404, B2 => 
                           n31164, ZN => n38065);
   U3492 : NAND4_X1 port map( A1 => n38068, A2 => n38067, A3 => n38066, A4 => 
                           n38065, ZN => n38069);
   U3493 : AOI22_X1 port map( A1 => n38159, A2 => n38070, B1 => n38337, B2 => 
                           n38069, ZN => n38071);
   U3494 : OAI21_X1 port map( B1 => n38342, B2 => n38072, A => n38071, ZN => 
                           OUT1(12));
   U3495 : AOI22_X1 port map( A1 => n29327, A2 => n31173, B1 => n29498, B2 => 
                           n31189, ZN => n38076);
   U3496 : AOI22_X1 port map( A1 => n29324, A2 => n31178, B1 => n29493, B2 => 
                           n30053, ZN => n38075);
   U3497 : AOI22_X1 port map( A1 => n29494, A2 => n30068, B1 => n29495, B2 => 
                           n31188, ZN => n38074);
   U3498 : AOI22_X1 port map( A1 => n30014, A2 => n31185, B1 => n29497, B2 => 
                           n31195, ZN => n38073);
   U3499 : NAND4_X1 port map( A1 => n38076, A2 => n38075, A3 => n38074, A4 => 
                           n38073, ZN => n38082);
   U3500 : AOI22_X1 port map( A1 => n29971, A2 => n31176, B1 => n29996, B2 => 
                           n30055, ZN => n38080);
   U3501 : AOI22_X1 port map( A1 => n29476, A2 => n31183, B1 => n29496, B2 => 
                           n30058, ZN => n38079);
   U3502 : AOI22_X1 port map( A1 => n29499, A2 => n30062, B1 => n29943, B2 => 
                           n30054, ZN => n38078);
   U3503 : AOI22_X1 port map( A1 => n29951, A2 => n30059, B1 => n29990, B2 => 
                           n30057, ZN => n38077);
   U3504 : NAND4_X1 port map( A1 => n38080, A2 => n38079, A3 => n38078, A4 => 
                           n38077, ZN => n38081);
   U3505 : NOR2_X1 port map( A1 => n38082, A2 => n38081, ZN => n38094);
   U3506 : AOI22_X1 port map( A1 => n29870, A2 => n31166, B1 => n29867, B2 => 
                           n31171, ZN => n38086);
   U3507 : AOI22_X1 port map( A1 => n29865, A2 => n31159, B1 => n29857, B2 => 
                           n31191, ZN => n38085);
   U3508 : AOI22_X1 port map( A1 => n29864, A2 => n31164, B1 => n29869, B2 => 
                           n30126, ZN => n38084);
   U3509 : AOI22_X1 port map( A1 => n29868, A2 => n31182, B1 => n29871, B2 => 
                           n31180, ZN => n38083);
   U3510 : NAND4_X1 port map( A1 => n38086, A2 => n38085, A3 => n38084, A4 => 
                           n38083, ZN => n38092);
   U3511 : AOI22_X1 port map( A1 => n29683, A2 => n31166, B1 => n29399, B2 => 
                           n30125, ZN => n38090);
   U3512 : AOI22_X1 port map( A1 => n29357, A2 => n31191, B1 => n29445, B2 => 
                           n31159, ZN => n38089);
   U3513 : AOI22_X1 port map( A1 => n29592, A2 => n30127, B1 => n29700, B2 => 
                           n31170, ZN => n38088);
   U3514 : AOI22_X1 port map( A1 => n29703, A2 => n30126, B1 => n29396, B2 => 
                           n31180, ZN => n38087);
   U3515 : NAND4_X1 port map( A1 => n38090, A2 => n38089, A3 => n38088, A4 => 
                           n38087, ZN => n38091);
   U3516 : AOI22_X1 port map( A1 => n38159, A2 => n38092, B1 => n38337, B2 => 
                           n38091, ZN => n38093);
   U3517 : OAI21_X1 port map( B1 => n38342, B2 => n38094, A => n38093, ZN => 
                           OUT1(11));
   U3518 : AOI22_X1 port map( A1 => n29718, A2 => n31181, B1 => n29326, B2 => 
                           n31173, ZN => n38098);
   U3519 : AOI22_X1 port map( A1 => n29251, A2 => n30067, B1 => n29490, B2 => 
                           n30062, ZN => n38097);
   U3520 : AOI22_X1 port map( A1 => n29485, A2 => n31175, B1 => n29716, B2 => 
                           n30055, ZN => n38096);
   U3521 : AOI22_X1 port map( A1 => n29530, A2 => n30061, B1 => n29714, B2 => 
                           n31176, ZN => n38095);
   U3522 : NAND4_X1 port map( A1 => n38098, A2 => n38097, A3 => n38096, A4 => 
                           n38095, ZN => n38104);
   U3523 : AOI22_X1 port map( A1 => n29715, A2 => n30054, B1 => n29486, B2 => 
                           n31184, ZN => n38102);
   U3524 : AOI22_X1 port map( A1 => n29477, A2 => n31183, B1 => n29719, B2 => 
                           n30065, ZN => n38101);
   U3525 : AOI22_X1 port map( A1 => n29489, A2 => n30064, B1 => n29487, B2 => 
                           n31188, ZN => n38100);
   U3526 : AOI22_X1 port map( A1 => n29488, A2 => n31177, B1 => n29717, B2 => 
                           n31198, ZN => n38099);
   U3527 : NAND4_X1 port map( A1 => n38102, A2 => n38101, A3 => n38100, A4 => 
                           n38099, ZN => n38103);
   U3528 : NOR2_X1 port map( A1 => n38104, A2 => n38103, ZN => n38116);
   U3529 : AOI22_X1 port map( A1 => n29259, A2 => n30125, B1 => n29252, B2 => 
                           n31182, ZN => n38108);
   U3530 : AOI22_X1 port map( A1 => n29249, A2 => n31167, B1 => n29250, B2 => 
                           n31166, ZN => n38107);
   U3531 : AOI22_X1 port map( A1 => n29256, A2 => n31171, B1 => n29253, B2 => 
                           n31159, ZN => n38106);
   U3532 : AOI22_X1 port map( A1 => n29257, A2 => n31180, B1 => n29254, B2 => 
                           n31179, ZN => n38105);
   U3533 : NAND4_X1 port map( A1 => n38108, A2 => n38107, A3 => n38106, A4 => 
                           n38105, ZN => n38114);
   U3534 : AOI22_X1 port map( A1 => n29258, A2 => n31164, B1 => n29442, B2 => 
                           n31159, ZN => n38112);
   U3535 : AOI22_X1 port map( A1 => n29590, A2 => n31194, B1 => n29686, B2 => 
                           n31166, ZN => n38111);
   U3536 : AOI22_X1 port map( A1 => n29676, A2 => n31167, B1 => n29255, B2 => 
                           n31180, ZN => n38110);
   U3537 : AOI22_X1 port map( A1 => n29710, A2 => n31182, B1 => n29354, B2 => 
                           n31179, ZN => n38109);
   U3538 : NAND4_X1 port map( A1 => n38112, A2 => n38111, A3 => n38110, A4 => 
                           n38109, ZN => n38113);
   U3539 : AOI22_X1 port map( A1 => n38159, A2 => n38114, B1 => n38337, B2 => 
                           n38113, ZN => n38115);
   U3540 : OAI21_X1 port map( B1 => n38295, B2 => n38116, A => n38115, ZN => 
                           OUT1(10));
   U3541 : AOI22_X1 port map( A1 => n29533, A2 => n30068, B1 => n30015, B2 => 
                           n30065, ZN => n38120);
   U3542 : AOI22_X1 port map( A1 => n29534, A2 => n31178, B1 => n29484, B2 => 
                           n31175, ZN => n38119);
   U3543 : AOI22_X1 port map( A1 => n29522, A2 => n30064, B1 => n29994, B2 => 
                           n31174, ZN => n38118);
   U3544 : AOI22_X1 port map( A1 => n29317, A2 => n30056, B1 => n29535, B2 => 
                           n30062, ZN => n38117);
   U3545 : NAND4_X1 port map( A1 => n38120, A2 => n38119, A3 => n38118, A4 => 
                           n38117, ZN => n38126);
   U3546 : AOI22_X1 port map( A1 => n29492, A2 => n30058, B1 => n29992, B2 => 
                           n30057, ZN => n38124);
   U3547 : AOI22_X1 port map( A1 => n29532, A2 => n31188, B1 => n29970, B2 => 
                           n30060, ZN => n38123);
   U3548 : AOI22_X1 port map( A1 => n29478, A2 => n30066, B1 => n29531, B2 => 
                           n30067, ZN => n38122);
   U3549 : AOI22_X1 port map( A1 => n29950, A2 => n30059, B1 => n29962, B2 => 
                           n30054, ZN => n38121);
   U3550 : NAND4_X1 port map( A1 => n38124, A2 => n38123, A3 => n38122, A4 => 
                           n38121, ZN => n38125);
   U3551 : NOR2_X1 port map( A1 => n38126, A2 => n38125, ZN => n38138);
   U3552 : AOI22_X1 port map( A1 => n29935, A2 => n31164, B1 => n29940, B2 => 
                           n31186, ZN => n38130);
   U3553 : AOI22_X1 port map( A1 => n29937, A2 => n31159, B1 => n29933, B2 => 
                           n31191, ZN => n38129);
   U3554 : AOI22_X1 port map( A1 => n29934, A2 => n31169, B1 => n29939, B2 => 
                           n30127, ZN => n38128);
   U3555 : AOI22_X1 port map( A1 => n29936, A2 => n30126, B1 => n29938, B2 => 
                           n31170, ZN => n38127);
   U3556 : NAND4_X1 port map( A1 => n38130, A2 => n38129, A3 => n38128, A4 => 
                           n38127, ZN => n38136);
   U3557 : AOI22_X1 port map( A1 => n29711, A2 => n31166, B1 => n29702, B2 => 
                           n31170, ZN => n38134);
   U3558 : AOI22_X1 port map( A1 => n29677, A2 => n31167, B1 => n29580, B2 => 
                           n31194, ZN => n38133);
   U3559 : AOI22_X1 port map( A1 => n29355, A2 => n31191, B1 => n29398, B2 => 
                           n31187, ZN => n38132);
   U3560 : AOI22_X1 port map( A1 => n29402, A2 => n30128, B1 => n29440, B2 => 
                           n31193, ZN => n38131);
   U3561 : NAND4_X1 port map( A1 => n38134, A2 => n38133, A3 => n38132, A4 => 
                           n38131, ZN => n38135);
   U3562 : AOI22_X1 port map( A1 => n38159, A2 => n38136, B1 => n38337, B2 => 
                           n38135, ZN => n38137);
   U3563 : OAI21_X1 port map( B1 => n38342, B2 => n38138, A => n38137, ZN => 
                           OUT1(9));
   U3564 : AOI22_X1 port map( A1 => n29968, A2 => n31176, B1 => n29546, B2 => 
                           n30062, ZN => n38142);
   U3565 : AOI22_X1 port map( A1 => n29521, A2 => n30064, B1 => n29542, B2 => 
                           n30068, ZN => n38141);
   U3566 : AOI22_X1 port map( A1 => n29545, A2 => n31178, B1 => n29543, B2 => 
                           n31175, ZN => n38140);
   U3567 : AOI22_X1 port map( A1 => n29985, A2 => n31174, B1 => n30016, B2 => 
                           n30065, ZN => n38139);
   U3568 : NAND4_X1 port map( A1 => n38142, A2 => n38141, A3 => n38140, A4 => 
                           n38139, ZN => n38148);
   U3569 : AOI22_X1 port map( A1 => n29547, A2 => n30067, B1 => n29973, B2 => 
                           n30054, ZN => n38146);
   U3570 : AOI22_X1 port map( A1 => n29491, A2 => n30058, B1 => n29479, B2 => 
                           n30066, ZN => n38145);
   U3571 : AOI22_X1 port map( A1 => n29993, A2 => n30057, B1 => n29948, B2 => 
                           n30059, ZN => n38144);
   U3572 : AOI22_X1 port map( A1 => n29316, A2 => n30056, B1 => n29541, B2 => 
                           n31188, ZN => n38143);
   U3573 : NAND4_X1 port map( A1 => n38146, A2 => n38145, A3 => n38144, A4 => 
                           n38143, ZN => n38147);
   U3574 : NOR2_X1 port map( A1 => n38148, A2 => n38147, ZN => n38161);
   U3575 : AOI22_X1 port map( A1 => n29923, A2 => n31170, B1 => n29919, B2 => 
                           n31187, ZN => n38152);
   U3576 : AOI22_X1 port map( A1 => n29922, A2 => n31186, B1 => n29925, B2 => 
                           n31180, ZN => n38151);
   U3577 : AOI22_X1 port map( A1 => n29920, A2 => n31171, B1 => n29921, B2 => 
                           n30126, ZN => n38150);
   U3578 : AOI22_X1 port map( A1 => n29918, A2 => n31179, B1 => n29924, B2 => 
                           n31193, ZN => n38149);
   U3579 : NAND4_X1 port map( A1 => n38152, A2 => n38151, A3 => n38150, A4 => 
                           n38149, ZN => n38158);
   U3580 : AOI22_X1 port map( A1 => n29678, A2 => n31166, B1 => n29705, B2 => 
                           n31182, ZN => n38156);
   U3581 : AOI22_X1 port map( A1 => n29397, A2 => n30125, B1 => n29438, B2 => 
                           n31193, ZN => n38155);
   U3582 : AOI22_X1 port map( A1 => n29582, A2 => n31171, B1 => n29673, B2 => 
                           n31192, ZN => n38154);
   U3583 : AOI22_X1 port map( A1 => n29356, A2 => n31191, B1 => n29403, B2 => 
                           n31169, ZN => n38153);
   U3584 : NAND4_X1 port map( A1 => n38156, A2 => n38155, A3 => n38154, A4 => 
                           n38153, ZN => n38157);
   U3585 : AOI22_X1 port map( A1 => n38159, A2 => n38158, B1 => n38337, B2 => 
                           n38157, ZN => n38160);
   U3586 : OAI21_X1 port map( B1 => n38342, B2 => n38161, A => n38160, ZN => 
                           OUT1(8));
   U3587 : AOI22_X1 port map( A1 => n29018, A2 => n30067, B1 => n29023, B2 => 
                           n30053, ZN => n38165);
   U3588 : AOI22_X1 port map( A1 => n29668, A2 => n31176, B1 => n29038, B2 => 
                           n30056, ZN => n38164);
   U3589 : AOI22_X1 port map( A1 => n29663, A2 => n31174, B1 => n29035, B2 => 
                           n30058, ZN => n38163);
   U3590 : AOI22_X1 port map( A1 => n29665, A2 => n30059, B1 => n29020, B2 => 
                           n30061, ZN => n38162);
   U3591 : NAND4_X1 port map( A1 => n38165, A2 => n38164, A3 => n38163, A4 => 
                           n38162, ZN => n38171);
   U3592 : AOI22_X1 port map( A1 => n29019, A2 => n31195, B1 => n29028, B2 => 
                           n31196, ZN => n38169);
   U3593 : AOI22_X1 port map( A1 => n29047, A2 => n31183, B1 => n29666, B2 => 
                           n30057, ZN => n38168);
   U3594 : AOI22_X1 port map( A1 => n29664, A2 => n31197, B1 => n29667, B2 => 
                           n30065, ZN => n38167);
   U3595 : AOI22_X1 port map( A1 => n29033, A2 => n30063, B1 => n29024, B2 => 
                           n30068, ZN => n38166);
   U3596 : NAND4_X1 port map( A1 => n38169, A2 => n38168, A3 => n38167, A4 => 
                           n38166, ZN => n38170);
   U3597 : NOR2_X1 port map( A1 => n38171, A2 => n38170, ZN => n38184);
   U3598 : CLKBUF_X1 port map( A => n38172, Z => n38339);
   U3599 : AOI22_X1 port map( A1 => n29239, A2 => n31187, B1 => n29246, B2 => 
                           n31179, ZN => n38176);
   U3600 : AOI22_X1 port map( A1 => n29247, A2 => n31159, B1 => n29244, B2 => 
                           n31167, ZN => n38175);
   U3601 : AOI22_X1 port map( A1 => n29245, A2 => n30128, B1 => n29233, B2 => 
                           n31166, ZN => n38174);
   U3602 : AOI22_X1 port map( A1 => n29237, A2 => n31182, B1 => n29236, B2 => 
                           n30127, ZN => n38173);
   U3603 : NAND4_X1 port map( A1 => n38176, A2 => n38175, A3 => n38174, A4 => 
                           n38173, ZN => n38182);
   U3604 : AOI22_X1 port map( A1 => n29114, A2 => n31191, B1 => n29152, B2 => 
                           n30126, ZN => n38180);
   U3605 : AOI22_X1 port map( A1 => n29155, A2 => n31186, B1 => n29021, B2 => 
                           n31193, ZN => n38179);
   U3606 : AOI22_X1 port map( A1 => n29111, A2 => n30125, B1 => n29086, B2 => 
                           n30128, ZN => n38178);
   U3607 : AOI22_X1 port map( A1 => n29150, A2 => n31170, B1 => n29124, B2 => 
                           n31171, ZN => n38177);
   U3608 : NAND4_X1 port map( A1 => n38180, A2 => n38179, A3 => n38178, A4 => 
                           n38177, ZN => n38181);
   U3609 : AOI22_X1 port map( A1 => n38339, A2 => n38182, B1 => n38337, B2 => 
                           n38181, ZN => n38183);
   U3610 : OAI21_X1 port map( B1 => n38342, B2 => n38184, A => n38183, ZN => 
                           OUT1(7));
   U3611 : AOI22_X1 port map( A1 => n29745, A2 => n30054, B1 => n29728, B2 => 
                           n30065, ZN => n38188);
   U3612 : AOI22_X1 port map( A1 => n29726, A2 => n30055, B1 => n29754, B2 => 
                           n31198, ZN => n38187);
   U3613 : AOI22_X1 port map( A1 => n29744, A2 => n30060, B1 => n29022, B2 => 
                           n30061, ZN => n38186);
   U3614 : AOI22_X1 port map( A1 => n29029, A2 => n30053, B1 => n29026, B2 => 
                           n30063, ZN => n38185);
   U3615 : NAND4_X1 port map( A1 => n38188, A2 => n38187, A3 => n38186, A4 => 
                           n38185, ZN => n38194);
   U3616 : AOI22_X1 port map( A1 => n29048, A2 => n31196, B1 => n29044, B2 => 
                           n30056, ZN => n38192);
   U3617 : AOI22_X1 port map( A1 => n29054, A2 => n31177, B1 => n29050, B2 => 
                           n30068, ZN => n38191);
   U3618 : AOI22_X1 port map( A1 => n29051, A2 => n30064, B1 => n29736, B2 => 
                           n30057, ZN => n38190);
   U3619 : AOI22_X1 port map( A1 => n29041, A2 => n30066, B1 => n29049, B2 => 
                           n30067, ZN => n38189);
   U3620 : NAND4_X1 port map( A1 => n38192, A2 => n38191, A3 => n38190, A4 => 
                           n38189, ZN => n38193);
   U3621 : NOR2_X1 port map( A1 => n38194, A2 => n38193, ZN => n38206);
   U3622 : AOI22_X1 port map( A1 => n29813, A2 => n30052, B1 => n29805, B2 => 
                           n31192, ZN => n38198);
   U3623 : AOI22_X1 port map( A1 => n29820, A2 => n30125, B1 => n29819, B2 => 
                           n31191, ZN => n38197);
   U3624 : AOI22_X1 port map( A1 => n29784, A2 => n31186, B1 => n29822, B2 => 
                           n31193, ZN => n38196);
   U3625 : AOI22_X1 port map( A1 => n29818, A2 => n31180, B1 => n29823, B2 => 
                           n31171, ZN => n38195);
   U3626 : NAND4_X1 port map( A1 => n38198, A2 => n38197, A3 => n38196, A4 => 
                           n38195, ZN => n38204);
   U3627 : AOI22_X1 port map( A1 => n29156, A2 => n31186, B1 => n29039, B2 => 
                           n31193, ZN => n38202);
   U3628 : AOI22_X1 port map( A1 => n29115, A2 => n31179, B1 => n29140, B2 => 
                           n31170, ZN => n38201);
   U3629 : AOI22_X1 port map( A1 => n29120, A2 => n31194, B1 => n29105, B2 => 
                           n31187, ZN => n38200);
   U3630 : AOI22_X1 port map( A1 => n29141, A2 => n31167, B1 => n29040, B2 => 
                           n31169, ZN => n38199);
   U3631 : NAND4_X1 port map( A1 => n38202, A2 => n38201, A3 => n38200, A4 => 
                           n38199, ZN => n38203);
   U3632 : AOI22_X1 port map( A1 => n38339, A2 => n38204, B1 => n38337, B2 => 
                           n38203, ZN => n38205);
   U3633 : OAI21_X1 port map( B1 => n38342, B2 => n38206, A => n38205, ZN => 
                           OUT1(6));
   U3634 : AOI22_X1 port map( A1 => n29723, A2 => n30055, B1 => n29057, B2 => 
                           n30063, ZN => n38210);
   U3635 : AOI22_X1 port map( A1 => n29061, A2 => n30061, B1 => n29732, B2 => 
                           n30054, ZN => n38209);
   U3636 : AOI22_X1 port map( A1 => n29071, A2 => n31189, B1 => n29734, B2 => 
                           n30060, ZN => n38208);
   U3637 : AOI22_X1 port map( A1 => n29068, A2 => n31173, B1 => n29052, B2 => 
                           n30064, ZN => n38207);
   U3638 : NAND4_X1 port map( A1 => n38210, A2 => n38209, A3 => n38208, A4 => 
                           n38207, ZN => n38216);
   U3639 : AOI22_X1 port map( A1 => n29069, A2 => n30062, B1 => n29060, B2 => 
                           n31175, ZN => n38214);
   U3640 : AOI22_X1 port map( A1 => n29046, A2 => n30066, B1 => n29751, B2 => 
                           n30059, ZN => n38213);
   U3641 : AOI22_X1 port map( A1 => n29737, A2 => n31181, B1 => n29752, B2 => 
                           n30065, ZN => n38212);
   U3642 : AOI22_X1 port map( A1 => n29058, A2 => n30068, B1 => n29073, B2 => 
                           n30058, ZN => n38211);
   U3643 : NAND4_X1 port map( A1 => n38214, A2 => n38213, A3 => n38212, A4 => 
                           n38211, ZN => n38215);
   U3644 : NOR2_X1 port map( A1 => n38216, A2 => n38215, ZN => n38228);
   U3645 : AOI22_X1 port map( A1 => n29806, A2 => n30126, B1 => n29826, B2 => 
                           n31193, ZN => n38220);
   U3646 : AOI22_X1 port map( A1 => n29827, A2 => n31164, B1 => n29824, B2 => 
                           n31194, ZN => n38219);
   U3647 : AOI22_X1 port map( A1 => n29814, A2 => n31170, B1 => n29825, B2 => 
                           n31179, ZN => n38218);
   U3648 : AOI22_X1 port map( A1 => n29809, A2 => n31186, B1 => n29817, B2 => 
                           n30128, ZN => n38217);
   U3649 : NAND4_X1 port map( A1 => n38220, A2 => n38219, A3 => n38218, A4 => 
                           n38217, ZN => n38226);
   U3650 : AOI22_X1 port map( A1 => n29151, A2 => n31167, B1 => n29110, B2 => 
                           n31160, ZN => n38224);
   U3651 : AOI22_X1 port map( A1 => n29138, A2 => n30051, B1 => n29137, B2 => 
                           n31182, ZN => n38223);
   U3652 : AOI22_X1 port map( A1 => n29109, A2 => n30125, B1 => n29063, B2 => 
                           n31180, ZN => n38222);
   U3653 : AOI22_X1 port map( A1 => n29121, A2 => n31171, B1 => n29065, B2 => 
                           n31193, ZN => n38221);
   U3654 : NAND4_X1 port map( A1 => n38224, A2 => n38223, A3 => n38222, A4 => 
                           n38221, ZN => n38225);
   U3655 : AOI22_X1 port map( A1 => n38339, A2 => n38226, B1 => n38337, B2 => 
                           n38225, ZN => n38227);
   U3656 : OAI21_X1 port map( B1 => n38295, B2 => n38228, A => n38227, ZN => 
                           OUT1(5));
   U3657 : AOI22_X1 port map( A1 => n29056, A2 => n31188, B1 => n29080, B2 => 
                           n31184, ZN => n38232);
   U3658 : AOI22_X1 port map( A1 => n29077, A2 => n31175, B1 => n29101, B2 => 
                           n31173, ZN => n38231);
   U3659 : AOI22_X1 port map( A1 => n29730, A2 => n31185, B1 => n29750, B2 => 
                           n30059, ZN => n38230);
   U3660 : AOI22_X1 port map( A1 => n29729, A2 => n30054, B1 => n29078, B2 => 
                           n31178, ZN => n38229);
   U3661 : NAND4_X1 port map( A1 => n38232, A2 => n38231, A3 => n38230, A4 => 
                           n38229, ZN => n38238);
   U3662 : AOI22_X1 port map( A1 => n29735, A2 => n30060, B1 => n29738, B2 => 
                           n31181, ZN => n38236);
   U3663 : AOI22_X1 port map( A1 => n29100, A2 => n30062, B1 => n29079, B2 => 
                           n30058, ZN => n38235);
   U3664 : AOI22_X1 port map( A1 => n29733, A2 => n30055, B1 => n29096, B2 => 
                           n31189, ZN => n38234);
   U3665 : AOI22_X1 port map( A1 => n29053, A2 => n30064, B1 => n29025, B2 => 
                           n30066, ZN => n38233);
   U3666 : NAND4_X1 port map( A1 => n38236, A2 => n38235, A3 => n38234, A4 => 
                           n38233, ZN => n38237);
   U3667 : NOR2_X1 port map( A1 => n38238, A2 => n38237, ZN => n38250);
   U3668 : AOI22_X1 port map( A1 => n29798, A2 => n30051, B1 => n29791, B2 => 
                           n31167, ZN => n38242);
   U3669 : AOI22_X1 port map( A1 => n29802, A2 => n31187, B1 => n29792, B2 => 
                           n31182, ZN => n38241);
   U3670 : AOI22_X1 port map( A1 => n29771, A2 => n31194, B1 => n29803, B2 => 
                           n31191, ZN => n38240);
   U3671 : AOI22_X1 port map( A1 => n29775, A2 => n31169, B1 => n29785, B2 => 
                           n31159, ZN => n38239);
   U3672 : NAND4_X1 port map( A1 => n38242, A2 => n38241, A3 => n38240, A4 => 
                           n38239, ZN => n38248);
   U3673 : AOI22_X1 port map( A1 => n29117, A2 => n31171, B1 => n29066, B2 => 
                           n31159, ZN => n38246);
   U3674 : AOI22_X1 port map( A1 => n29112, A2 => n31191, B1 => n29153, B2 => 
                           n30126, ZN => n38245);
   U3675 : AOI22_X1 port map( A1 => n29102, A2 => n30125, B1 => n29085, B2 => 
                           n30128, ZN => n38244);
   U3676 : AOI22_X1 port map( A1 => n29144, A2 => n31170, B1 => n29142, B2 => 
                           n30051, ZN => n38243);
   U3677 : NAND4_X1 port map( A1 => n38246, A2 => n38245, A3 => n38244, A4 => 
                           n38243, ZN => n38247);
   U3678 : AOI22_X1 port map( A1 => n38339, A2 => n38248, B1 => n38337, B2 => 
                           n38247, ZN => n38249);
   U3679 : OAI21_X1 port map( B1 => n38342, B2 => n38250, A => n38249, ZN => 
                           OUT1(4));
   U3680 : AOI22_X1 port map( A1 => n29088, A2 => n30053, B1 => n29092, B2 => 
                           n30062, ZN => n38254);
   U3681 : AOI22_X1 port map( A1 => n29740, A2 => n30057, B1 => n29727, B2 => 
                           n30055, ZN => n38253);
   U3682 : AOI22_X1 port map( A1 => n29721, A2 => n30060, B1 => n29082, B2 => 
                           n31184, ZN => n38252);
   U3683 : AOI22_X1 port map( A1 => n29089, A2 => n31178, B1 => n29081, B2 => 
                           n31177, ZN => n38251);
   U3684 : NAND4_X1 port map( A1 => n38254, A2 => n38253, A3 => n38252, A4 => 
                           n38251, ZN => n38260);
   U3685 : AOI22_X1 port map( A1 => n29724, A2 => n31185, B1 => n29055, B2 => 
                           n31188, ZN => n38258);
   U3686 : AOI22_X1 port map( A1 => n29091, A2 => n30067, B1 => n29749, B2 => 
                           n30059, ZN => n38257);
   U3687 : AOI22_X1 port map( A1 => n29755, A2 => n30054, B1 => n29059, B2 => 
                           n31195, ZN => n38256);
   U3688 : AOI22_X1 port map( A1 => n29094, A2 => n31173, B1 => n29027, B2 => 
                           n31183, ZN => n38255);
   U3689 : NAND4_X1 port map( A1 => n38258, A2 => n38257, A3 => n38256, A4 => 
                           n38255, ZN => n38259);
   U3690 : NOR2_X1 port map( A1 => n38260, A2 => n38259, ZN => n38272);
   U3691 : AOI22_X1 port map( A1 => n29793, A2 => n31193, B1 => n29804, B2 => 
                           n31192, ZN => n38264);
   U3692 : AOI22_X1 port map( A1 => n29796, A2 => n31169, B1 => n29787, B2 => 
                           n30051, ZN => n38263);
   U3693 : AOI22_X1 port map( A1 => n29808, A2 => n30127, B1 => n29795, B2 => 
                           n31179, ZN => n38262);
   U3694 : AOI22_X1 port map( A1 => n29794, A2 => n30125, B1 => n29807, B2 => 
                           n30052, ZN => n38261);
   U3695 : NAND4_X1 port map( A1 => n38264, A2 => n38263, A3 => n38262, A4 => 
                           n38261, ZN => n38270);
   U3696 : AOI22_X1 port map( A1 => n29154, A2 => n30051, B1 => n29147, B2 => 
                           n31170, ZN => n38268);
   U3697 : AOI22_X1 port map( A1 => n29158, A2 => n31167, B1 => n29104, B2 => 
                           n31191, ZN => n38267);
   U3698 : AOI22_X1 port map( A1 => n29106, A2 => n31164, B1 => n29067, B2 => 
                           n31193, ZN => n38266);
   U3699 : AOI22_X1 port map( A1 => n29076, A2 => n31169, B1 => n29125, B2 => 
                           n31194, ZN => n38265);
   U3700 : NAND4_X1 port map( A1 => n38268, A2 => n38267, A3 => n38266, A4 => 
                           n38265, ZN => n38269);
   U3701 : AOI22_X1 port map( A1 => n38339, A2 => n38270, B1 => n38337, B2 => 
                           n38269, ZN => n38271);
   U3702 : OAI21_X1 port map( B1 => n38342, B2 => n38272, A => n38271, ZN => 
                           OUT1(3));
   U3703 : AOI22_X1 port map( A1 => n29043, A2 => n31196, B1 => n29045, B2 => 
                           n30061, ZN => n38276);
   U3704 : AOI22_X1 port map( A1 => n29741, A2 => n31197, B1 => n29090, B2 => 
                           n30056, ZN => n38275);
   U3705 : AOI22_X1 port map( A1 => n29036, A2 => n31195, B1 => n29725, B2 => 
                           n30065, ZN => n38274);
   U3706 : AOI22_X1 port map( A1 => n29743, A2 => n31181, B1 => n29030, B2 => 
                           n31184, ZN => n38273);
   U3707 : NAND4_X1 port map( A1 => n38276, A2 => n38275, A3 => n38274, A4 => 
                           n38273, ZN => n38282);
   U3708 : AOI22_X1 port map( A1 => n29720, A2 => n31176, B1 => n29037, B2 => 
                           n30053, ZN => n38280);
   U3709 : AOI22_X1 port map( A1 => n29034, A2 => n30058, B1 => n29731, B2 => 
                           n30055, ZN => n38279);
   U3710 : AOI22_X1 port map( A1 => n29748, A2 => n30059, B1 => n29093, B2 => 
                           n31183, ZN => n38278);
   U3711 : AOI22_X1 port map( A1 => n29042, A2 => n31189, B1 => n29031, B2 => 
                           n30063, ZN => n38277);
   U3712 : NAND4_X1 port map( A1 => n38280, A2 => n38279, A3 => n38278, A4 => 
                           n38277, ZN => n38281);
   U3713 : NOR2_X1 port map( A1 => n38282, A2 => n38281, ZN => n38294);
   U3714 : AOI22_X1 port map( A1 => n29777, A2 => n31190, B1 => n29776, B2 => 
                           n31164, ZN => n38286);
   U3715 : AOI22_X1 port map( A1 => n29800, A2 => n31180, B1 => n29788, B2 => 
                           n31166, ZN => n38285);
   U3716 : AOI22_X1 port map( A1 => n29797, A2 => n31167, B1 => n29789, B2 => 
                           n31182, ZN => n38284);
   U3717 : AOI22_X1 port map( A1 => n29779, A2 => n31171, B1 => n29801, B2 => 
                           n31179, ZN => n38283);
   U3718 : NAND4_X1 port map( A1 => n38286, A2 => n38285, A3 => n38284, A4 => 
                           n38283, ZN => n38292);
   U3719 : AOI22_X1 port map( A1 => n29070, A2 => n31193, B1 => n29123, B2 => 
                           n31171, ZN => n38290);
   U3720 : AOI22_X1 port map( A1 => n29165, A2 => n31192, B1 => n29159, B2 => 
                           n30051, ZN => n38289);
   U3721 : AOI22_X1 port map( A1 => n29075, A2 => n31180, B1 => n29107, B2 => 
                           n31191, ZN => n38288);
   U3722 : AOI22_X1 port map( A1 => n29113, A2 => n30125, B1 => n29166, B2 => 
                           n31182, ZN => n38287);
   U3723 : NAND4_X1 port map( A1 => n38290, A2 => n38289, A3 => n38288, A4 => 
                           n38287, ZN => n38291);
   U3724 : AOI22_X1 port map( A1 => n38339, A2 => n38292, B1 => n38337, B2 => 
                           n38291, ZN => n38293);
   U3725 : OAI21_X1 port map( B1 => n38295, B2 => n38294, A => n38293, ZN => 
                           OUT1(2));
   U3726 : AOI22_X1 port map( A1 => n29722, A2 => n30055, B1 => n29099, B2 => 
                           n31183, ZN => n38299);
   U3727 : AOI22_X1 port map( A1 => n29742, A2 => n31197, B1 => n29097, B2 => 
                           n30062, ZN => n38298);
   U3728 : AOI22_X1 port map( A1 => n29064, A2 => n30064, B1 => n29746, B2 => 
                           n31198, ZN => n38297);
   U3729 : AOI22_X1 port map( A1 => n29095, A2 => n30067, B1 => n29083, B2 => 
                           n31177, ZN => n38296);
   U3730 : NAND4_X1 port map( A1 => n38299, A2 => n38298, A3 => n38297, A4 => 
                           n38296, ZN => n38305);
   U3731 : AOI22_X1 port map( A1 => n29739, A2 => n30060, B1 => n29098, B2 => 
                           n30056, ZN => n38303);
   U3732 : AOI22_X1 port map( A1 => n29087, A2 => n31175, B1 => n29062, B2 => 
                           n30061, ZN => n38302);
   U3733 : AOI22_X1 port map( A1 => n29084, A2 => n31184, B1 => n29753, B2 => 
                           n30057, ZN => n38301);
   U3734 : AOI22_X1 port map( A1 => n29032, A2 => n30063, B1 => n29747, B2 => 
                           n30065, ZN => n38300);
   U3735 : NAND4_X1 port map( A1 => n38303, A2 => n38302, A3 => n38301, A4 => 
                           n38300, ZN => n38304);
   U3736 : NOR2_X1 port map( A1 => n38305, A2 => n38304, ZN => n38317);
   U3737 : AOI22_X1 port map( A1 => n29783, A2 => n31193, B1 => n29767, B2 => 
                           n31186, ZN => n38309);
   U3738 : AOI22_X1 port map( A1 => n29790, A2 => n31191, B1 => n29781, B2 => 
                           n30052, ZN => n38308);
   U3739 : AOI22_X1 port map( A1 => n29773, A2 => n31169, B1 => n29782, B2 => 
                           n30127, ZN => n38307);
   U3740 : AOI22_X1 port map( A1 => n29780, A2 => n31167, B1 => n29786, B2 => 
                           n30125, ZN => n38306);
   U3741 : NAND4_X1 port map( A1 => n38309, A2 => n38308, A3 => n38307, A4 => 
                           n38306, ZN => n38315);
   U3742 : AOI22_X1 port map( A1 => n29116, A2 => n31194, B1 => n29149, B2 => 
                           n31166, ZN => n38313);
   U3743 : AOI22_X1 port map( A1 => n29108, A2 => n31191, B1 => n29143, B2 => 
                           n30126, ZN => n38312);
   U3744 : AOI22_X1 port map( A1 => n29072, A2 => n31159, B1 => n29139, B2 => 
                           n31182, ZN => n38311);
   U3745 : AOI22_X1 port map( A1 => n29074, A2 => n31169, B1 => n29103, B2 => 
                           n30125, ZN => n38310);
   U3746 : NAND4_X1 port map( A1 => n38313, A2 => n38312, A3 => n38311, A4 => 
                           n38310, ZN => n38314);
   U3747 : AOI22_X1 port map( A1 => n38339, A2 => n38315, B1 => n38337, B2 => 
                           n38314, ZN => n38316);
   U3748 : OAI21_X1 port map( B1 => n38342, B2 => n38317, A => n38316, ZN => 
                           OUT1(1));
   U3749 : AOI22_X1 port map( A1 => n29833, A2 => n31185, B1 => n29127, B2 => 
                           n30068, ZN => n38321);
   U3750 : AOI22_X1 port map( A1 => n29130, A2 => n31178, B1 => n29135, B2 => 
                           n30063, ZN => n38320);
   U3751 : AOI22_X1 port map( A1 => n29131, A2 => n30066, B1 => n29215, B2 => 
                           n30056, ZN => n38319);
   U3752 : AOI22_X1 port map( A1 => n29829, A2 => n30059, B1 => n29832, B2 => 
                           n31181, ZN => n38318);
   U3753 : NAND4_X1 port map( A1 => n38321, A2 => n38320, A3 => n38319, A4 => 
                           n38318, ZN => n38327);
   U3754 : AOI22_X1 port map( A1 => n29128, A2 => n31175, B1 => n29126, B2 => 
                           n31177, ZN => n38325);
   U3755 : AOI22_X1 port map( A1 => n29136, A2 => n30062, B1 => n29831, B2 => 
                           n31197, ZN => n38324);
   U3756 : AOI22_X1 port map( A1 => n29830, A2 => n31174, B1 => n29828, B2 => 
                           n30060, ZN => n38323);
   U3757 : AOI22_X1 port map( A1 => n29201, A2 => n31189, B1 => n29132, B2 => 
                           n30064, ZN => n38322);
   U3758 : NAND4_X1 port map( A1 => n38325, A2 => n38324, A3 => n38323, A4 => 
                           n38322, ZN => n38326);
   U3759 : NOR2_X1 port map( A1 => n38327, A2 => n38326, ZN => n38341);
   U3760 : AOI22_X1 port map( A1 => n29757, A2 => n31193, B1 => n29758, B2 => 
                           n30125, ZN => n38331);
   U3761 : AOI22_X1 port map( A1 => n29759, A2 => n31194, B1 => n29761, B2 => 
                           n30051, ZN => n38330);
   U3762 : AOI22_X1 port map( A1 => n29756, A2 => n31180, B1 => n29760, B2 => 
                           n31167, ZN => n38329);
   U3763 : AOI22_X1 port map( A1 => n29762, A2 => n31191, B1 => n29763, B2 => 
                           n31182, ZN => n38328);
   U3764 : NAND4_X1 port map( A1 => n38331, A2 => n38330, A3 => n38329, A4 => 
                           n38328, ZN => n38338);
   U3765 : AOI22_X1 port map( A1 => n29134, A2 => n30125, B1 => n29260, B2 => 
                           n31166, ZN => n38335);
   U3766 : AOI22_X1 port map( A1 => n29262, A2 => n31167, B1 => n29210, B2 => 
                           n30128, ZN => n38334);
   U3767 : AOI22_X1 port map( A1 => n29133, A2 => n31193, B1 => n29261, B2 => 
                           n31170, ZN => n38333);
   U3768 : AOI22_X1 port map( A1 => n29248, A2 => n30127, B1 => n29129, B2 => 
                           n31160, ZN => n38332);
   U3769 : NAND4_X1 port map( A1 => n38335, A2 => n38334, A3 => n38333, A4 => 
                           n38332, ZN => n38336);
   U3770 : AOI22_X1 port map( A1 => n38339, A2 => n38338, B1 => n38337, B2 => 
                           n38336, ZN => n38340);
   U3771 : OAI21_X1 port map( B1 => n38342, B2 => n38341, A => n38340, ZN => 
                           OUT1(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_17_port, curr_instruction_to_cu_i_16_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n151, cu_i_n135, 
      cu_i_N279, cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, 
      cu_i_N273, cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, 
      cu_i_cmd_alu_op_type_0_port, cu_i_cmd_alu_op_type_1_port, 
      cu_i_cmd_alu_op_type_2_port, cu_i_cmd_alu_op_type_3_port, 
      cu_i_cmd_word_3_port, cu_i_cmd_word_6_port, cu_i_cmd_word_8_port, 
      datapath_i_alu_output_val_i_0_port, datapath_i_alu_output_val_i_1_port, 
      datapath_i_alu_output_val_i_2_port, datapath_i_alu_output_val_i_3_port, 
      datapath_i_alu_output_val_i_4_port, datapath_i_alu_output_val_i_5_port, 
      datapath_i_alu_output_val_i_6_port, datapath_i_alu_output_val_i_7_port, 
      datapath_i_alu_output_val_i_8_port, datapath_i_alu_output_val_i_9_port, 
      datapath_i_alu_output_val_i_10_port, datapath_i_alu_output_val_i_11_port,
      datapath_i_alu_output_val_i_12_port, datapath_i_alu_output_val_i_13_port,
      datapath_i_alu_output_val_i_14_port, datapath_i_alu_output_val_i_15_port,
      datapath_i_alu_output_val_i_16_port, datapath_i_alu_output_val_i_17_port,
      datapath_i_alu_output_val_i_18_port, datapath_i_alu_output_val_i_19_port,
      datapath_i_alu_output_val_i_20_port, datapath_i_alu_output_val_i_21_port,
      datapath_i_alu_output_val_i_22_port, datapath_i_alu_output_val_i_23_port,
      datapath_i_alu_output_val_i_24_port, datapath_i_alu_output_val_i_25_port,
      datapath_i_alu_output_val_i_26_port, datapath_i_alu_output_val_i_27_port,
      datapath_i_alu_output_val_i_28_port, datapath_i_alu_output_val_i_29_port,
      datapath_i_alu_output_val_i_30_port, datapath_i_alu_output_val_i_31_port,
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_decode_stage_dp_n44, datapath_i_decode_stage_dp_n43, 
      datapath_i_decode_stage_dp_n42, datapath_i_decode_stage_dp_n41, 
      datapath_i_decode_stage_dp_n40, datapath_i_decode_stage_dp_n39, 
      datapath_i_decode_stage_dp_n38, datapath_i_decode_stage_dp_n37, 
      datapath_i_decode_stage_dp_n36, datapath_i_decode_stage_dp_n35, 
      datapath_i_decode_stage_dp_n34, datapath_i_decode_stage_dp_n33, 
      datapath_i_decode_stage_dp_n32, datapath_i_decode_stage_dp_n31, 
      datapath_i_decode_stage_dp_n30, datapath_i_decode_stage_dp_n29, 
      datapath_i_decode_stage_dp_n28, datapath_i_decode_stage_dp_n27, 
      datapath_i_decode_stage_dp_n26, datapath_i_decode_stage_dp_n25, 
      datapath_i_decode_stage_dp_n24, datapath_i_decode_stage_dp_n23, 
      datapath_i_decode_stage_dp_n22, datapath_i_decode_stage_dp_n21, 
      datapath_i_decode_stage_dp_n20, datapath_i_decode_stage_dp_n19, 
      datapath_i_decode_stage_dp_n18, datapath_i_decode_stage_dp_n17, 
      datapath_i_decode_stage_dp_n16, datapath_i_decode_stage_dp_n15, 
      datapath_i_decode_stage_dp_n14, datapath_i_decode_stage_dp_n13, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, n301, n302, n474, n477, n492, 
      n1427, n1429, n1431, n1433, n1435, n1437, n1439, n1441, n1443, n1445, 
      n1447, n1449, n1453, n1613, n1614, n1615, n1617, n1619, n1621, n1623, 
      n1625, n1627, n1629, n1631, n1633, n1635, n1637, n1639, n1641, n1643, 
      n1645, n1647, n1649, n1651, n1653, n1655, n1657, n1659, n1661, n1663, 
      n1665, n1667, n1669, n1671, n1673, n2299, n3112, n3119, n3120, n3121, 
      n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
      n3132, n3133, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3155, n3160, n3161, n5478, 
      n5479, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, 
      n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
      n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
      n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
      n3205, n3206, n3207, n3209, n3210, n3211, n3227, n3229, n3231, n3233, 
      n3235, n3236, n3238, n3239, n3241, n3242, n3243, n3248, n3252, n3254, 
      n3257, n3261, n3269, n3281, n3284, n3288, n3291, n3294, n3297, n3300, 
      n3303, n3306, n3309, n3312, n3315, n3318, n3321, n3324, n3327, n3330, 
      n3333, n3336, n3339, n3342, n3345, n3348, n3351, n3354, n3357, n3360, 
      n3363, n3366, n3369, n3372, n3375, n3378, n3381, n3543, n3555, n3692, 
      n3596, n4048, n4052, n4060, n4128, n4133, n4155, n4187, n4193, n4228, 
      n4230, n4231, n4268, n4280, n4337, n4341, n4344, n4417, n5542, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4992, n4993, 
      n4995, IRAM_ADDRESS_29_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_25_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_13_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_11_port, n5006, n5007, n6233, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n6232, IRAM_ADDRESS_6_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_2_port, n5065, n5066, n5067, n5068, 
      n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, 
      n5079, n5081, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, 
      n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, 
      n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, 
      n5113, n5115, n5116, n5117, n5119, n5120, n5121, n5122, n5123, n5125, 
      n5126, n5127, n5128, n5129, n5130, n5131, n5134, n5135, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, 
      n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, 
      n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, 
      n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, 
      n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, 
      n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, 
      n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, 
      n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, 
      n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, 
      n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, 
      n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, 
      n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, 
      n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, 
      n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, 
      n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5288, 
      n5290, n5291, n5293, n5294, n5296, n5297, n5299, n5300, n5302, n5303, 
      n5305, n5306, n5308, n5309, n5311, n5312, n5314, n5315, n5317, n5319, 
      n5320, n5322, n5323, n5324, n5325, n5326, n5328, n5329, n5330, n5331, 
      n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, 
      n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, 
      n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, 
      n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, 
      n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, 
      n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5392, 
      IRAM_ADDRESS_12_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_8_port, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5442, n5443, n5444, n5445, n5448, 
      n5449, n5450, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, 
      n5461, n5462, n5463, n5465, n5481, n5482, n5483, n5484, n5485, n5486, 
      n5487, n5488, n5489, n5501, n5502, n5503, n5504, n5505, n5506, n5507, 
      n5508, n5509, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, 
      n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, 
      n5529, n5530, n5531, n5532, n5534, n5537, n5538, n5539, n5540, n5541, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5860, n5861, n5862, n5863, n5864, n5865, 
      n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, 
      n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, 
      n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, 
      n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, 
      n5906, n5907, n5908, IRAM_ADDRESS_14_port, IRAM_ADDRESS_16_port, 
      IRAM_ADDRESS_18_port, IRAM_ADDRESS_20_port, IRAM_ADDRESS_22_port, 
      IRAM_ADDRESS_24_port, IRAM_ADDRESS_26_port, IRAM_ADDRESS_28_port, 
      IRAM_ADDRESS_30_port, n5918, n5919, n5920, n5921, n5922, n5923, n5924, 
      n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, 
      n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, 
      n5945, n5946, n5947, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, 
      IRAM_ADDRESS_31_port, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, 
      n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
      n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, 
      n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, 
      n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, 
      n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, 
      n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
      n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
      n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
      n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, 
      n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, 
      n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6230, n6231, n_3831, n_3832, n_3833, n_3834, n_3835, 
      n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, 
      n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, 
      n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, 
      n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, 
      n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, 
      n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, 
      n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, 
      n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, 
      n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, 
      n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, 
      n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, 
      n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, 
      n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, 
      n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, 
      n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, 
      n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, 
      n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, 
      n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, 
      n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, 
      n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, 
      n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, 
      n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033, 
      n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, 
      n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, 
      n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, 
      n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, 
      n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, 
      n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, 
      n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, 
      n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, 
      n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, 
      n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, 
      n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, 
      n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, 
      n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, 
      n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, 
      n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, 
      n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177, 
      n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, 
      n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, 
      n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, 
      n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, 
      n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, 
      n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, 
      n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, 
      n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, 
      n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, 
      n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, 
      n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, 
      n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, 
      n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, 
      n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, 
      n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, 
      n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, 
      n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330 : 
      std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => n3284);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => n4417);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_n151);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => n3281);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n5358, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n5406, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n5406, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n5406, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n5406, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n5406, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n5406, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n5406, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n5406, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n5406, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n5406, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n5406, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n4993, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n4993, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n4993, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n4993, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n4993, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n5406, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n5358, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n5358, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n5358, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n5358, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n5358, Z 
                           => DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n5358, Z 
                           => DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n5358, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n5358, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n5358, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n5358, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n5358, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n5358, Z 
                           => DRAM_ADDRESS_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n301, D => n5078, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n301, D => n5458, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n301, D => n5457, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n301, D => n5077, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n301, D => n5076, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n301, D => n5449, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n301, D => n5041, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n301, D => n5042, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n301, D => n5043, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n301, D => n5044, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n301, D => n5045, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n301, D => n5071, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n301, D => n5065, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n301, D => n5459, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n301, D => n5067, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n301, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n5882, D => n5078, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n5882, D => n5458, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n5882, D => n5457, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n5882, D => n5077, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n5882, D => n5076, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n5882, D => n5449, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n5882, D => n5041, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n5882, D => n5042, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n5882, D => n5043, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n5882, D => n5044, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n5882, D => n5045, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n5882, D => n5071, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n5882, D => n5065, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n6229, D => n5459, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n5882, D => n5067, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n5882, D => n5069, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n5882, D => n5072, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n6229, D => n5066, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n5882, D => n5453, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n6229, D => n5068, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n5882, D => n5070, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n6229, D => n5046, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n5882, D => n5047, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n5882, D => n5079, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n6229, D => n5048, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n5882, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n6229, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n6229, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n6229, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n5882, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n6229, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n5882, D => n5049, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   clk_r_REG10041_S2 : DFFR_X1 port map( D => n6229, CK => CLK, RN => RST, Q =>
                           n5462, QN => n_3831);
   clk_r_REG10127_S6 : DFFR_X1 port map( D => n3555, CK => CLK, RN => RST, Q =>
                           n_3832, QN => n5461);
   clk_r_REG10092_S3 : DFFR_X1 port map( D => n4133, CK => CLK, RN => RST, Q =>
                           n_3833, QN => n5460);
   clk_r_REG10255_S7 : DFFR_X1 port map( D => n5877, CK => CLK, RN => RST, Q =>
                           n5459, QN => n_3834);
   clk_r_REG10263_S7 : DFFR_X1 port map( D => n5878, CK => CLK, RN => RST, Q =>
                           n5458, QN => n5532);
   clk_r_REG10265_S7 : DFFR_X1 port map( D => n5879, CK => CLK, RN => RST, Q =>
                           n5457, QN => n5509);
   clk_r_REG10268_S7 : DFFR_X1 port map( D => n5884, CK => CLK, RN => RST, Q =>
                           n5456, QN => n_3835);
   clk_r_REG10273_S7 : DFFR_X1 port map( D => n5886, CK => CLK, RN => RST, Q =>
                           n5455, QN => n_3836);
   clk_r_REG10272_S1 : DFFR_X1 port map( D => n5883, CK => CLK, RN => RST, Q =>
                           n5454, QN => n_3837);
   clk_r_REG10256_S7 : DFFR_X1 port map( D => n5876, CK => CLK, RN => RST, Q =>
                           n5453, QN => n_3838);
   clk_r_REG10274_S7 : DFFR_X1 port map( D => n5887, CK => CLK, RN => RST, Q =>
                           n6226, QN => n5537);
   clk_r_REG10276_S7 : DFFR_X1 port map( D => n5888, CK => CLK, RN => RST, Q =>
                           n_3839, QN => n5538);
   clk_r_REG10300_S1 : DFFR_X1 port map( D => n5890, CK => CLK, RN => RST, Q =>
                           n5450, QN => n_3840);
   clk_r_REG10279_S7 : DFFR_X1 port map( D => n5891, CK => CLK, RN => RST, Q =>
                           n5449, QN => n_3841);
   clk_r_REG10278_S7 : DFFR_X1 port map( D => n5892, CK => CLK, RN => RST, Q =>
                           n5448, QN => n_3842);
   clk_r_REG10118_S2 : DFFR_X1 port map( D => n5873, CK => CLK, RN => RST, Q =>
                           DRAM_READNOTWRITE, QN => n_3843);
   clk_r_REG10111_S2 : DFFS_X1 port map( D => n3543, CK => CLK, SN => RST, Q =>
                           n_3844, QN => DRAM_ENABLE);
   clk_r_REG8055_S7 : DFFS_X1 port map( D => n5908, CK => CLK, SN => RST, Q => 
                           n5445, QN => n_3845);
   clk_r_REG8158_S8 : DFFS_X1 port map( D => n5445, CK => CLK, SN => RST, Q => 
                           n5444, QN => n_3846);
   clk_r_REG8061_S6 : DFFS_X1 port map( D => n5907, CK => CLK, SN => RST, Q => 
                           n5443, QN => n_3847);
   clk_r_REG8151_S7 : DFFS_X1 port map( D => n5443, CK => CLK, SN => RST, Q => 
                           n5442, QN => n_3848);
   clk_r_REG10123_S4 : DFFS_X1 port map( D => n5867, CK => CLK, SN => RST, Q =>
                           n_3849, QN => n5540);
   clk_r_REG10040_S2 : DFFR_X1 port map( D => n6229, CK => CLK, RN => RST, Q =>
                           n5440, QN => n6217);
   clk_r_REG10063_S3 : DFFR_X1 port map( D => n5440, CK => CLK, RN => RST, Q =>
                           n5439, QN => n_3850);
   clk_r_REG10053_S2 : DFFR_X1 port map( D => n5864, CK => CLK, RN => RST, Q =>
                           n5438, QN => n_3851);
   clk_r_REG10054_S2 : DFFR_X1 port map( D => n5863, CK => CLK, RN => RST, Q =>
                           n5437, QN => n_3852);
   clk_r_REG10058_S2 : DFFR_X1 port map( D => n5862, CK => CLK, RN => RST, Q =>
                           n5436, QN => n_3853);
   clk_r_REG10062_S2 : DFFR_X1 port map( D => n5861, CK => CLK, RN => RST, Q =>
                           n5435, QN => n_3854);
   clk_r_REG8043_S7 : DFFS_X1 port map( D => n5945, CK => CLK, SN => RST, Q => 
                           n5434, QN => n_3855);
   clk_r_REG8182_S8 : DFFS_X1 port map( D => n5434, CK => CLK, SN => RST, Q => 
                           n5433, QN => n_3856);
   clk_r_REG8047_S7 : DFFS_X1 port map( D => n5906, CK => CLK, SN => RST, Q => 
                           n5432, QN => n_3857);
   clk_r_REG8166_S8 : DFFS_X1 port map( D => n5432, CK => CLK, SN => RST, Q => 
                           n5431, QN => n_3858);
   clk_r_REG8067_S6 : DFFS_X1 port map( D => n5905, CK => CLK, SN => RST, Q => 
                           n5430, QN => n_3859);
   clk_r_REG8143_S7 : DFFS_X1 port map( D => n5430, CK => CLK, SN => RST, Q => 
                           n5429, QN => n_3860);
   clk_r_REG10101_S1 : DFFR_X1 port map( D => n301, CK => CLK, RN => RST, Q => 
                           n5428, QN => n_3861);
   clk_r_REG8074_S6 : DFFS_X1 port map( D => n5904, CK => CLK, SN => RST, Q => 
                           n5427, QN => n_3862);
   clk_r_REG8136_S7 : DFFS_X1 port map( D => n5427, CK => CLK, SN => RST, Q => 
                           n5426, QN => n_3863);
   clk_r_REG7506_S6 : DFFS_X1 port map( D => n5893, CK => CLK, SN => RST, Q => 
                           n5425, QN => n_3864);
   clk_r_REG7507_S7 : DFFS_X1 port map( D => n5425, CK => CLK, SN => RST, Q => 
                           n5424, QN => n_3865);
   clk_r_REG7508_S8 : DFFS_X1 port map( D => n5424, CK => CLK, SN => RST, Q => 
                           n5423, QN => n_3866);
   clk_r_REG8027_S7 : DFFS_X1 port map( D => n5894, CK => CLK, SN => RST, Q => 
                           n5422, QN => n_3867);
   clk_r_REG8028_S8 : DFFS_X1 port map( D => n5422, CK => CLK, SN => RST, Q => 
                           n5421, QN => n_3868);
   clk_r_REG8184_S9 : DFFS_X1 port map( D => n5421, CK => CLK, SN => RST, Q => 
                           n5420, QN => n_3869);
   clk_r_REG8080_S6 : DFFS_X1 port map( D => n5903, CK => CLK, SN => RST, Q => 
                           n5419, QN => n_3870);
   clk_r_REG8129_S7 : DFFS_X1 port map( D => n5419, CK => CLK, SN => RST, Q => 
                           n5418, QN => n_3871);
   clk_r_REG8086_S6 : DFFS_X1 port map( D => n5902, CK => CLK, SN => RST, Q => 
                           n5417, QN => n_3872);
   clk_r_REG8121_S7 : DFFS_X1 port map( D => n5417, CK => CLK, SN => RST, Q => 
                           n5416, QN => n_3873);
   clk_r_REG8092_S6 : DFFS_X1 port map( D => n5901, CK => CLK, SN => RST, Q => 
                           n5415, QN => n_3874);
   clk_r_REG8114_S7 : DFFS_X1 port map( D => n5415, CK => CLK, SN => RST, Q => 
                           n5414, QN => n_3875);
   clk_r_REG8098_S6 : DFFS_X1 port map( D => n5900, CK => CLK, SN => RST, Q => 
                           n5413, QN => n_3876);
   clk_r_REG8107_S7 : DFFS_X1 port map( D => n5413, CK => CLK, SN => RST, Q => 
                           n5412, QN => n_3877);
   clk_r_REG8100_S6 : DFFS_X1 port map( D => n5899, CK => CLK, SN => RST, Q => 
                           n5411, QN => n_3878);
   clk_r_REG8104_S7 : DFFS_X1 port map( D => n5411, CK => CLK, SN => RST, Q => 
                           n5410, QN => n_3879);
   clk_r_REG9914_S5 : DFFR_X1 port map( D => n5408, CK => CLK, RN => RST, Q => 
                           n5407, QN => n_3880);
   clk_r_REG10115_S2 : DFFS_X1 port map( D => n3543, CK => CLK, SN => RST, Q =>
                           n5406, QN => n_3881);
   clk_r_REG10113_S2 : DFFS_X1 port map( D => n3254, CK => CLK, SN => RST, Q =>
                           n5405, QN => n_3882);
   clk_r_REG8185_S5 : DFFR_X1 port map( D => n1449, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_8_port, QN => n_3883);
   clk_r_REG8183_S5 : DFFR_X1 port map( D => n1447, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_10_port, QN => n_3884);
   clk_r_REG8181_S5 : DFFR_X1 port map( D => n1445, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_12_port, QN => n_3885);
   clk_r_REG8165_S5 : DFFR_X1 port map( D => n1443, CK => CLK, RN => RST, Q => 
                           n_3886, QN => n5484);
   clk_r_REG8157_S5 : DFFR_X1 port map( D => n1441, CK => CLK, RN => RST, Q => 
                           n_3887, QN => n5485);
   clk_r_REG8150_S5 : DFFR_X1 port map( D => n1439, CK => CLK, RN => RST, Q => 
                           n_3888, QN => n5486);
   clk_r_REG8142_S5 : DFFR_X1 port map( D => n1437, CK => CLK, RN => RST, Q => 
                           n_3889, QN => n5483);
   clk_r_REG8135_S5 : DFFR_X1 port map( D => n1435, CK => CLK, RN => RST, Q => 
                           n_3890, QN => n5481);
   clk_r_REG8128_S5 : DFFR_X1 port map( D => n1433, CK => CLK, RN => RST, Q => 
                           n_3891, QN => n5487);
   clk_r_REG8120_S5 : DFFR_X1 port map( D => n1431, CK => CLK, RN => RST, Q => 
                           n_3892, QN => n5488);
   clk_r_REG8113_S5 : DFFR_X1 port map( D => n1429, CK => CLK, RN => RST, Q => 
                           n_3893, QN => n5489);
   clk_r_REG8106_S5 : DFFR_X1 port map( D => n1427, CK => CLK, RN => RST, Q => 
                           n_3894, QN => n5482);
   clk_r_REG10087_S4 : DFFR_X1 port map( D => n3241, CK => CLK, RN => RST, Q =>
                           n5392, QN => n_3895);
   clk_r_REG7948_S7 : DFFR_X1 port map( D => n5531, CK => CLK, RN => RST, Q => 
                           n6221, QN => n5503);
   clk_r_REG8037_S8 : DFFS_X1 port map( D => n5529, CK => CLK, SN => RST, Q => 
                           n5390, QN => n_3896);
   clk_r_REG9917_S4 : DFFS_X1 port map( D => n5528, CK => CLK, SN => RST, Q => 
                           n5389, QN => n_3897);
   clk_r_REG9913_S5 : DFFS_X1 port map( D => n5385, CK => CLK, SN => RST, Q => 
                           n5384, QN => n_3898);
   clk_r_REG9907_S4 : DFFR_X1 port map( D => n5516, CK => CLK, RN => RST, Q => 
                           n5383, QN => n6215);
   clk_r_REG9910_S4 : DFFS_X1 port map( D => n5515, CK => CLK, SN => RST, Q => 
                           n5382, QN => n6216);
   clk_r_REG8096_S6 : DFFR_X1 port map( D => n5939, CK => CLK, RN => RST, Q => 
                           n5381, QN => n_3899);
   clk_r_REG8097_S6 : DFFS_X1 port map( D => n5939, CK => CLK, SN => RST, Q => 
                           n5380, QN => n_3900);
   clk_r_REG8090_S6 : DFFR_X1 port map( D => n5937, CK => CLK, RN => RST, Q => 
                           n5379, QN => n_3901);
   clk_r_REG8091_S6 : DFFS_X1 port map( D => n5937, CK => CLK, SN => RST, Q => 
                           n5378, QN => n_3902);
   clk_r_REG8084_S6 : DFFR_X1 port map( D => n5935, CK => CLK, RN => RST, Q => 
                           n5377, QN => n_3903);
   clk_r_REG8085_S6 : DFFS_X1 port map( D => n5935, CK => CLK, SN => RST, Q => 
                           n5376, QN => n_3904);
   clk_r_REG8078_S6 : DFFR_X1 port map( D => n5933, CK => CLK, RN => RST, Q => 
                           n5375, QN => n_3905);
   clk_r_REG8079_S6 : DFFS_X1 port map( D => n5933, CK => CLK, SN => RST, Q => 
                           n5374, QN => n_3906);
   clk_r_REG8052_S6 : DFFR_X1 port map( D => n5925, CK => CLK, RN => RST, Q => 
                           n5373, QN => n_3907);
   clk_r_REG8053_S6 : DFFS_X1 port map( D => n5925, CK => CLK, SN => RST, Q => 
                           n5372, QN => n_3908);
   clk_r_REG8170_S7 : DFFR_X1 port map( D => n5923, CK => CLK, RN => RST, Q => 
                           n5371, QN => n_3909);
   clk_r_REG8171_S7 : DFFS_X1 port map( D => n5923, CK => CLK, SN => RST, Q => 
                           n5370, QN => n_3910);
   clk_r_REG8059_S6 : DFFR_X1 port map( D => n5927, CK => CLK, RN => RST, Q => 
                           n5369, QN => n_3911);
   clk_r_REG8060_S6 : DFFS_X1 port map( D => n5927, CK => CLK, SN => RST, Q => 
                           n5368, QN => n_3912);
   clk_r_REG8065_S6 : DFFR_X1 port map( D => n5929, CK => CLK, RN => RST, Q => 
                           n5367, QN => n_3913);
   clk_r_REG8066_S6 : DFFS_X1 port map( D => n5929, CK => CLK, SN => RST, Q => 
                           n5366, QN => n_3914);
   clk_r_REG8071_S6 : DFFR_X1 port map( D => n5931, CK => CLK, RN => RST, Q => 
                           n5365, QN => n_3915);
   clk_r_REG8072_S6 : DFFS_X1 port map( D => n5931, CK => CLK, SN => RST, Q => 
                           n5364, QN => n_3916);
   clk_r_REG9892_S5 : DFFS_X1 port map( D => n5896, CK => CLK, SN => RST, Q => 
                           n5363, QN => n_3917);
   clk_r_REG9893_S6 : DFFS_X1 port map( D => n5363, CK => CLK, SN => RST, Q => 
                           n5362, QN => n_3918);
   clk_r_REG9894_S7 : DFFS_X1 port map( D => n5362, CK => CLK, SN => RST, Q => 
                           n5361, QN => n_3919);
   clk_r_REG9908_S3 : DFFR_X1 port map( D => n5870, CK => CLK, RN => RST, Q => 
                           n5360, QN => n5515);
   clk_r_REG9909_S4 : DFFS_X1 port map( D => n5515, CK => CLK, SN => RST, Q => 
                           n_3920, QN => n5359);
   clk_r_REG10114_S2 : DFFS_X1 port map( D => n3543, CK => CLK, SN => RST, Q =>
                           n5358, QN => n_3921);
   clk_r_REG8418_S5 : DFFS_X1 port map( D => n5919, CK => CLK, SN => RST, Q => 
                           n5357, QN => n_3922);
   clk_r_REG8419_S6 : DFFS_X1 port map( D => n5357, CK => CLK, SN => RST, Q => 
                           n5356, QN => n_3923);
   clk_r_REG8420_S7 : DFFS_X1 port map( D => n5356, CK => CLK, SN => RST, Q => 
                           n5355, QN => n_3924);
   clk_r_REG9898_S5 : DFFS_X1 port map( D => n5918, CK => CLK, SN => RST, Q => 
                           n5354, QN => n_3925);
   clk_r_REG9899_S6 : DFFS_X1 port map( D => n5354, CK => CLK, SN => RST, Q => 
                           n5353, QN => n_3926);
   clk_r_REG9900_S7 : DFFS_X1 port map( D => n5353, CK => CLK, SN => RST, Q => 
                           n5352, QN => n_3927);
   clk_r_REG10097_S3 : DFFS_X1 port map( D => n5875, CK => CLK, SN => RST, Q =>
                           n5351, QN => n_3928);
   clk_r_REG10093_S3 : DFFR_X1 port map( D => n4133, CK => CLK, RN => RST, Q =>
                           n5350, QN => n_3929);
   clk_r_REG8099_S5 : DFFR_X1 port map( D => n1427, CK => CLK, RN => RST, Q => 
                           n5349, QN => n_3930);
   clk_r_REG8093_S5 : DFFR_X1 port map( D => n1429, CK => CLK, RN => RST, Q => 
                           n5348, QN => n_3931);
   clk_r_REG8087_S5 : DFFR_X1 port map( D => n1431, CK => CLK, RN => RST, Q => 
                           n5347, QN => n_3932);
   clk_r_REG8081_S5 : DFFR_X1 port map( D => n1433, CK => CLK, RN => RST, Q => 
                           n5346, QN => n_3933);
   clk_r_REG8075_S5 : DFFR_X1 port map( D => n1435, CK => CLK, RN => RST, Q => 
                           n5345, QN => n_3934);
   clk_r_REG8068_S5 : DFFR_X1 port map( D => n1437, CK => CLK, RN => RST, Q => 
                           n5344, QN => n_3935);
   clk_r_REG8062_S5 : DFFR_X1 port map( D => n1439, CK => CLK, RN => RST, Q => 
                           n5343, QN => n_3936);
   clk_r_REG8056_S5 : DFFR_X1 port map( D => n1441, CK => CLK, RN => RST, Q => 
                           n5342, QN => n_3937);
   clk_r_REG8048_S5 : DFFR_X1 port map( D => n1443, CK => CLK, RN => RST, Q => 
                           n5341, QN => n_3938);
   clk_r_REG10281_S7 : DFFS_X1 port map( D => n5944, CK => CLK, SN => RST, Q =>
                           n5340, QN => n6222);
   clk_r_REG6931_S5 : DFFS_X1 port map( D => n5895, CK => CLK, SN => RST, Q => 
                           n5339, QN => n_3939);
   clk_r_REG6932_S6 : DFFS_X1 port map( D => n5339, CK => CLK, SN => RST, Q => 
                           n5338, QN => n_3940);
   clk_r_REG6933_S7 : DFFS_X1 port map( D => n5338, CK => CLK, SN => RST, Q => 
                           n5337, QN => n_3941);
   clk_r_REG10016_S1 : DFFS_X1 port map( D => n5512, CK => CLK, SN => RST, Q =>
                           n5336, QN => n_3942);
   clk_r_REG6926_S3 : DFFR_X1 port map( D => n5505, CK => CLK, RN => RST, Q => 
                           n5335, QN => n5514);
   clk_r_REG6927_S4 : DFFS_X1 port map( D => n5514, CK => CLK, SN => RST, Q => 
                           n_3943, QN => n5334);
   clk_r_REG7724_S6 : DFFS_X1 port map( D => n5897, CK => CLK, SN => RST, Q => 
                           n5333, QN => n_3944);
   clk_r_REG7725_S7 : DFFS_X1 port map( D => n5333, CK => CLK, SN => RST, Q => 
                           n5332, QN => n_3945);
   clk_r_REG7726_S8 : DFFS_X1 port map( D => n5332, CK => CLK, SN => RST, Q => 
                           n5331, QN => n_3946);
   clk_r_REG7525_S6 : DFFS_X1 port map( D => n5898, CK => CLK, SN => RST, Q => 
                           n5330, QN => n_3947);
   clk_r_REG7526_S7 : DFFS_X1 port map( D => n5330, CK => CLK, SN => RST, Q => 
                           n5329, QN => n_3948);
   clk_r_REG7527_S8 : DFFS_X1 port map( D => n5329, CK => CLK, SN => RST, Q => 
                           n5328, QN => n_3949);
   clk_r_REG7946_S6 : DFFS_X1 port map( D => n5920, CK => CLK, SN => RST, Q => 
                           n_3950, QN => n5531);
   clk_r_REG7947_S7 : DFFR_X1 port map( D => n5531, CK => CLK, RN => RST, Q => 
                           n_3951, QN => n5326);
   clk_r_REG10023_S4 : DFFR_X1 port map( D => n5530, CK => CLK, RN => RST, Q =>
                           n5325, QN => n_3952);
   clk_r_REG10124_S4 : DFFR_X1 port map( D => n5866, CK => CLK, RN => RST, Q =>
                           n5324, QN => n_3953);
   clk_r_REG10104_S2 : DFFR_X1 port map( D => n4187, CK => CLK, RN => RST, Q =>
                           n5323, QN => n_3954);
   clk_r_REG10019_S1 : DFFS_X1 port map( D => n5513, CK => CLK, SN => RST, Q =>
                           n5322, QN => n_3955);
   clk_r_REG7633_S6 : DFFR_X1 port map( D => n5507, CK => CLK, RN => RST, Q => 
                           n_3956, QN => n5517);
   clk_r_REG7634_S7 : DFFS_X1 port map( D => n5517, CK => CLK, SN => RST, Q => 
                           n_3957, QN => n5320);
   clk_r_REG7514_S8 : DFFS_X1 port map( D => n5527, CK => CLK, SN => RST, Q => 
                           n5319, QN => n_3958);
   clk_r_REG7512_S7 : DFFR_X1 port map( D => n5506, CK => CLK, RN => RST, Q => 
                           n_3959, QN => n5527);
   clk_r_REG7513_S8 : DFFS_X1 port map( D => n5527, CK => CLK, SN => RST, Q => 
                           n_3960, QN => n5317);
   clk_r_REG8035_S7 : DFFR_X1 port map( D => n5508, CK => CLK, RN => RST, Q => 
                           n_3961, QN => n5529);
   clk_r_REG8036_S8 : DFFS_X1 port map( D => n5529, CK => CLK, SN => RST, Q => 
                           n_3962, QN => n5315);
   clk_r_REG8178_S8 : DFFS_X1 port map( D => n5526, CK => CLK, SN => RST, Q => 
                           n5314, QN => n_3963);
   clk_r_REG8176_S7 : DFFR_X1 port map( D => n5922, CK => CLK, RN => RST, Q => 
                           n_3964, QN => n5526);
   clk_r_REG8177_S8 : DFFS_X1 port map( D => n5526, CK => CLK, SN => RST, Q => 
                           n_3965, QN => n5312);
   clk_r_REG8164_S7 : DFFS_X1 port map( D => n5525, CK => CLK, SN => RST, Q => 
                           n5311, QN => n_3966);
   clk_r_REG8162_S6 : DFFR_X1 port map( D => n5924, CK => CLK, RN => RST, Q => 
                           n_3967, QN => n5525);
   clk_r_REG8163_S7 : DFFS_X1 port map( D => n5525, CK => CLK, SN => RST, Q => 
                           n_3968, QN => n5309);
   clk_r_REG8156_S7 : DFFS_X1 port map( D => n5524, CK => CLK, SN => RST, Q => 
                           n5308, QN => n_3969);
   clk_r_REG8154_S6 : DFFR_X1 port map( D => n5926, CK => CLK, RN => RST, Q => 
                           n_3970, QN => n5524);
   clk_r_REG8155_S7 : DFFS_X1 port map( D => n5524, CK => CLK, SN => RST, Q => 
                           n_3971, QN => n5306);
   clk_r_REG8148_S7 : DFFS_X1 port map( D => n5523, CK => CLK, SN => RST, Q => 
                           n5305, QN => n_3972);
   clk_r_REG8146_S6 : DFFR_X1 port map( D => n5928, CK => CLK, RN => RST, Q => 
                           n_3973, QN => n5523);
   clk_r_REG8147_S7 : DFFS_X1 port map( D => n5523, CK => CLK, SN => RST, Q => 
                           n_3974, QN => n5303);
   clk_r_REG8140_S7 : DFFS_X1 port map( D => n5522, CK => CLK, SN => RST, Q => 
                           n5302, QN => n_3975);
   clk_r_REG8138_S6 : DFFR_X1 port map( D => n5930, CK => CLK, RN => RST, Q => 
                           n_3976, QN => n5522);
   clk_r_REG8139_S7 : DFFS_X1 port map( D => n5522, CK => CLK, SN => RST, Q => 
                           n_3977, QN => n5300);
   clk_r_REG8133_S7 : DFFS_X1 port map( D => n5521, CK => CLK, SN => RST, Q => 
                           n5299, QN => n_3978);
   clk_r_REG8131_S6 : DFFR_X1 port map( D => n5932, CK => CLK, RN => RST, Q => 
                           n_3979, QN => n5521);
   clk_r_REG8132_S7 : DFFS_X1 port map( D => n5521, CK => CLK, SN => RST, Q => 
                           n_3980, QN => n5297);
   clk_r_REG8126_S7 : DFFS_X1 port map( D => n5520, CK => CLK, SN => RST, Q => 
                           n5296, QN => n_3981);
   clk_r_REG8124_S6 : DFFR_X1 port map( D => n5934, CK => CLK, RN => RST, Q => 
                           n_3982, QN => n5520);
   clk_r_REG8125_S7 : DFFS_X1 port map( D => n5520, CK => CLK, SN => RST, Q => 
                           n_3983, QN => n5294);
   clk_r_REG8118_S7 : DFFS_X1 port map( D => n5519, CK => CLK, SN => RST, Q => 
                           n5293, QN => n_3984);
   clk_r_REG8116_S6 : DFFR_X1 port map( D => n5936, CK => CLK, RN => RST, Q => 
                           n_3985, QN => n5519);
   clk_r_REG8117_S7 : DFFS_X1 port map( D => n5519, CK => CLK, SN => RST, Q => 
                           n_3986, QN => n5291);
   clk_r_REG8111_S7 : DFFS_X1 port map( D => n5518, CK => CLK, SN => RST, Q => 
                           n5290, QN => n_3987);
   clk_r_REG8109_S6 : DFFR_X1 port map( D => n5938, CK => CLK, RN => RST, Q => 
                           n_3988, QN => n5518);
   clk_r_REG8110_S7 : DFFS_X1 port map( D => n5518, CK => CLK, SN => RST, Q => 
                           n_3989, QN => n5288);
   clk_r_REG9915_S3 : DFFR_X1 port map( D => n5870, CK => CLK, RN => RST, Q => 
                           n_3990, QN => n5528);
   clk_r_REG9916_S4 : DFFS_X1 port map( D => n5528, CK => CLK, SN => RST, Q => 
                           n6220, QN => n5286);
   clk_r_REG10098_S4 : DFFS_X1 port map( D => n5868, CK => CLK, SN => RST, Q =>
                           n5285, QN => n_3991);
   clk_r_REG10257_S6 : DFFS_X1 port map( D => n5874, CK => CLK, SN => RST, Q =>
                           n5284, QN => n_3992);
   clk_r_REG7012_S3 : DFFR_X1 port map( D => n5283, CK => CLK, RN => RST, Q => 
                           n5282, QN => n_3993);
   clk_r_REG9376_S2 : DFF_X1 port map( D => n1671, CK => CLK, Q => n5281, QN =>
                           n_3994);
   clk_r_REG9377_S3 : DFFR_X1 port map( D => n5281, CK => CLK, RN => RST, Q => 
                           n5280, QN => n_3995);
   clk_r_REG9440_S2 : DFF_X1 port map( D => n1669, CK => CLK, Q => n5279, QN =>
                           n_3996);
   clk_r_REG9441_S3 : DFFR_X1 port map( D => n5279, CK => CLK, RN => RST, Q => 
                           n5278, QN => n_3997);
   clk_r_REG9504_S2 : DFF_X1 port map( D => n1667, CK => CLK, Q => n5277, QN =>
                           n_3998);
   clk_r_REG9505_S3 : DFFR_X1 port map( D => n5277, CK => CLK, RN => RST, Q => 
                           n5276, QN => n_3999);
   clk_r_REG9568_S2 : DFF_X1 port map( D => n1665, CK => CLK, Q => n5275, QN =>
                           n_4000);
   clk_r_REG9569_S3 : DFFR_X1 port map( D => n5275, CK => CLK, RN => RST, Q => 
                           n5274, QN => n_4001);
   clk_r_REG9632_S2 : DFF_X1 port map( D => n1663, CK => CLK, Q => n5273, QN =>
                           n_4002);
   clk_r_REG9633_S3 : DFFR_X1 port map( D => n5273, CK => CLK, RN => RST, Q => 
                           n5272, QN => n_4003);
   clk_r_REG9696_S2 : DFF_X1 port map( D => n1661, CK => CLK, Q => n5271, QN =>
                           n_4004);
   clk_r_REG9697_S3 : DFFR_X1 port map( D => n5271, CK => CLK, RN => RST, Q => 
                           n5270, QN => n_4005);
   clk_r_REG7112_S2 : DFF_X1 port map( D => n1659, CK => CLK, Q => n5269, QN =>
                           n_4006);
   clk_r_REG7113_S3 : DFFR_X1 port map( D => n5269, CK => CLK, RN => RST, Q => 
                           n5268, QN => n_4007);
   clk_r_REG7032_S2 : DFF_X1 port map( D => n1657, CK => CLK, Q => n5267, QN =>
                           n_4008);
   clk_r_REG7033_S3 : DFFR_X1 port map( D => n5267, CK => CLK, RN => RST, Q => 
                           n5266, QN => n_4009);
   clk_r_REG9248_S2 : DFF_X1 port map( D => n1655, CK => CLK, Q => n5265, QN =>
                           n_4010);
   clk_r_REG9249_S3 : DFFR_X1 port map( D => n5265, CK => CLK, RN => RST, Q => 
                           n5264, QN => n_4011);
   clk_r_REG7152_S2 : DFF_X1 port map( D => n1653, CK => CLK, Q => n5263, QN =>
                           n_4012);
   clk_r_REG7153_S3 : DFFR_X1 port map( D => n5263, CK => CLK, RN => RST, Q => 
                           n5262, QN => n_4013);
   clk_r_REG9760_S2 : DFF_X1 port map( D => n1651, CK => CLK, Q => n5261, QN =>
                           n_4014);
   clk_r_REG9761_S3 : DFFR_X1 port map( D => n5261, CK => CLK, RN => RST, Q => 
                           n5260, QN => n_4015);
   clk_r_REG8739_S2 : DFF_X1 port map( D => n1649, CK => CLK, Q => n5259, QN =>
                           n_4016);
   clk_r_REG8740_S3 : DFFR_X1 port map( D => n5259, CK => CLK, RN => RST, Q => 
                           n5258, QN => n_4017);
   clk_r_REG8803_S2 : DFF_X1 port map( D => n1647, CK => CLK, Q => n5257, QN =>
                           n_4018);
   clk_r_REG8804_S3 : DFFR_X1 port map( D => n5257, CK => CLK, RN => RST, Q => 
                           n5256, QN => n_4019);
   clk_r_REG8867_S2 : DFF_X1 port map( D => n1645, CK => CLK, Q => n5255, QN =>
                           n_4020);
   clk_r_REG8868_S3 : DFFR_X1 port map( D => n5255, CK => CLK, RN => RST, Q => 
                           n5254, QN => n_4021);
   clk_r_REG8931_S2 : DFF_X1 port map( D => n1643, CK => CLK, Q => n5253, QN =>
                           n_4022);
   clk_r_REG8932_S3 : DFFR_X1 port map( D => n5253, CK => CLK, RN => RST, Q => 
                           n5252, QN => n_4023);
   clk_r_REG8484_S2 : DFF_X1 port map( D => n1641, CK => CLK, Q => n5251, QN =>
                           n_4024);
   clk_r_REG8485_S3 : DFFR_X1 port map( D => n5251, CK => CLK, RN => RST, Q => 
                           n5250, QN => n_4025);
   clk_r_REG7267_S2 : DFF_X1 port map( D => n1639, CK => CLK, Q => n5249, QN =>
                           n_4026);
   clk_r_REG7268_S3 : DFFR_X1 port map( D => n5249, CK => CLK, RN => RST, Q => 
                           n5248, QN => n_4027);
   clk_r_REG8548_S2 : DFF_X1 port map( D => n1637, CK => CLK, Q => n5247, QN =>
                           n_4028);
   clk_r_REG8549_S3 : DFFR_X1 port map( D => n5247, CK => CLK, RN => RST, Q => 
                           n5246, QN => n_4029);
   clk_r_REG8612_S2 : DFF_X1 port map( D => n1635, CK => CLK, Q => n5245, QN =>
                           n_4030);
   clk_r_REG8613_S3 : DFFR_X1 port map( D => n5245, CK => CLK, RN => RST, Q => 
                           n5244, QN => n_4031);
   clk_r_REG9057_S2 : DFF_X1 port map( D => n1633, CK => CLK, Q => n5243, QN =>
                           n_4032);
   clk_r_REG9058_S3 : DFFR_X1 port map( D => n5243, CK => CLK, RN => RST, Q => 
                           n5242, QN => n_4033);
   clk_r_REG9121_S2 : DFF_X1 port map( D => n1631, CK => CLK, Q => n5241, QN =>
                           n_4034);
   clk_r_REG7366_S2 : DFF_X1 port map( D => n1629, CK => CLK, Q => n5240, QN =>
                           n_4035);
   clk_r_REG7406_S2 : DFF_X1 port map( D => n1627, CK => CLK, Q => n5239, QN =>
                           n_4036);
   clk_r_REG7560_S2 : DFF_X1 port map( D => n1625, CK => CLK, Q => n5238, QN =>
                           n_4037);
   clk_r_REG7651_S2 : DFF_X1 port map( D => n1623, CK => CLK, Q => n5237, QN =>
                           n_4038);
   clk_r_REG7954_S2 : DFF_X1 port map( D => n1621, CK => CLK, Q => n5236, QN =>
                           n_4039);
   clk_r_REG7872_S2 : DFF_X1 port map( D => n1619, CK => CLK, Q => n5235, QN =>
                           n_4040);
   clk_r_REG9824_S2 : DFF_X1 port map( D => n1617, CK => CLK, Q => n5234, QN =>
                           n_4041);
   clk_r_REG8204_S2 : DFF_X1 port map( D => n1615, CK => CLK, Q => n5233, QN =>
                           n_4042);
   clk_r_REG8346_S2 : DFF_X1 port map( D => n1614, CK => CLK, Q => n5232, QN =>
                           n_4043);
   clk_r_REG6924_S2 : DFF_X1 port map( D => n1613, CK => CLK, Q => n5231, QN =>
                           n_4044);
   clk_r_REG7006_S2 : DFF_X1 port map( D => n3381, CK => CLK, Q => n5230, QN =>
                           n_4045);
   clk_r_REG7007_S3 : DFFR_X1 port map( D => n5230, CK => CLK, RN => RST, Q => 
                           n5229, QN => n_4046);
   clk_r_REG7008_S4 : DFFR_X1 port map( D => n5229, CK => CLK, RN => RST, Q => 
                           n5228, QN => n_4047);
   clk_r_REG6997_S2 : DFF_X1 port map( D => n3378, CK => CLK, Q => n5227, QN =>
                           n_4048);
   clk_r_REG6998_S3 : DFFR_X1 port map( D => n5227, CK => CLK, RN => RST, Q => 
                           n5226, QN => n_4049);
   clk_r_REG6999_S4 : DFFR_X1 port map( D => n5226, CK => CLK, RN => RST, Q => 
                           n5225, QN => n_4050);
   clk_r_REG6988_S2 : DFF_X1 port map( D => n3375, CK => CLK, Q => n5224, QN =>
                           n_4051);
   clk_r_REG6989_S3 : DFFR_X1 port map( D => n5224, CK => CLK, RN => RST, Q => 
                           n5223, QN => n_4052);
   clk_r_REG6990_S4 : DFFR_X1 port map( D => n5223, CK => CLK, RN => RST, Q => 
                           n5222, QN => n_4053);
   clk_r_REG6981_S2 : DFF_X1 port map( D => n3372, CK => CLK, Q => n5221, QN =>
                           n_4054);
   clk_r_REG6982_S3 : DFFR_X1 port map( D => n5221, CK => CLK, RN => RST, Q => 
                           n5220, QN => n_4055);
   clk_r_REG6983_S4 : DFFR_X1 port map( D => n5220, CK => CLK, RN => RST, Q => 
                           n5219, QN => n_4056);
   clk_r_REG6974_S2 : DFF_X1 port map( D => n3369, CK => CLK, Q => n5218, QN =>
                           n_4057);
   clk_r_REG6975_S3 : DFFR_X1 port map( D => n5218, CK => CLK, RN => RST, Q => 
                           n5217, QN => n_4058);
   clk_r_REG6976_S4 : DFFR_X1 port map( D => n5217, CK => CLK, RN => RST, Q => 
                           n5216, QN => n_4059);
   clk_r_REG6967_S2 : DFF_X1 port map( D => n3366, CK => CLK, Q => n5215, QN =>
                           n_4060);
   clk_r_REG6968_S3 : DFFR_X1 port map( D => n5215, CK => CLK, RN => RST, Q => 
                           n5214, QN => n_4061);
   clk_r_REG6969_S4 : DFFR_X1 port map( D => n5214, CK => CLK, RN => RST, Q => 
                           n5213, QN => n_4062);
   clk_r_REG6959_S2 : DFF_X1 port map( D => n3363, CK => CLK, Q => n5212, QN =>
                           n_4063);
   clk_r_REG6960_S3 : DFFR_X1 port map( D => n5212, CK => CLK, RN => RST, Q => 
                           n5211, QN => n_4064);
   clk_r_REG6961_S4 : DFFR_X1 port map( D => n5211, CK => CLK, RN => RST, Q => 
                           n5210, QN => n_4065);
   clk_r_REG7107_S2 : DFF_X1 port map( D => n3360, CK => CLK, Q => n5209, QN =>
                           n_4066);
   clk_r_REG7108_S3 : DFFR_X1 port map( D => n5209, CK => CLK, RN => RST, Q => 
                           n5208, QN => n_4067);
   clk_r_REG7109_S4 : DFFR_X1 port map( D => n5208, CK => CLK, RN => RST, Q => 
                           n5207, QN => n_4068);
   clk_r_REG7028_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n5206, QN =>
                           n_4069);
   clk_r_REG7029_S2 : DFFR_X1 port map( D => n5206, CK => CLK, RN => RST, Q => 
                           n5205, QN => n_4070);
   clk_r_REG7030_S3 : DFFR_X1 port map( D => n5205, CK => CLK, RN => RST, Q => 
                           n5204, QN => n_4071);
   clk_r_REG7020_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n5203, QN =>
                           n_4072);
   clk_r_REG7021_S2 : DFFR_X1 port map( D => n5203, CK => CLK, RN => RST, Q => 
                           n5202, QN => n_4073);
   clk_r_REG7022_S3 : DFFR_X1 port map( D => n5202, CK => CLK, RN => RST, Q => 
                           n5201, QN => n_4074);
   clk_r_REG7147_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n5200, QN =>
                           n_4075);
   clk_r_REG7148_S2 : DFFR_X1 port map( D => n5200, CK => CLK, RN => RST, Q => 
                           n5199, QN => n_4076);
   clk_r_REG7149_S3 : DFFR_X1 port map( D => n5199, CK => CLK, RN => RST, Q => 
                           n5198, QN => n_4077);
   clk_r_REG6952_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n5197, QN =>
                           n_4078);
   clk_r_REG6953_S2 : DFFR_X1 port map( D => n5197, CK => CLK, RN => RST, Q => 
                           n5196, QN => n_4079);
   clk_r_REG6954_S3 : DFFR_X1 port map( D => n5196, CK => CLK, RN => RST, Q => 
                           n5195, QN => n_4080);
   clk_r_REG7140_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n5194, QN =>
                           n_4081);
   clk_r_REG7141_S2 : DFFR_X1 port map( D => n5194, CK => CLK, RN => RST, Q => 
                           n5193, QN => n_4082);
   clk_r_REG7142_S3 : DFFR_X1 port map( D => n5193, CK => CLK, RN => RST, Q => 
                           n5192, QN => n_4083);
   clk_r_REG7133_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n5191, QN =>
                           n_4084);
   clk_r_REG7134_S2 : DFFR_X1 port map( D => n5191, CK => CLK, RN => RST, Q => 
                           n5190, QN => n_4085);
   clk_r_REG7135_S3 : DFFR_X1 port map( D => n5190, CK => CLK, RN => RST, Q => 
                           n5189, QN => n_4086);
   clk_r_REG7126_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n5188, QN =>
                           n_4087);
   clk_r_REG7127_S2 : DFFR_X1 port map( D => n5188, CK => CLK, RN => RST, Q => 
                           n5187, QN => n_4088);
   clk_r_REG7128_S3 : DFFR_X1 port map( D => n5187, CK => CLK, RN => RST, Q => 
                           n5186, QN => n_4089);
   clk_r_REG7119_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n5185, QN =>
                           n_4090);
   clk_r_REG7120_S2 : DFFR_X1 port map( D => n5185, CK => CLK, RN => RST, Q => 
                           n5184, QN => n_4091);
   clk_r_REG7121_S3 : DFFR_X1 port map( D => n5184, CK => CLK, RN => RST, Q => 
                           n5183, QN => n_4092);
   clk_r_REG7238_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n5182, QN =>
                           n_4093);
   clk_r_REG7239_S2 : DFFR_X1 port map( D => n5182, CK => CLK, RN => RST, Q => 
                           n5181, QN => n_4094);
   clk_r_REG7240_S3 : DFFR_X1 port map( D => n5181, CK => CLK, RN => RST, Q => 
                           n5180, QN => n_4095);
   clk_r_REG7257_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n5179, QN =>
                           n_4096);
   clk_r_REG7258_S2 : DFFR_X1 port map( D => n5179, CK => CLK, RN => RST, Q => 
                           n5178, QN => n_4097);
   clk_r_REG7259_S3 : DFFR_X1 port map( D => n5178, CK => CLK, RN => RST, Q => 
                           n5177, QN => n_4098);
   clk_r_REG7187_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n5176, QN =>
                           n_4099);
   clk_r_REG7188_S2 : DFFR_X1 port map( D => n5176, CK => CLK, RN => RST, Q => 
                           n5175, QN => n_4100);
   clk_r_REG7189_S3 : DFFR_X1 port map( D => n5175, CK => CLK, RN => RST, Q => 
                           n5174, QN => n_4101);
   clk_r_REG7169_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n5173, QN =>
                           n_4102);
   clk_r_REG7170_S2 : DFFR_X1 port map( D => n5173, CK => CLK, RN => RST, Q => 
                           n5172, QN => n_4103);
   clk_r_REG7171_S3 : DFFR_X1 port map( D => n5172, CK => CLK, RN => RST, Q => 
                           n5171, QN => n_4104);
   clk_r_REG7066_S2 : DFF_X1 port map( D => n3321, CK => CLK, Q => n5170, QN =>
                           n_4105);
   clk_r_REG7067_S3 : DFFR_X1 port map( D => n5170, CK => CLK, RN => RST, Q => 
                           n5169, QN => n_4106);
   clk_r_REG7068_S4 : DFFR_X1 port map( D => n5169, CK => CLK, RN => RST, Q => 
                           n5168, QN => n_4107);
   clk_r_REG7047_S2 : DFF_X1 port map( D => n3318, CK => CLK, Q => n5167, QN =>
                           n_4108);
   clk_r_REG7048_S3 : DFFR_X1 port map( D => n5167, CK => CLK, RN => RST, Q => 
                           n5166, QN => n_4109);
   clk_r_REG7049_S4 : DFFR_X1 port map( D => n5166, CK => CLK, RN => RST, Q => 
                           n5165, QN => n_4110);
   clk_r_REG7330_S2 : DFF_X1 port map( D => n3315, CK => CLK, Q => n5164, QN =>
                           n_4111);
   clk_r_REG7331_S3 : DFFR_X1 port map( D => n5164, CK => CLK, RN => RST, Q => 
                           n5163, QN => n_4112);
   clk_r_REG7332_S4 : DFFR_X1 port map( D => n5163, CK => CLK, RN => RST, Q => 
                           n5162, QN => n_4113);
   clk_r_REG7400_S2 : DFF_X1 port map( D => n3312, CK => CLK, Q => n5161, QN =>
                           n_4114);
   clk_r_REG7401_S3 : DFFR_X1 port map( D => n5161, CK => CLK, RN => RST, Q => 
                           n5160, QN => n_4115);
   clk_r_REG7402_S4 : DFFR_X1 port map( D => n5160, CK => CLK, RN => RST, Q => 
                           n5159, QN => n_4116);
   clk_r_REG7549_S2 : DFF_X1 port map( D => n3309, CK => CLK, Q => n5158, QN =>
                           n_4117);
   clk_r_REG7550_S3 : DFFR_X1 port map( D => n5158, CK => CLK, RN => RST, Q => 
                           n5157, QN => n_4118);
   clk_r_REG7551_S4 : DFFR_X1 port map( D => n5157, CK => CLK, RN => RST, Q => 
                           n5156, QN => n_4119);
   clk_r_REG7644_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n5155, QN =>
                           n_4120);
   clk_r_REG7645_S2 : DFFR_X1 port map( D => n5155, CK => CLK, RN => RST, Q => 
                           n5154, QN => n_4121);
   clk_r_REG7646_S3 : DFFR_X1 port map( D => n5154, CK => CLK, RN => RST, Q => 
                           n5153, QN => n_4122);
   clk_r_REG7535_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n5152, QN =>
                           n_4123);
   clk_r_REG7536_S2 : DFFR_X1 port map( D => n5152, CK => CLK, RN => RST, Q => 
                           n5151, QN => n_4124);
   clk_r_REG7537_S3 : DFFR_X1 port map( D => n5151, CK => CLK, RN => RST, Q => 
                           n5150, QN => n_4125);
   clk_r_REG7745_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n5149, QN =>
                           n_4126);
   clk_r_REG7746_S2 : DFFR_X1 port map( D => n5149, CK => CLK, RN => RST, Q => 
                           n5148, QN => n_4127);
   clk_r_REG7747_S3 : DFFR_X1 port map( D => n5148, CK => CLK, RN => RST, Q => 
                           n5147, QN => n_4128);
   clk_r_REG6937_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n5146, QN =>
                           n_4129);
   clk_r_REG6938_S2 : DFFR_X1 port map( D => n5146, CK => CLK, RN => RST, Q => 
                           n5145, QN => n_4130);
   clk_r_REG6939_S3 : DFFR_X1 port map( D => n5145, CK => CLK, RN => RST, Q => 
                           n5144, QN => n_4131);
   clk_r_REG7387_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n5143, QN =>
                           n_4132);
   clk_r_REG7388_S2 : DFFR_X1 port map( D => n5143, CK => CLK, RN => RST, Q => 
                           n5142, QN => n_4133);
   clk_r_REG7389_S3 : DFFR_X1 port map( D => n5142, CK => CLK, RN => RST, Q => 
                           n5141, QN => n_4134);
   clk_r_REG7311_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n5140, QN =>
                           n_4135);
   clk_r_REG7312_S2 : DFFR_X1 port map( D => n5140, CK => CLK, RN => RST, Q => 
                           n5139, QN => n_4136);
   clk_r_REG7313_S3 : DFFR_X1 port map( D => n5139, CK => CLK, RN => RST, Q => 
                           n5138, QN => n_4137);
   clk_r_REG6911_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n5137, QN =>
                           n_4138);
   clk_r_REG6912_S2 : DFFR_X1 port map( D => n5137, CK => CLK, RN => RST, Q => 
                           n5136, QN => n_4139);
   clk_r_REG6913_S3 : DFFR_X1 port map( D => n5136, CK => CLK, RN => RST, Q => 
                           n5135, QN => n_4140);
   clk_r_REG10264_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port, CK 
                           => CLK, RN => RST, Q => n5134, QN => n_4141);
   clk_r_REG10297_S4 : DFFR_X1 port map( D => n3284, CK => CLK, RN => RST, Q =>
                           n_4142, QN => n5539);
   clk_r_REG10298_S4 : DFFR_X1 port map( D => n4417, CK => CLK, RN => RST, Q =>
                           n_4143, QN => n6225);
   clk_r_REG10296_S4 : DFFR_X1 port map( D => n3281, CK => CLK, RN => RST, Q =>
                           n5131, QN => n6224);
   clk_r_REG10259_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port, CK 
                           => CLK, RN => RST, Q => n5130, QN => n_4144);
   clk_r_REG10262_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port, CK 
                           => CLK, RN => RST, Q => n5129, QN => n_4145);
   clk_r_REG10260_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port, CK 
                           => CLK, RN => RST, Q => n5128, QN => n_4146);
   clk_r_REG10109_S2 : DFFS_X1 port map( D => n5885, CK => CLK, SN => RST, Q =>
                           n_4147, QN => n5126);
   clk_r_REG10117_S2 : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => CLK, 
                           RN => RST, Q => n5125, QN => n_4148);
   clk_r_REG10275_S7 : DFFS_X1 port map( D => n5889, CK => CLK, SN => RST, Q =>
                           n5534, QN => n_4149);
   clk_r_REG10121_S2 : DFFS_X1 port map( D => n5881, CK => CLK, SN => RST, Q =>
                           n_4150, QN => n5123);
   clk_r_REG10095_S2 : DFFR_X1 port map( D => n3269, CK => CLK, RN => RST, Q =>
                           n5122, QN => n_4151);
   clk_r_REG8180_S5 : DFFS_X1 port map( D => n4231, CK => CLK, SN => RST, Q => 
                           n5121, QN => n_4152);
   clk_r_REG8172_S7 : DFFR_X1 port map( D => n4230, CK => CLK, RN => RST, Q => 
                           n5120, QN => n_4153);
   clk_r_REG8049_S5 : DFFS_X1 port map( D => n4228, CK => CLK, SN => RST, Q => 
                           n5119, QN => n_4154);
   clk_r_REG10277_S7 : DFFS_X1 port map( D => n474, CK => CLK, SN => RST, Q => 
                           n_4155, QN => n5504);
   clk_r_REG10122_S2 : DFFS_X1 port map( D => n4048, CK => CLK, SN => RST, Q =>
                           n5117, QN => n_4156);
   clk_r_REG10089_S2 : DFFR_X1 port map( D => cu_i_n135, CK => CLK, RN => RST, 
                           Q => n5116, QN => n_4157);
   clk_r_REG10261_S7 : DFFS_X1 port map( D => n477, CK => CLK, SN => RST, Q => 
                           n5115, QN => n_4158);
   clk_r_REG7510_S6 : DFFR_X1 port map( D => n5501, CK => CLK, RN => RST, Q => 
                           n5506, QN => n_4159);
   clk_r_REG7511_S7 : DFFR_X1 port map( D => n5506, CK => CLK, RN => RST, Q => 
                           n_4160, QN => n5113);
   clk_r_REG7631_S5 : DFFR_X1 port map( D => n5502, CK => CLK, RN => RST, Q => 
                           n5507, QN => n_4161);
   clk_r_REG7632_S6 : DFFR_X1 port map( D => n5507, CK => CLK, RN => RST, Q => 
                           n_4162, QN => n5111);
   clk_r_REG8094_S6 : DFFR_X1 port map( D => n5938, CK => CLK, RN => RST, Q => 
                           n_4163, QN => n5110);
   clk_r_REG8088_S6 : DFFR_X1 port map( D => n5936, CK => CLK, RN => RST, Q => 
                           n_4164, QN => n5109);
   clk_r_REG8082_S6 : DFFR_X1 port map( D => n5934, CK => CLK, RN => RST, Q => 
                           n_4165, QN => n5108);
   clk_r_REG8076_S6 : DFFR_X1 port map( D => n5932, CK => CLK, RN => RST, Q => 
                           n_4166, QN => n5107);
   clk_r_REG8069_S6 : DFFR_X1 port map( D => n5930, CK => CLK, RN => RST, Q => 
                           n_4167, QN => n5106);
   clk_r_REG8063_S6 : DFFR_X1 port map( D => n5928, CK => CLK, RN => RST, Q => 
                           n_4168, QN => n5105);
   clk_r_REG8057_S6 : DFFR_X1 port map( D => n5926, CK => CLK, RN => RST, Q => 
                           n_4169, QN => n5104);
   clk_r_REG8050_S6 : DFFR_X1 port map( D => n5924, CK => CLK, RN => RST, Q => 
                           n_4170, QN => n5103);
   clk_r_REG8168_S7 : DFFR_X1 port map( D => n5922, CK => CLK, RN => RST, Q => 
                           n_4171, QN => n5102);
   clk_r_REG8031_S6 : DFFS_X1 port map( D => n4128, CK => CLK, SN => RST, Q => 
                           n_4172, QN => n5508);
   clk_r_REG8032_S7 : DFFR_X1 port map( D => n5508, CK => CLK, RN => RST, Q => 
                           n_4173, QN => n5100);
   clk_r_REG10018_S1 : DFFS_X1 port map( D => n5513, CK => CLK, SN => RST, Q =>
                           n6218, QN => n5099);
   clk_r_REG10085_S4 : DFFS_X1 port map( D => n3261, CK => CLK, SN => RST, Q =>
                           n5098, QN => n_4174);
   clk_r_REG7723_S6 : DFFS_X1 port map( D => n5897, CK => CLK, SN => RST, Q => 
                           n_4175, QN => n5096);
   clk_r_REG9905_S3 : DFFS_X1 port map( D => n3257, CK => CLK, SN => RST, Q => 
                           n5095, QN => n5516);
   clk_r_REG9906_S4 : DFFR_X1 port map( D => n5516, CK => CLK, RN => RST, Q => 
                           n_4176, QN => n5094);
   clk_r_REG10299_S1 : DFFS_X1 port map( D => n3252, CK => CLK, SN => RST, Q =>
                           n5092, QN => n_4177);
   clk_r_REG8044_S5 : DFFS_X1 port map( D => n4341, CK => CLK, SN => RST, Q => 
                           n5091, QN => n_4178);
   clk_r_REG8045_S5 : DFFR_X1 port map( D => n4344, CK => CLK, RN => RST, Q => 
                           n5090, QN => n_4179);
   clk_r_REG10258_S7 : DFFR_X1 port map( D => n3248, CK => CLK, RN => RST, Q =>
                           n5089, QN => n_4180);
   clk_r_REG10283_S7 : DFFS_X1 port map( D => n492, CK => CLK, SN => RST, Q => 
                           n5088, QN => n_4181);
   clk_r_REG10015_S1 : DFFS_X1 port map( D => n5512, CK => CLK, SN => RST, Q =>
                           n_4182, QN => n5087);
   clk_r_REG10017_S2 : DFFR_X1 port map( D => n5087, CK => CLK, RN => RST, Q =>
                           n5086, QN => n_4183);
   clk_r_REG8103_S6 : DFFS_X1 port map( D => n3243, CK => CLK, SN => RST, Q => 
                           n5085, QN => n_4184);
   clk_r_REG6925_S2 : DFF_X1 port map( D => n3242, CK => CLK, Q => n5084, QN =>
                           n_4185);
   clk_r_REG6930_S5 : DFFS_X1 port map( D => n5895, CK => CLK, SN => RST, Q => 
                           n_4186, QN => n5083);
   clk_r_REG10021_S3 : DFFS_X1 port map( D => n3596, CK => CLK, SN => RST, Q =>
                           n_4187, QN => n5530);
   clk_r_REG10266_S7 : DFFS_X1 port map( D => n2299, CK => CLK, SN => RST, Q =>
                           n_4188, QN => n5511);
   clk_r_REG10129_S7 : DFFR_X1 port map( D => n3205, CK => CLK, RN => RST, Q =>
                           n5079, QN => n_4189);
   clk_r_REG10280_S7 : DFFS_X1 port map( D => n5944, CK => CLK, SN => RST, Q =>
                           n_4190, QN => n5078);
   clk_r_REG10282_S7 : DFFR_X1 port map( D => n3236, CK => CLK, RN => RST, Q =>
                           n5077, QN => n_4191);
   clk_r_REG10284_S7 : DFFR_X1 port map( D => n3238, CK => CLK, RN => RST, Q =>
                           n5076, QN => n_4192);
   clk_r_REG10269_S7 : DFFR_X1 port map( D => n3155, CK => CLK, RN => RST, Q =>
                           n5075, QN => n_4193);
   clk_r_REG10088_S2 : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK => CLK, 
                           RN => RST, Q => n5074, QN => n_4194);
   clk_r_REG10125_S4 : DFFS_X1 port map( D => n3235, CK => CLK, SN => RST, Q =>
                           n5073, QN => n_4195);
   clk_r_REG10186_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_16_port,
                           CK => CLK, RN => RST, Q => n5072, QN => n_4196);
   clk_r_REG10285_S7 : DFFR_X1 port map( D => n3227, CK => CLK, RN => RST, Q =>
                           n5071, QN => n_4197);
   clk_r_REG10243_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_20_port,
                           CK => CLK, RN => RST, Q => n5070, QN => n_4198);
   clk_r_REG10246_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_19_port,
                           CK => CLK, RN => RST, Q => n5068, QN => n_4199);
   clk_r_REG10249_S7 : DFFR_X1 port map( D => n3233, CK => CLK, RN => RST, Q =>
                           n5067, QN => n_4200);
   clk_r_REG10250_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_17_port,
                           CK => CLK, RN => RST, Q => n5066, QN => n_4201);
   clk_r_REG10251_S7 : DFFR_X1 port map( D => n3231, CK => CLK, RN => RST, Q =>
                           n5065, QN => n_4202);
   clk_r_REG6929_S5 : DFFS_X1 port map( D => n5921, CK => CLK, SN => RST, Q => 
                           n_4203, QN => IRAM_ADDRESS_2_port);
   clk_r_REG10105_S2 : DFFR_X1 port map( D => n5865, CK => CLK, RN => RST, Q =>
                           n_4204, QN => IRAM_ENABLE);
   clk_r_REG7945_S5 : DFFS_X1 port map( D => n5943, CK => CLK, SN => RST, Q => 
                           n_4205, QN => IRAM_ADDRESS_5_port);
   clk_r_REG7515_S7 : DFFS_X1 port map( D => n5942, CK => CLK, SN => RST, Q => 
                           n_4206, QN => IRAM_ADDRESS_9_port);
   clk_r_REG7629_S4 : DFFS_X1 port map( D => n5941, CK => CLK, SN => RST, Q => 
                           n_4207, QN => IRAM_ADDRESS_7_port);
   clk_r_REG7935_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_4208);
   clk_r_REG7521_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_4209);
   clk_r_REG7721_S5 : DFFR_X1 port map( D => n1453, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_6_port, QN => n_4210);
   clk_r_REG8416_S5 : DFFR_X1 port map( D => n5478, CK => CLK, RN => RST, Q => 
                           n6232, QN => n_4211);
   clk_r_REG8417_S5 : DFFS_X1 port map( D => n5919, CK => CLK, SN => RST, Q => 
                           n_4212, QN => n5055);
   clk_r_REG7524_S6 : DFFS_X1 port map( D => n5898, CK => CLK, SN => RST, Q => 
                           n_4213, QN => n5054);
   clk_r_REG10119_S3 : DFFR_X1 port map( D => n3211, CK => CLK, RN => RST, Q =>
                           n5053, QN => n_4214);
   clk_r_REG10120_S3 : DFFR_X1 port map( D => n3210, CK => CLK, RN => RST, Q =>
                           n5052, QN => n_4215);
   clk_r_REG10099_S3 : DFFR_X1 port map( D => n3209, CK => CLK, RN => RST, Q =>
                           n5051, QN => n_4216);
   clk_r_REG10096_S3 : DFFS_X1 port map( D => n5875, CK => CLK, SN => RST, Q =>
                           n_4217, QN => n5050);
   clk_r_REG10286_S7 : DFFR_X1 port map( D => n3207, CK => CLK, RN => RST, Q =>
                           n5049, QN => n_4218);
   clk_r_REG10288_S7 : DFFR_X1 port map( D => n3206, CK => CLK, RN => RST, Q =>
                           n5048, QN => n_4219);
   clk_r_REG10252_S7 : DFFR_X1 port map( D => n3204, CK => CLK, RN => RST, Q =>
                           n5047, QN => n_4220);
   clk_r_REG10253_S7 : DFFR_X1 port map( D => n3203, CK => CLK, RN => RST, Q =>
                           n5046, QN => n_4221);
   clk_r_REG10291_S7 : DFFR_X1 port map( D => n3202, CK => CLK, RN => RST, Q =>
                           n5045, QN => n_4222);
   clk_r_REG10292_S7 : DFFR_X1 port map( D => n3201, CK => CLK, RN => RST, Q =>
                           n5044, QN => n_4223);
   clk_r_REG10293_S7 : DFFR_X1 port map( D => n3200, CK => CLK, RN => RST, Q =>
                           n5043, QN => n_4224);
   clk_r_REG10294_S7 : DFFR_X1 port map( D => n3199, CK => CLK, RN => RST, Q =>
                           n5042, QN => n_4225);
   clk_r_REG10295_S7 : DFFR_X1 port map( D => n3198, CK => CLK, RN => RST, Q =>
                           n5041, QN => n_4226);
   clk_r_REG10042_S3 : DFFR_X1 port map( D => n3197, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5040, QN => n_4227);
   clk_r_REG10043_S3 : DFFR_X1 port map( D => n3196, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5039, QN => n_4228);
   clk_r_REG10044_S3 : DFFR_X1 port map( D => n3195, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5038, QN => n_4229);
   clk_r_REG10045_S3 : DFFR_X1 port map( D => n3194, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5037, QN => n_4230);
   clk_r_REG10064_S3 : DFFR_X1 port map( D => n3193, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5036, QN => n_4231);
   clk_r_REG10065_S3 : DFFR_X1 port map( D => n3192, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5035, QN => n_4232);
   clk_r_REG10066_S3 : DFFR_X1 port map( D => n3191, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5034, QN => n_4233);
   clk_r_REG10067_S3 : DFFR_X1 port map( D => n3190, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5033, QN => n_4234);
   clk_r_REG10068_S3 : DFFR_X1 port map( D => n3189, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5032, QN => n_4235);
   clk_r_REG10069_S3 : DFFR_X1 port map( D => n3188, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5031, QN => n_4236);
   clk_r_REG10070_S3 : DFFR_X1 port map( D => n3187, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5030, QN => n_4237);
   clk_r_REG10071_S3 : DFFR_X1 port map( D => n3186, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5029, QN => n_4238);
   clk_r_REG10072_S3 : DFFR_X1 port map( D => n3185, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5028, QN => n_4239);
   clk_r_REG10073_S3 : DFFR_X1 port map( D => n3184, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5027, QN => n_4240);
   clk_r_REG10046_S3 : DFFR_X1 port map( D => n3183, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5026, QN => n_4241);
   clk_r_REG10047_S3 : DFFR_X1 port map( D => n3182, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5025, QN => n_4242);
   clk_r_REG10048_S3 : DFFR_X1 port map( D => n3181, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5024, QN => n_4243);
   clk_r_REG10049_S3 : DFFR_X1 port map( D => n3180, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5023, QN => n_4244);
   clk_r_REG10050_S3 : DFFR_X1 port map( D => n3179, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5022, QN => n_4245);
   clk_r_REG10051_S3 : DFFR_X1 port map( D => n3178, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5021, QN => n_4246);
   clk_r_REG10074_S3 : DFFR_X1 port map( D => n3177, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5020, QN => n_4247);
   clk_r_REG10075_S3 : DFFR_X1 port map( D => n3176, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5019, QN => n_4248);
   clk_r_REG10076_S3 : DFFR_X1 port map( D => n3175, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5018, QN => n_4249);
   clk_r_REG10077_S3 : DFFR_X1 port map( D => n3174, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5017, QN => n_4250);
   clk_r_REG10078_S3 : DFFR_X1 port map( D => n3173, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5016, QN => n_4251);
   clk_r_REG10079_S3 : DFFR_X1 port map( D => n3172, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5015, QN => n_4252);
   clk_r_REG10080_S3 : DFFR_X1 port map( D => n3171, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5014, QN => n_4253);
   clk_r_REG10081_S3 : DFFR_X1 port map( D => n3170, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5013, QN => n_4254);
   clk_r_REG10082_S3 : DFFR_X1 port map( D => n3169, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5012, QN => n_4255);
   clk_r_REG10083_S3 : DFFR_X1 port map( D => n3168, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5011, QN => n_4256);
   clk_r_REG10084_S3 : DFFR_X1 port map( D => n3167, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5010, QN => n_4257);
   clk_r_REG10052_S3 : DFFR_X1 port map( D => n3166, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n5009, QN => n_4258);
   clk_r_REG9896_S5 : DFFR_X1 port map( D => n5479, CK => CLK, RN => RST, Q => 
                           n6233, QN => n_4259);
   clk_r_REG9897_S5 : DFFS_X1 port map( D => n5918, CK => CLK, SN => RST, Q => 
                           n_4260, QN => n5007);
   clk_r_REG10100_S4 : DFFR_X1 port map( D => n3160, CK => CLK, RN => RST, Q =>
                           n5006, QN => n_4261);
   clk_r_REG8038_S7 : DFFS_X1 port map( D => n5940, CK => CLK, SN => RST, Q => 
                           n_4262, QN => IRAM_ADDRESS_11_port);
   clk_r_REG8070_S6 : DFFS_X1 port map( D => n5931, CK => CLK, SN => RST, Q => 
                           n_4263, QN => IRAM_ADDRESS_21_port);
   clk_r_REG8064_S6 : DFFS_X1 port map( D => n5929, CK => CLK, SN => RST, Q => 
                           n_4264, QN => IRAM_ADDRESS_19_port);
   clk_r_REG8058_S6 : DFFS_X1 port map( D => n5927, CK => CLK, SN => RST, Q => 
                           n_4265, QN => IRAM_ADDRESS_17_port);
   clk_r_REG8169_S7 : DFFS_X1 port map( D => n5923, CK => CLK, SN => RST, Q => 
                           n_4266, QN => IRAM_ADDRESS_13_port);
   clk_r_REG8051_S6 : DFFS_X1 port map( D => n5925, CK => CLK, SN => RST, Q => 
                           n_4267, QN => IRAM_ADDRESS_15_port);
   clk_r_REG8077_S6 : DFFS_X1 port map( D => n5933, CK => CLK, SN => RST, Q => 
                           n_4268, QN => IRAM_ADDRESS_23_port);
   clk_r_REG8083_S6 : DFFS_X1 port map( D => n5935, CK => CLK, SN => RST, Q => 
                           n_4269, QN => IRAM_ADDRESS_25_port);
   clk_r_REG8089_S6 : DFFS_X1 port map( D => n5937, CK => CLK, SN => RST, Q => 
                           n_4270, QN => IRAM_ADDRESS_27_port);
   clk_r_REG8095_S6 : DFFS_X1 port map( D => n5939, CK => CLK, SN => RST, Q => 
                           n_4271, QN => IRAM_ADDRESS_29_port);
   clk_r_REG10270_S7 : DFFS_X1 port map( D => n5880, CK => CLK, SN => RST, Q =>
                           n6227, QN => n4995);
   clk_r_REG10271_S1 : DFFR_X1 port map( D => n4060, CK => CLK, RN => RST, Q =>
                           n_4272, QN => n5541);
   clk_r_REG10110_S2 : DFFR_X1 port map( D => n5872, CK => CLK, RN => RST, Q =>
                           n_4273, QN => n4993);
   clk_r_REG8179_S5 : DFFS_X1 port map( D => n4155, CK => CLK, SN => RST, Q => 
                           n4992, QN => n_4274);
   clk_r_REG7944_S4 : DFFS_X1 port map( D => n4193, CK => CLK, SN => RST, Q => 
                           n_4275, QN => n6223);
   clk_r_REG10014_S1 : DFFR_X1 port map( D => n4052, CK => CLK, RN => RST, Q =>
                           n4990, QN => n_4276);
   clk_r_REG7367_S3 : DFFS_X1 port map( D => n4268, CK => CLK, SN => RST, Q => 
                           n4989, QN => n_4277);
   clk_r_REG7516_S7 : DFFS_X1 port map( D => n4280, CK => CLK, SN => RST, Q => 
                           n4988, QN => n_4278);
   clk_r_REG7630_S4 : DFFR_X1 port map( D => n3148, CK => CLK, RN => RST, Q => 
                           n4987, QN => n_4279);
   clk_r_REG7936_S5 : DFFR_X1 port map( D => n3147, CK => CLK, RN => RST, Q => 
                           n4986, QN => n_4280);
   clk_r_REG7509_S5 : DFFR_X1 port map( D => n3146, CK => CLK, RN => RST, Q => 
                           n4985, QN => n_4281);
   clk_r_REG8030_S5 : DFFR_X1 port map( D => n3145, CK => CLK, RN => RST, Q => 
                           n4984, QN => n_4282);
   clk_r_REG8167_S6 : DFFR_X1 port map( D => n3144, CK => CLK, RN => RST, Q => 
                           n4983, QN => n_4283);
   clk_r_REG8159_S6 : DFFR_X1 port map( D => n3143, CK => CLK, RN => RST, Q => 
                           n4982, QN => n_4284);
   clk_r_REG8152_S7 : DFFR_X1 port map( D => n3142, CK => CLK, RN => RST, Q => 
                           n4981, QN => n_4285);
   clk_r_REG8144_S7 : DFFR_X1 port map( D => n3141, CK => CLK, RN => RST, Q => 
                           n4980, QN => n_4286);
   clk_r_REG8137_S7 : DFFR_X1 port map( D => n3140, CK => CLK, RN => RST, Q => 
                           n4979, QN => n_4287);
   clk_r_REG8130_S7 : DFFR_X1 port map( D => n3139, CK => CLK, RN => RST, Q => 
                           n4978, QN => n_4288);
   clk_r_REG8122_S7 : DFFR_X1 port map( D => n3138, CK => CLK, RN => RST, Q => 
                           n4977, QN => n_4289);
   clk_r_REG8115_S7 : DFFR_X1 port map( D => n3137, CK => CLK, RN => RST, Q => 
                           n4976, QN => n_4290);
   clk_r_REG8108_S7 : DFFR_X1 port map( D => n3136, CK => CLK, RN => RST, Q => 
                           n4975, QN => n_4291);
   clk_r_REG10106_S2 : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK => CLK, 
                           RN => RST, Q => n4973, QN => n_4292);
   clk_r_REG7522_S5 : DFFS_X1 port map( D => n3133, CK => CLK, SN => RST, Q => 
                           n4972, QN => n_4293);
   clk_r_REG7523_S5 : DFFS_X1 port map( D => n3132, CK => CLK, SN => RST, Q => 
                           n4971, QN => n_4294);
   clk_r_REG7722_S5 : DFFS_X1 port map( D => n3131, CK => CLK, SN => RST, Q => 
                           n4970, QN => n_4295);
   clk_r_REG7505_S5 : DFFS_X1 port map( D => n3130, CK => CLK, SN => RST, Q => 
                           n4969, QN => n_4296);
   clk_r_REG8029_S5 : DFFS_X1 port map( D => n3129, CK => CLK, SN => RST, Q => 
                           n4968, QN => n_4297);
   clk_r_REG8039_S5 : DFFS_X1 port map( D => n3128, CK => CLK, SN => RST, Q => 
                           n4967, QN => n_4298);
   clk_r_REG8040_S6 : DFFS_X1 port map( D => n4967, CK => CLK, SN => RST, Q => 
                           n4966, QN => n_4299);
   clk_r_REG8046_S6 : DFFS_X1 port map( D => n3127, CK => CLK, SN => RST, Q => 
                           n4965, QN => n_4300);
   clk_r_REG8054_S6 : DFFS_X1 port map( D => n3126, CK => CLK, SN => RST, Q => 
                           n4964, QN => n_4301);
   clk_r_REG8149_S6 : DFFS_X1 port map( D => n3125, CK => CLK, SN => RST, Q => 
                           n4963, QN => n_4302);
   clk_r_REG8141_S6 : DFFS_X1 port map( D => n3124, CK => CLK, SN => RST, Q => 
                           n4962, QN => n_4303);
   clk_r_REG8134_S6 : DFFS_X1 port map( D => n3123, CK => CLK, SN => RST, Q => 
                           n4961, QN => n_4304);
   clk_r_REG8127_S6 : DFFS_X1 port map( D => n3122, CK => CLK, SN => RST, Q => 
                           n4960, QN => n_4305);
   clk_r_REG8119_S6 : DFFS_X1 port map( D => n3121, CK => CLK, SN => RST, Q => 
                           n4959, QN => n_4306);
   clk_r_REG8112_S6 : DFFS_X1 port map( D => n3120, CK => CLK, SN => RST, Q => 
                           n4958, QN => n_4307);
   clk_r_REG8105_S6 : DFFS_X1 port map( D => n3119, CK => CLK, SN => RST, Q => 
                           n4957, QN => n_4308);
   clk_r_REG9895_S5 : DFFR_X1 port map( D => n3161, CK => CLK, RN => RST, Q => 
                           n4956, QN => n_4309);
   clk_r_REG9891_S5 : DFFS_X1 port map( D => n5896, CK => CLK, SN => RST, Q => 
                           n_4310, QN => n4955);
   clk_r_REG10267_S7 : DFFS_X1 port map( D => n3239, CK => CLK, SN => RST, Q =>
                           n4954, QN => n_4311);
   clk_r_REG10020_S2 : DFFR_X1 port map( D => n3112, CK => CLK, RN => RST, Q =>
                           n4953, QN => n_4312);
   clk_r_REG10094_S2 : DFFR_X1 port map( D => n302, CK => CLK, RN => RST, Q => 
                           n4952, QN => n_4313);
   clk_r_REG8101_S5 : DFFR_X1 port map( D => n3692, CK => CLK, RN => RST, Q => 
                           n5542, QN => n_4314);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => n5437, ADD_WR(3) => n5436, ADD_WR(2) =>
                           n4953, ADD_WR(1) => n5435, ADD_WR(0) => n5438, 
                           ADD_RD1(4) => n3207, ADD_RD1(3) => n3206, ADD_RD1(2)
                           => n3205, ADD_RD1(1) => n3204, ADD_RD1(0) => n3203, 
                           ADD_RD2(4) => curr_instruction_to_cu_i_20_port, 
                           ADD_RD2(3) => curr_instruction_to_cu_i_19_port, 
                           ADD_RD2(2) => n5876, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n43, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n44, OUT1(31) => n1673, 
                           OUT1(30) => n1671, OUT1(29) => n1669, OUT1(28) => 
                           n1667, OUT1(27) => n1665, OUT1(26) => n1663, 
                           OUT1(25) => n1661, OUT1(24) => n1659, OUT1(23) => 
                           n1657, OUT1(22) => n1655, OUT1(21) => n1653, 
                           OUT1(20) => n1651, OUT1(19) => n1649, OUT1(18) => 
                           n1647, OUT1(17) => n1645, OUT1(16) => n1643, 
                           OUT1(15) => n1641, OUT1(14) => n1639, OUT1(13) => 
                           n1637, OUT1(12) => n1635, OUT1(11) => n1633, 
                           OUT1(10) => n1631, OUT1(9) => n1629, OUT1(8) => 
                           n1627, OUT1(7) => n1625, OUT1(6) => n1623, OUT1(5) 
                           => n1621, OUT1(4) => n1619, OUT1(3) => n1617, 
                           OUT1(2) => n1615, OUT1(1) => n1614, OUT1(0) => n1613
                           , OUT2(31) => n3381, OUT2(30) => n3378, OUT2(29) => 
                           n3375, OUT2(28) => n3372, OUT2(27) => n3369, 
                           OUT2(26) => n3366, OUT2(25) => n3363, OUT2(24) => 
                           n3360, OUT2(23) => n3357, OUT2(22) => n3354, 
                           OUT2(21) => n3351, OUT2(20) => n3348, OUT2(19) => 
                           n3345, OUT2(18) => n3342, OUT2(17) => n3339, 
                           OUT2(16) => n3336, OUT2(15) => n3333, OUT2(14) => 
                           n3330, OUT2(13) => n3327, OUT2(12) => n3324, 
                           OUT2(11) => n3321, OUT2(10) => n3318, OUT2(9) => 
                           n3315, OUT2(8) => n3312, OUT2(7) => n3309, OUT2(6) 
                           => n3306, OUT2(5) => n3303, OUT2(4) => n3300, 
                           OUT2(3) => n3297, OUT2(2) => n3294, OUT2(1) => n3291
                           , OUT2(0) => n3288, RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_4315, mul_exeception => 
                           n_4316, FUNC(0) => n5860, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_4317, 
                           OUTALU(31) => datapath_i_alu_output_val_i_31_port, 
                           OUTALU(30) => datapath_i_alu_output_val_i_30_port, 
                           OUTALU(29) => datapath_i_alu_output_val_i_29_port, 
                           OUTALU(28) => datapath_i_alu_output_val_i_28_port, 
                           OUTALU(27) => datapath_i_alu_output_val_i_27_port, 
                           OUTALU(26) => datapath_i_alu_output_val_i_26_port, 
                           OUTALU(25) => datapath_i_alu_output_val_i_25_port, 
                           OUTALU(24) => datapath_i_alu_output_val_i_24_port, 
                           OUTALU(23) => datapath_i_alu_output_val_i_23_port, 
                           OUTALU(22) => datapath_i_alu_output_val_i_22_port, 
                           OUTALU(21) => datapath_i_alu_output_val_i_21_port, 
                           OUTALU(20) => datapath_i_alu_output_val_i_20_port, 
                           OUTALU(19) => datapath_i_alu_output_val_i_19_port, 
                           OUTALU(18) => datapath_i_alu_output_val_i_18_port, 
                           OUTALU(17) => datapath_i_alu_output_val_i_17_port, 
                           OUTALU(16) => datapath_i_alu_output_val_i_16_port, 
                           OUTALU(15) => datapath_i_alu_output_val_i_15_port, 
                           OUTALU(14) => datapath_i_alu_output_val_i_14_port, 
                           OUTALU(13) => datapath_i_alu_output_val_i_13_port, 
                           OUTALU(12) => datapath_i_alu_output_val_i_12_port, 
                           OUTALU(11) => datapath_i_alu_output_val_i_11_port, 
                           OUTALU(10) => datapath_i_alu_output_val_i_10_port, 
                           OUTALU(9) => datapath_i_alu_output_val_i_9_port, 
                           OUTALU(8) => datapath_i_alu_output_val_i_8_port, 
                           OUTALU(7) => datapath_i_alu_output_val_i_7_port, 
                           OUTALU(6) => datapath_i_alu_output_val_i_6_port, 
                           OUTALU(5) => datapath_i_alu_output_val_i_5_port, 
                           OUTALU(4) => datapath_i_alu_output_val_i_4_port, 
                           OUTALU(3) => datapath_i_alu_output_val_i_3_port, 
                           OUTALU(2) => datapath_i_alu_output_val_i_2_port, 
                           OUTALU(1) => datapath_i_alu_output_val_i_1_port, 
                           OUTALU(0) => datapath_i_alu_output_val_i_0_port, 
                           rst_BAR => RST);
   U2333 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_31_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(31), ZN => n5683
                           );
   U2335 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_30_port, A2 => 
                           n5715, B1 => n6231, B2 => DRAM_DATA(30), ZN => n5684
                           );
   U2337 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_29_port, A2 => 
                           n6230, B1 => n6231, B2 => DRAM_DATA(29), ZN => n5685
                           );
   U2339 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_28_port, A2 => 
                           n6230, B1 => n6231, B2 => DRAM_DATA(28), ZN => n5686
                           );
   U2341 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_27_port, A2 => 
                           n6230, B1 => n6231, B2 => DRAM_DATA(27), ZN => n5687
                           );
   U2343 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_26_port, A2 => 
                           n6230, B1 => n6231, B2 => DRAM_DATA(26), ZN => n5688
                           );
   U2345 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_25_port, A2 => 
                           n5715, B1 => n6231, B2 => DRAM_DATA(25), ZN => n5689
                           );
   U2347 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_24_port, A2 => 
                           n6230, B1 => n6231, B2 => DRAM_DATA(24), ZN => n5690
                           );
   U2349 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_23_port, A2 => 
                           n6230, B1 => n6231, B2 => DRAM_DATA(23), ZN => n5691
                           );
   U2351 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(22), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_22_port, ZN => n5692)
                           ;
   U2353 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(21), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_21_port, ZN => n5693)
                           ;
   U2355 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(20), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_20_port, ZN => n5694)
                           ;
   U2357 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(19), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_19_port, ZN => n5695)
                           ;
   U2359 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(18), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_18_port, ZN => n5696)
                           ;
   U2361 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(17), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_17_port, ZN => n5697)
                           ;
   U2363 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(16), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_16_port, ZN => n5698)
                           ;
   U2365 : AOI22_X1 port map( A1 => n5714, A2 => DRAM_DATA(15), B1 => n6230, B2
                           => datapath_i_alu_output_val_i_15_port, ZN => n5699)
                           ;
   U2367 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_14_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(14), ZN => n5700
                           );
   U2369 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_13_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(13), ZN => n5701
                           );
   U2371 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_12_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(12), ZN => n5702
                           );
   U2373 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_11_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(11), ZN => n5703
                           );
   U2375 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_10_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(10), ZN => n5704
                           );
   U2377 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_9_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(9), ZN => n5705)
                           ;
   U2379 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_8_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(8), ZN => n5706)
                           ;
   U2381 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_7_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(7), ZN => n5707)
                           ;
   U2383 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_6_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(6), ZN => n5708)
                           ;
   U2385 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_5_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(5), ZN => n5709)
                           ;
   U2387 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_4_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(4), ZN => n5710)
                           ;
   U2389 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_3_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(3), ZN => n5711)
                           ;
   U2391 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_2_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(2), ZN => n5712)
                           ;
   U2393 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_1_port, A2 => 
                           n5715, B1 => n5714, B2 => DRAM_DATA(1), ZN => n5713)
                           ;
   U2395 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_0_port, A2 => 
                           n6230, B1 => n5714, B2 => DRAM_DATA(0), ZN => n5716)
                           ;
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   clk_r_REG8102_S5 : DFFR_X1 port map( D => n3692, CK => CLK, RN => RST, Q => 
                           n5465, QN => n_4318);
   clk_r_REG10103_S1 : DFFS_X1 port map( D => n3135, CK => CLK, SN => RST, Q =>
                           n5463, QN => n_4319);
   clk_r_REG7011_S2 : DFF_X1 port map( D => n1673, CK => CLK, Q => n5283, QN =>
                           n_4320);
   clk_r_REG9912_S4 : DFFS_X1 port map( D => n5947, CK => CLK, SN => RST, Q => 
                           n5385, QN => n6219);
   clk_r_REG10112_S2 : DFFR_X1 port map( D => n5871, CK => CLK, RN => RST, Q =>
                           n_4321, QN => n5093);
   clk_r_REG10022_S4 : DFFR_X1 port map( D => n5530, CK => CLK, RN => RST, Q =>
                           n_4322, QN => n5081);
   clk_r_REG10126_S6 : DFFS_X1 port map( D => n5874, CK => CLK, SN => RST, Q =>
                           n6214, QN => n5127);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => n5073, Q => 
                           n3555);
   clk_r_REG10245_S7 : DFFR_X1 port map( D => n3229, CK => CLK, RN => RST, Q =>
                           n5069, QN => n_4323);
   clk_r_REG9911_S4 : DFFS_X1 port map( D => n5947, CK => CLK, SN => RST, Q => 
                           n_4324, QN => n5408);
   clk_r_REG6928_S4 : DFFS_X1 port map( D => n5514, CK => CLK, SN => RST, Q => 
                           n5386, QN => n_4325);
   clk_r_REG10090_S2 : DFFS_X1 port map( D => n5869, CK => CLK, SN => RST, Q =>
                           n5409, QN => n_4326);
   clk_r_REG10091_S2 : DFFS_X1 port map( D => n5869, CK => CLK, SN => RST, Q =>
                           n5387, QN => n_4327);
   clk_r_REG10086_S4 : DFFR_X1 port map( D => n3241, CK => CLK, RN => RST, Q =>
                           n5097, QN => n_4328);
   clk_r_REG10128_S6 : DFFR_X1 port map( D => n3555, CK => CLK, RN => RST, Q =>
                           n5388, QN => n_4329);
   clk_r_REG10102_S1 : DFFS_X1 port map( D => n3135, CK => CLK, SN => RST, Q =>
                           n4974, QN => n_4330);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X2 port map( A => 
                           n5192, EN => n6228, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X2 port map( A => 
                           n5189, EN => n5093, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X2 port map( A => 
                           n5186, EN => n5405, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X2 port map( A => 
                           n5201, EN => n6228, Z => DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X2 port map( A => 
                           n5195, EN => n6228, Z => DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X2 port map( A => 
                           n5183, EN => n6228, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X2 port map( A => 
                           n5180, EN => n6228, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X2 port map( A => 
                           n5198, EN => n5093, Z => DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X2 port map( A => 
                           n5225, EN => n6228, Z => DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X2 port map( A => 
                           n5222, EN => n6228, Z => DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X2 port map( A => 
                           n5219, EN => n6228, Z => DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X2 port map( A => 
                           n5216, EN => n6228, Z => DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X2 port map( A => 
                           n5174, EN => n6228, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X2 port map( A => 
                           n5159, EN => n6228, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X2 port map( A => 
                           n5150, EN => n6228, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X2 port map( A => 
                           n5147, EN => n6228, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X2 port map( A => 
                           n5228, EN => n5093, Z => DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X2 port map( A => 
                           n5213, EN => n5093, Z => DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X2 port map( A => 
                           n5207, EN => n5093, Z => DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X2 port map( A => 
                           n5204, EN => n5093, Z => DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X2 port map( A => 
                           n5168, EN => n5093, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X2 port map( A => 
                           n5162, EN => n5093, Z => DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X2 port map( A => 
                           n5156, EN => n5093, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X2 port map( A => 
                           n5135, EN => n5093, Z => DRAM_DATA(0));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X2 port map( A => 
                           n5210, EN => n5405, Z => DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X2 port map( A => 
                           n5177, EN => n5405, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X2 port map( A => 
                           n5171, EN => n5405, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X2 port map( A => 
                           n5165, EN => n5405, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X2 port map( A => 
                           n5153, EN => n5405, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X2 port map( A => 
                           n5144, EN => n5405, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X2 port map( A => 
                           n5141, EN => n5405, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X2 port map( A => 
                           n5138, EN => n5405, Z => DRAM_DATA(1));
   U2622 : OAI21_X2 port map( B1 => n5420, B2 => n5098, A => n4988, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U2623 : INV_X1 port map( A => n4337, ZN => n5946);
   U2624 : INV_X1 port map( A => n5946, ZN => n5947);
   U2625 : OAI21_X2 port map( B1 => n5098, B2 => n5390, A => n6065, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U2626 : AOI22_X2 port map( A1 => n3555, A2 => cu_i_n135, B1 => n5116, B2 => 
                           n5874, ZN => n5869);
   U2627 : CLKBUF_X1 port map( A => n6232, Z => IRAM_ADDRESS_1_port);
   U2628 : CLKBUF_X1 port map( A => n6233, Z => IRAM_ADDRESS_0_port);
   U2629 : CLKBUF_X1 port map( A => n5542, Z => IRAM_ADDRESS_31_port);
   U2630 : AOI22_X1 port map( A1 => n5388, A2 => cu_i_cmd_alu_op_type_3_port, 
                           B1 => n5461, B2 => n5134, ZN => n6017);
   U2631 : AOI22_X1 port map( A1 => n5388, A2 => cu_i_cmd_alu_op_type_2_port, 
                           B1 => n5461, B2 => n5128, ZN => n6019);
   U2632 : AOI22_X1 port map( A1 => n5388, A2 => cu_i_cmd_alu_op_type_0_port, 
                           B1 => n5461, B2 => n5130, ZN => n6021);
   U2633 : NOR2_X1 port map( A1 => n6019, A2 => n6015, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U2634 : NOR2_X1 port map( A1 => n6021, A2 => n6020, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U2635 : NOR2_X1 port map( A1 => n6018, A2 => n6014, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U2636 : CLKBUF_X1 port map( A => n5081, Z => n6183);
   U2637 : MUX2_X1 port map( A => IRAM_DATA(22), B => n5047, S => n5388, Z => 
                           n3204);
   U2638 : INV_X1 port map( A => n3555, ZN => n5874);
   U2639 : AOI22_X1 port map( A1 => n5388, A2 => n5459, B1 => n5461, B2 => 
                           IRAM_DATA(13), ZN => n6179);
   U2640 : INV_X1 port map( A => n6179, ZN => n5877);
   U2641 : AOI22_X1 port map( A1 => n5127, A2 => n5455, B1 => n5284, B2 => 
                           IRAM_DATA(30), ZN => n5973);
   U2642 : INV_X1 port map( A => n5973, ZN => n5886);
   U2643 : AOI22_X1 port map( A1 => n5127, A2 => n5456, B1 => n5284, B2 => 
                           IRAM_DATA(29), ZN => n6177);
   U2644 : INV_X1 port map( A => n6177, ZN => n5884);
   U2645 : AOI22_X1 port map( A1 => n5127, A2 => n5450, B1 => n5284, B2 => 
                           IRAM_DATA(31), ZN => n5959);
   U2646 : NAND3_X1 port map( A1 => n5886, A2 => n5884, A3 => n5959, ZN => 
                           n5960);
   U2647 : INV_X1 port map( A => n5960, ZN => n5883);
   U2648 : NAND2_X1 port map( A1 => n5284, A2 => IRAM_DATA(26), ZN => n5951);
   U2649 : OAI21_X1 port map( B1 => n6214, B2 => n5538, A => n5951, ZN => n5888
                           );
   U2650 : NAND2_X1 port map( A1 => n5284, A2 => IRAM_DATA(28), ZN => n5952);
   U2651 : OAI21_X1 port map( B1 => n6214, B2 => n5537, A => n5952, ZN => n5887
                           );
   U2652 : AOI22_X1 port map( A1 => n5127, A2 => n5448, B1 => n5284, B2 => 
                           IRAM_DATA(27), ZN => n6148);
   U2653 : INV_X1 port map( A => n6148, ZN => n5892);
   U2654 : INV_X1 port map( A => n5888, ZN => n6212);
   U2655 : INV_X1 port map( A => n5887, ZN => n6144);
   U2656 : NAND3_X1 port map( A1 => n6144, A2 => n5973, A3 => n5892, ZN => 
                           n5953);
   U2657 : NOR3_X1 port map( A1 => n6212, A2 => n5959, A3 => n5953, ZN => n5975
                           );
   U2658 : NAND2_X1 port map( A1 => n5975, A2 => n6218, ZN => n5885);
   U2659 : NOR2_X1 port map( A1 => n5884, A2 => n5885, ZN => 
                           cu_i_cmd_word_3_port);
   U2660 : OAI22_X1 port map( A1 => n5874, A2 => cu_i_cmd_word_3_port, B1 => 
                           n5053, B2 => n3555, ZN => n5954);
   U2661 : INV_X1 port map( A => n5954, ZN => n5873);
   U2662 : INV_X1 port map( A => n5885, ZN => n6029);
   U2663 : OAI22_X1 port map( A1 => n5874, A2 => n6029, B1 => n5052, B2 => 
                           n3555, ZN => n3543);
   U2664 : INV_X1 port map( A => n3543, ZN => n5872);
   U2665 : NAND2_X1 port map( A1 => n5872, A2 => n5954, ZN => n3254);
   U2666 : INV_X1 port map( A => n3254, ZN => n5871);
   U2667 : NOR2_X1 port map( A1 => n5119, A2 => n5372, ZN => n6058);
   U2668 : NAND2_X1 port map( A1 => n6058, A2 => n5342, ZN => n6050);
   U2669 : OAI211_X1 port map( C1 => n6058, C2 => n5342, A => n5407, B => n6050
                           , ZN => n5955);
   U2670 : NAND2_X1 port map( A1 => n4964, A2 => n5955, ZN => n6099);
   U2671 : INV_X1 port map( A => n6099, ZN => n5908);
   U2672 : NOR2_X1 port map( A1 => n5368, A2 => n6050, ZN => n6049);
   U2673 : NAND2_X1 port map( A1 => n6049, A2 => n5343, ZN => n6056);
   U2674 : OAI211_X1 port map( C1 => n6049, C2 => n5343, A => n5407, B => n6056
                           , ZN => n5956);
   U2675 : NAND2_X1 port map( A1 => n4963, A2 => n5956, ZN => n6094);
   U2676 : INV_X1 port map( A => n6094, ZN => n5907);
   U2677 : NOR2_X1 port map( A1 => n5892, A2 => n5888, ZN => n5889);
   U2678 : INV_X1 port map( A => n5889, ZN => n6013);
   U2679 : NAND2_X1 port map( A1 => n6177, A2 => n5959, ZN => n5961);
   U2680 : NOR4_X1 port map( A1 => n6013, A2 => n5887, A3 => n5886, A4 => n5961
                           , ZN => n5880);
   U2681 : NAND2_X1 port map( A1 => n5880, A2 => n6218, ZN => n5881);
   U2682 : AOI22_X1 port map( A1 => n5127, A2 => n6222, B1 => IRAM_DATA(0), B2 
                           => n6214, ZN => n5944);
   U2683 : MUX2_X1 port map( A => IRAM_DATA(4), B => n5076, S => n5127, Z => 
                           n3238);
   U2684 : NAND2_X1 port map( A1 => n5284, A2 => IRAM_DATA(2), ZN => n5957);
   U2685 : OAI21_X1 port map( B1 => n6214, B2 => n5509, A => n5957, ZN => n5879
                           );
   U2686 : MUX2_X1 port map( A => IRAM_DATA(3), B => n5077, S => n5127, Z => 
                           n3236);
   U2687 : NAND2_X1 port map( A1 => n5284, A2 => IRAM_DATA(1), ZN => n5958);
   U2688 : OAI21_X1 port map( B1 => n6214, B2 => n5532, A => n5958, ZN => n5878
                           );
   U2689 : INV_X1 port map( A => n5959, ZN => n5890);
   U2690 : AOI211_X1 port map( C1 => n6144, C2 => n6212, A => n5892, B => n5960
                           , ZN => n4060);
   U2691 : NOR2_X1 port map( A1 => n5890, A2 => n6144, ZN => n5976);
   U2692 : AND2_X1 port map( A1 => n6177, A2 => n5976, ZN => n5972);
   U2693 : AND3_X1 port map( A1 => n6212, A2 => n5972, A3 => n5886, ZN => n3155
                           );
   U2694 : NOR4_X1 port map( A1 => n6148, A2 => n5887, A3 => n5886, A4 => n5961
                           , ZN => n5977);
   U2695 : NAND2_X1 port map( A1 => n5322, A2 => n5977, ZN => n6178);
   U2696 : AOI22_X1 port map( A1 => n5127, A2 => n5449, B1 => n5284, B2 => 
                           IRAM_DATA(5), ZN => n5964);
   U2697 : NAND4_X1 port map( A1 => n3238, A2 => n5879, A3 => n3236, A4 => 
                           n5878, ZN => n5962);
   U2698 : NOR3_X1 port map( A1 => n5964, A2 => n5944, A3 => n5962, ZN => n5992
                           );
   U2699 : NOR3_X1 port map( A1 => n6177, A2 => n5886, A3 => n5890, ZN => n6213
                           );
   U2700 : OAI21_X1 port map( B1 => n6144, B2 => n5892, A => n5888, ZN => n5963
                           );
   U2701 : AOI211_X1 port map( C1 => n6213, C2 => n5963, A => n4060, B => n3155
                           , ZN => n6028);
   U2702 : OAI222_X1 port map( A1 => n6178, A2 => n6212, B1 => n5881, B2 => 
                           n5992, C1 => n6028, C2 => n5099, ZN => n302);
   U2703 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n302, ZN => n3269
                           );
   U2704 : INV_X1 port map( A => n5964, ZN => n5891);
   U2705 : AND2_X1 port map( A1 => n5944, A2 => n5878, ZN => n3248);
   U2706 : NOR2_X1 port map( A1 => n5366, A2 => n6056, ZN => n6055);
   U2707 : NAND2_X1 port map( A1 => n6055, A2 => n5344, ZN => n6053);
   U2708 : OAI211_X1 port map( C1 => n6055, C2 => n5344, A => n5407, B => n6053
                           , ZN => n5965);
   U2709 : NAND2_X1 port map( A1 => n4962, A2 => n5965, ZN => n6111);
   U2710 : INV_X1 port map( A => n6111, ZN => n5905);
   U2711 : MUX2_X1 port map( A => IRAM_DATA(16), B => n5072, S => n5388, Z => 
                           curr_instruction_to_cu_i_16_port);
   U2712 : AOI22_X1 port map( A1 => n5388, A2 => n5453, B1 => n5461, B2 => 
                           IRAM_DATA(18), ZN => n6181);
   U2713 : INV_X1 port map( A => n6181, ZN => n5876);
   U2714 : NOR2_X1 port map( A1 => n5364, A2 => n6053, ZN => n6052);
   U2715 : NAND2_X1 port map( A1 => n6052, A2 => n5345, ZN => n6047);
   U2716 : OAI211_X1 port map( C1 => n6052, C2 => n5345, A => n5407, B => n6047
                           , ZN => n5966);
   U2717 : NAND2_X1 port map( A1 => n4961, A2 => n5966, ZN => n6197);
   U2718 : INV_X1 port map( A => n6197, ZN => n5904);
   U2719 : INV_X1 port map( A => cu_i_n151, ZN => n5867);
   U2720 : NOR2_X1 port map( A1 => n4417, A2 => n3284, ZN => n5967);
   U2721 : NOR2_X1 port map( A1 => n5967, A2 => n5867, ZN => n5866);
   U2722 : NAND3_X1 port map( A1 => cu_i_n151, A2 => n5967, A3 => n3281, ZN => 
                           n3235);
   U2723 : MUX2_X1 port map( A => IRAM_DATA(17), B => n5066, S => n5388, Z => 
                           curr_instruction_to_cu_i_17_port);
   U2724 : MUX2_X1 port map( A => IRAM_DATA(12), B => n5065, S => n5388, Z => 
                           n3231);
   U2725 : INV_X1 port map( A => n6178, ZN => n5882);
   U2726 : CLKBUF_X1 port map( A => n5882, Z => n6229);
   U2727 : INV_X1 port map( A => n5866, ZN => n5986);
   U2728 : NAND2_X1 port map( A1 => n5986, A2 => n3235, ZN => n5993);
   U2729 : AOI21_X1 port map( B1 => n5993, B2 => n5992, A => n5881, ZN => n6182
                           );
   U2730 : INV_X1 port map( A => n6182, ZN => n6180);
   U2731 : AOI221_X1 port map( B1 => n6180, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n6182, C2 =>
                           n3231, A => n6229, ZN => n5968);
   U2732 : INV_X1 port map( A => n5968, ZN => n5861);
   U2733 : MUX2_X1 port map( A => IRAM_DATA(19), B => n5068, S => n5388, Z => 
                           curr_instruction_to_cu_i_19_port);
   U2734 : MUX2_X1 port map( A => IRAM_DATA(14), B => n5067, S => n5388, Z => 
                           n3233);
   U2735 : AOI221_X1 port map( B1 => n6180, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n6182, C2 =>
                           n3233, A => n6229, ZN => n5969);
   U2736 : INV_X1 port map( A => n5969, ZN => n5862);
   U2737 : MUX2_X1 port map( A => IRAM_DATA(11), B => n5071, S => n5127, Z => 
                           n3227);
   U2738 : AOI221_X1 port map( B1 => n6180, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n6182, C2 =>
                           n3227, A => n6229, ZN => n5970);
   U2739 : INV_X1 port map( A => n5970, ZN => n5864);
   U2740 : MUX2_X1 port map( A => IRAM_DATA(20), B => n5070, S => n5388, Z => 
                           curr_instruction_to_cu_i_20_port);
   U2741 : MUX2_X1 port map( A => IRAM_DATA(15), B => n5069, S => n5388, Z => 
                           n3229);
   U2742 : AOI221_X1 port map( B1 => n6180, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n6182, C2 =>
                           n3229, A => n6229, ZN => n5971);
   U2743 : INV_X1 port map( A => n5971, ZN => n5863);
   U2744 : NAND2_X1 port map( A1 => n6148, A2 => n5888, ZN => n474);
   U2745 : NAND3_X1 port map( A1 => n5973, A2 => n5322, A3 => n5972, ZN => 
                           n6012);
   U2746 : NOR2_X1 port map( A1 => n6012, A2 => n474, ZN => n4187);
   U2747 : INV_X1 port map( A => n6028, ZN => n5974);
   U2748 : AOI211_X1 port map( C1 => n5976, C2 => n5889, A => n5975, B => n5974
                           , ZN => n5985);
   U2749 : INV_X1 port map( A => n5977, ZN => n5978);
   U2750 : NAND2_X1 port map( A1 => n5985, A2 => n5978, ZN => n6026);
   U2751 : AOI21_X1 port map( B1 => n6218, B2 => n6026, A => n4187, ZN => n5979
                           );
   U2752 : INV_X1 port map( A => n5979, ZN => n301);
   U2753 : NOR2_X1 port map( A1 => n5374, A2 => n6047, ZN => n6046);
   U2754 : NAND2_X1 port map( A1 => n6046, A2 => n5346, ZN => n6044);
   U2755 : OAI211_X1 port map( C1 => n6046, C2 => n5346, A => n5407, B => n6044
                           , ZN => n5980);
   U2756 : NAND2_X1 port map( A1 => n4960, A2 => n5980, ZN => n6092);
   U2757 : INV_X1 port map( A => n6092, ZN => n5903);
   U2758 : NOR2_X1 port map( A1 => n5376, A2 => n6044, ZN => n6043);
   U2759 : NAND2_X1 port map( A1 => n6043, A2 => n5347, ZN => n6038);
   U2760 : OAI211_X1 port map( C1 => n6043, C2 => n5347, A => n5407, B => n6038
                           , ZN => n5981);
   U2761 : NAND2_X1 port map( A1 => n4959, A2 => n5981, ZN => n6089);
   U2762 : INV_X1 port map( A => n6089, ZN => n5902);
   U2763 : INV_X1 port map( A => n5881, ZN => n5982);
   U2764 : NAND2_X1 port map( A1 => n5982, A2 => n5992, ZN => n4048);
   U2765 : NOR2_X1 port map( A1 => n5986, A2 => n4048, ZN => n5983);
   U2766 : NOR2_X1 port map( A1 => n5983, A2 => n5006, ZN => n5987);
   U2767 : AND3_X1 port map( A1 => n5987, A2 => n6183, A3 => DRAM_READY, ZN => 
                           n5714);
   U2768 : CLKBUF_X1 port map( A => n5714, Z => n6231);
   U2769 : INV_X1 port map( A => n4187, ZN => n5984);
   U2770 : OAI211_X1 port map( C1 => n5099, C2 => n5985, A => n6180, B => n5984
                           , ZN => enable_rf_i);
   U2771 : OAI21_X1 port map( B1 => n5986, B2 => n4048, A => n5285, ZN => 
                           write_rf_i);
   U2772 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U2773 : NOR2_X1 port map( A1 => n5987, A2 => n5325, ZN => n5715);
   U2774 : CLKBUF_X1 port map( A => n5715, Z => n6230);
   U2775 : NOR2_X1 port map( A1 => n5378, A2 => n6038, ZN => n6037);
   U2776 : NAND2_X1 port map( A1 => n6037, A2 => n5348, ZN => n6041);
   U2777 : OAI211_X1 port map( C1 => n6037, C2 => n5348, A => n5407, B => n6041
                           , ZN => n5988);
   U2778 : NAND2_X1 port map( A1 => n4958, A2 => n5988, ZN => n6087);
   U2779 : INV_X1 port map( A => n6087, ZN => n5901);
   U2780 : NOR2_X1 port map( A1 => n5380, A2 => n6041, ZN => n6040);
   U2781 : NAND2_X1 port map( A1 => n6040, A2 => n5349, ZN => n5990);
   U2782 : XOR2_X1 port map( A => n5542, B => n5990, Z => n5989);
   U2783 : AOI22_X1 port map( A1 => n5407, A2 => n5989, B1 => n5384, B2 => 
                           n5085, ZN => n6203);
   U2784 : INV_X1 port map( A => n6203, ZN => n5899);
   U2785 : OAI211_X1 port map( C1 => n6040, C2 => n5349, A => n5407, B => n5990
                           , ZN => n5991);
   U2786 : NAND2_X1 port map( A1 => n4957, A2 => n5991, ZN => n6085);
   U2787 : INV_X1 port map( A => n6085, ZN => n5900);
   U2788 : NAND2_X1 port map( A1 => n5880, A2 => n5992, ZN => n477);
   U2789 : INV_X1 port map( A => n5993, ZN => n5994);
   U2790 : OAI21_X1 port map( B1 => n5994, B2 => n5881, A => n5092, ZN => n5995
                           );
   U2791 : OAI221_X1 port map( B1 => n5995, B2 => n5322, C1 => n5995, C2 => 
                           n477, A => n5874, ZN => n5865);
   U2792 : INV_X1 port map( A => datapath_i_alu_output_val_i_2_port, ZN => 
                           n5996);
   U2793 : OAI22_X1 port map( A1 => n5386, A2 => n5361, B1 => n5996, B2 => 
                           n6220, ZN => n5997);
   U2794 : AOI21_X1 port map( B1 => n5094, B2 => n4955, A => n5997, ZN => n5921
                           );
   U2795 : INV_X1 port map( A => n5921, ZN => n6205);
   U2796 : AOI22_X1 port map( A1 => n4956, A2 => n5385, B1 => n5408, B2 => 
                           n6205, ZN => n6207);
   U2797 : INV_X1 port map( A => n6207, ZN => n5896);
   U2798 : AOI22_X1 port map( A1 => n5094, A2 => n5083, B1 => 
                           datapath_i_alu_output_val_i_3_port, B2 => n5286, ZN 
                           => n5998);
   U2799 : OAI21_X1 port map( B1 => n5386, B2 => n5337, A => n5998, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U2800 : NAND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_3_port,
                           A2 => n6205, ZN => n6118);
   U2801 : OAI211_X1 port map( C1 => n6205, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n5408, B => n6118, ZN => n5999);
   U2802 : NAND2_X1 port map( A1 => n4972, A2 => n5999, ZN => n6209);
   U2803 : INV_X1 port map( A => n6209, ZN => n5895);
   U2804 : AOI22_X1 port map( A1 => n5359, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n5094, B2 
                           => n5054, ZN => n6000);
   U2805 : OAI21_X1 port map( B1 => n5386, B2 => n5328, A => n6000, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U2806 : INV_X1 port map( A => n6118, ZN => n6001);
   U2807 : NAND2_X1 port map( A1 => n6001, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n6010);
   U2808 : OAI211_X1 port map( C1 => n6001, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n5408, B => n6010, ZN => n6002);
   U2809 : NAND2_X1 port map( A1 => n4971, A2 => n6002, ZN => n6113);
   U2810 : INV_X1 port map( A => n6113, ZN => n5898);
   U2811 : AOI22_X1 port map( A1 => n5094, A2 => n5055, B1 => n5286, B2 => 
                           datapath_i_alu_output_val_i_1_port, ZN => n6003);
   U2812 : OAI21_X1 port map( B1 => n5386, B2 => n5355, A => n6003, ZN => n5478
                           );
   U2813 : AOI22_X1 port map( A1 => n5385, A2 => IRAM_ADDRESS_1_port, B1 => 
                           n5478, B2 => n6219, ZN => n5919);
   U2814 : AOI21_X1 port map( B1 => datapath_i_alu_output_val_i_5_port, B2 => 
                           n6216, A => n6223, ZN => n5943);
   U2815 : AOI22_X1 port map( A1 => n5359, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n5094, B2 
                           => n5096, ZN => n6004);
   U2816 : OAI21_X1 port map( B1 => n5386, B2 => n5331, A => n6004, ZN => n1453
                           );
   U2817 : NOR2_X1 port map( A1 => n5943, A2 => n6010, ZN => n6009);
   U2818 : NAND2_X1 port map( A1 => n6009, A2 => n1453, ZN => n6035);
   U2819 : OAI211_X1 port map( C1 => n6009, C2 => n1453, A => n5408, B => n6035
                           , ZN => n6005);
   U2820 : NAND2_X1 port map( A1 => n4970, A2 => n6005, ZN => n6096);
   U2821 : INV_X1 port map( A => n6096, ZN => n5897);
   U2822 : AOI222_X1 port map( A1 => n5507, A2 => n6215, B1 => n5359, B2 => 
                           datapath_i_alu_output_val_i_7_port, C1 => n5320, C2 
                           => n5334, ZN => n5941);
   U2823 : INV_X1 port map( A => datapath_i_alu_output_val_i_8_port, ZN => 
                           n6006);
   U2824 : OAI222_X1 port map( A1 => n6006, A2 => n5382, B1 => n5383, B2 => 
                           n5425, C1 => n5423, C2 => n5386, ZN => n1449);
   U2825 : NOR2_X1 port map( A1 => n5941, A2 => n6035, ZN => n6034);
   U2826 : NAND2_X1 port map( A1 => n6034, A2 => n1449, ZN => n6061);
   U2827 : OAI211_X1 port map( C1 => n6034, C2 => n1449, A => n5408, B => n6061
                           , ZN => n6007);
   U2828 : NAND2_X1 port map( A1 => n4969, A2 => n6007, ZN => n6105);
   U2829 : INV_X1 port map( A => n6105, ZN => n5893);
   U2830 : AOI22_X1 port map( A1 => n5359, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n5094, B2 
                           => n5007, ZN => n6008);
   U2831 : OAI21_X1 port map( B1 => n5386, B2 => n5352, A => n6008, ZN => n5479
                           );
   U2832 : AOI22_X1 port map( A1 => n5385, A2 => IRAM_ADDRESS_0_port, B1 => 
                           n5479, B2 => n6219, ZN => n5918);
   U2833 : AOI211_X1 port map( C1 => n5943, C2 => n6010, A => n5385, B => n6009
                           , ZN => n6011);
   U2834 : NOR2_X1 port map( A1 => n4986, A2 => n6011, ZN => n5920);
   U2835 : OAI21_X1 port map( B1 => n6013, B2 => n6012, A => n6178, ZN => 
                           cu_i_cmd_word_6_port);
   U2836 : OR2_X1 port map( A1 => n4187, A2 => cu_i_cmd_word_6_port, ZN => 
                           cu_i_n135);
   U2837 : INV_X1 port map( A => n6017, ZN => n6015);
   U2838 : AOI22_X1 port map( A1 => n5388, A2 => cu_i_cmd_alu_op_type_1_port, 
                           B1 => n5461, B2 => n5129, ZN => n6018);
   U2839 : AOI21_X1 port map( B1 => n6019, B2 => n6021, A => n6017, ZN => n6014
                           );
   U2840 : OAI211_X1 port map( C1 => n6021, C2 => n6018, A => n6015, B => n6019
                           , ZN => n6016);
   U2841 : INV_X1 port map( A => n6016, ZN => n5860);
   U2842 : AOI21_X1 port map( B1 => n6019, B2 => n6018, A => n6017, ZN => n6020
                           );
   U2843 : AOI222_X1 port map( A1 => n5506, A2 => n6215, B1 => n5359, B2 => 
                           datapath_i_alu_output_val_i_9_port, C1 => n5317, C2 
                           => n5334, ZN => n5942);
   U2844 : INV_X1 port map( A => datapath_i_alu_output_val_i_10_port, ZN => 
                           n6022);
   U2845 : OAI222_X1 port map( A1 => n6022, A2 => n5382, B1 => n5383, B2 => 
                           n5422, C1 => n5420, C2 => n5386, ZN => n1447);
   U2846 : NOR2_X1 port map( A1 => n5942, A2 => n6061, ZN => n6060);
   U2847 : NAND2_X1 port map( A1 => n6060, A2 => n1447, ZN => n6082);
   U2848 : OAI211_X1 port map( C1 => n6060, C2 => n1447, A => n5408, B => n6082
                           , ZN => n6023);
   U2849 : NAND2_X1 port map( A1 => n4968, A2 => n6023, ZN => n6103);
   U2850 : INV_X1 port map( A => n6103, ZN => n5894);
   U2851 : AOI221_X1 port map( B1 => n5350, B2 => n5874, C1 => cu_i_n135, C2 =>
                           n3555, A => n5360, ZN => n4337);
   U2852 : OAI211_X1 port map( C1 => n5120, C2 => n5341, A => n5119, B => n5407
                           , ZN => n6024);
   U2853 : NAND2_X1 port map( A1 => n4965, A2 => n6024, ZN => n6066);
   U2854 : INV_X1 port map( A => n6066, ZN => n5906);
   U2855 : NAND2_X1 port map( A1 => n4992, A2 => n4966, ZN => n6101);
   U2856 : INV_X1 port map( A => n6101, ZN => n5945);
   U2857 : OR2_X1 port map( A1 => curr_instruction_to_cu_i_16_port, A2 => n5876
                           , ZN => n6025);
   U2858 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_20_port, A2 => 
                           curr_instruction_to_cu_i_17_port, A3 => 
                           curr_instruction_to_cu_i_19_port, A4 => n6025, ZN =>
                           n6027);
   U2859 : OAI22_X1 port map( A1 => n6028, A2 => n6027, B1 => n5880, B2 => 
                           n6026, ZN => n6033);
   U2860 : NOR4_X1 port map( A1 => n3229, A2 => n3227, A3 => n3231, A4 => n3233
                           , ZN => n6031);
   U2861 : AOI211_X1 port map( C1 => n5086, C2 => n4990, A => n6029, B => 
                           cu_i_n135, ZN => n6030);
   U2862 : OAI221_X1 port map( B1 => n5881, B2 => n6179, C1 => n5881, C2 => 
                           n6031, A => n6030, ZN => n6032);
   U2863 : AOI21_X1 port map( B1 => n6218, B2 => n6033, A => n6032, ZN => n4052
                           );
   U2864 : OR2_X1 port map( A1 => n4052, A2 => n5336, ZN => n5512);
   U2865 : AOI211_X1 port map( C1 => n5941, C2 => n6035, A => n5385, B => n6034
                           , ZN => n6036);
   U2866 : OR2_X1 port map( A1 => n4987, A2 => n6036, ZN => n5502);
   U2867 : CLKBUF_X1 port map( A => n5093, Z => n6228);
   U2868 : AOI211_X1 port map( C1 => n5379, C2 => n6038, A => n5384, B => n6037
                           , ZN => n6039);
   U2869 : OR2_X1 port map( A1 => n4976, A2 => n6039, ZN => n5936);
   U2870 : AOI211_X1 port map( C1 => n5381, C2 => n6041, A => n5384, B => n6040
                           , ZN => n6042);
   U2871 : OR2_X1 port map( A1 => n4975, A2 => n6042, ZN => n5938);
   U2872 : AOI211_X1 port map( C1 => n5377, C2 => n6044, A => n5384, B => n6043
                           , ZN => n6045);
   U2873 : OR2_X1 port map( A1 => n4977, A2 => n6045, ZN => n5934);
   U2874 : AOI211_X1 port map( C1 => n5375, C2 => n6047, A => n5384, B => n6046
                           , ZN => n6048);
   U2875 : OR2_X1 port map( A1 => n4978, A2 => n6048, ZN => n5932);
   U2876 : AOI211_X1 port map( C1 => n5369, C2 => n6050, A => n5384, B => n6049
                           , ZN => n6051);
   U2877 : OR2_X1 port map( A1 => n4981, A2 => n6051, ZN => n5926);
   U2878 : AOI211_X1 port map( C1 => n5365, C2 => n6053, A => n5384, B => n6052
                           , ZN => n6054);
   U2879 : OR2_X1 port map( A1 => n4979, A2 => n6054, ZN => n5930);
   U2880 : AOI211_X1 port map( C1 => n5367, C2 => n6056, A => n5384, B => n6055
                           , ZN => n6057);
   U2881 : OR2_X1 port map( A1 => n4980, A2 => n6057, ZN => n5928);
   U2882 : AOI211_X1 port map( C1 => n5119, C2 => n5373, A => n5384, B => n6058
                           , ZN => n6059);
   U2883 : OR2_X1 port map( A1 => n4982, A2 => n6059, ZN => n5924);
   U2884 : AOI211_X1 port map( C1 => n5942, C2 => n6061, A => n5385, B => n6060
                           , ZN => n6062);
   U2885 : OR2_X1 port map( A1 => n4985, A2 => n6062, ZN => n5501);
   U2886 : AOI211_X1 port map( C1 => n5121, C2 => n5371, A => n5384, B => n5120
                           , ZN => n6063);
   U2887 : OR2_X1 port map( A1 => n4983, A2 => n6063, ZN => n5922);
   U2888 : OR2_X1 port map( A1 => n5428, A2 => n5123, ZN => cu_i_N278);
   U2889 : INV_X1 port map( A => n5484, ZN => IRAM_ADDRESS_14_port);
   U2890 : INV_X1 port map( A => n5485, ZN => IRAM_ADDRESS_16_port);
   U2891 : INV_X1 port map( A => n5486, ZN => IRAM_ADDRESS_18_port);
   U2892 : INV_X1 port map( A => n5483, ZN => IRAM_ADDRESS_20_port);
   U2893 : INV_X1 port map( A => n5481, ZN => IRAM_ADDRESS_22_port);
   U2894 : INV_X1 port map( A => n5487, ZN => IRAM_ADDRESS_24_port);
   U2895 : INV_X1 port map( A => n5488, ZN => IRAM_ADDRESS_26_port);
   U2896 : INV_X1 port map( A => n5489, ZN => IRAM_ADDRESS_28_port);
   U2897 : INV_X1 port map( A => n5482, ZN => IRAM_ADDRESS_30_port);
   U2898 : INV_X1 port map( A => n5869, ZN => n6064);
   U2899 : NAND2_X1 port map( A1 => n5439, A2 => n6064, ZN => n3261);
   U2900 : OAI21_X1 port map( B1 => n5098, B2 => n5319, A => n4989, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U2901 : AOI22_X1 port map( A1 => n5242, A2 => n5387, B1 => n5097, B2 => 
                           n5508, ZN => n6065);
   U2902 : MUX2_X1 port map( A => n5013, B => n5142, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U2903 : MUX2_X1 port map( A => n5020, B => n5136, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U2904 : MUX2_X1 port map( A => n5011, B => n5148, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U2905 : MUX2_X1 port map( A => n5012, B => n5145, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U2906 : NOR2_X1 port map( A1 => n5439, A2 => n5869, ZN => n3241);
   U2907 : AOI22_X1 port map( A1 => n5097, A2 => n6066, B1 => n5409, B2 => 
                           n5248, ZN => n6067);
   U2908 : OAI21_X1 port map( B1 => n5098, B2 => n5431, A => n6067, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U2909 : AOI22_X1 port map( A1 => n5097, A2 => n5924, B1 => n5387, B2 => 
                           n5250, ZN => n6068);
   U2910 : OAI21_X1 port map( B1 => n5098, B2 => n5311, A => n6068, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U2911 : AOI22_X1 port map( A1 => n5097, A2 => n5928, B1 => n5409, B2 => 
                           n5258, ZN => n6069);
   U2912 : OAI21_X1 port map( B1 => n5098, B2 => n5305, A => n6069, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U2913 : MUX2_X1 port map( A => IRAM_DATA(23), B => n5079, S => n5388, Z => 
                           n3205);
   U2914 : NAND2_X1 port map( A1 => n5116, A2 => n5874, ZN => n6070);
   U2915 : OAI21_X1 port map( B1 => n5460, B2 => n5874, A => n6070, ZN => n4133
                           );
   U2916 : AOI222_X1 port map( A1 => n5922, A2 => n6215, B1 => n5286, B2 => 
                           datapath_i_alu_output_val_i_13_port, C1 => n5312, C2
                           => n5334, ZN => n5923);
   U2917 : AOI222_X1 port map( A1 => n5508, A2 => n6215, B1 => n5334, B2 => 
                           n5315, C1 => n5359, C2 => 
                           datapath_i_alu_output_val_i_11_port, ZN => n5940);
   U2918 : INV_X1 port map( A => datapath_i_alu_output_val_i_12_port, ZN => 
                           n6071);
   U2919 : OAI222_X1 port map( A1 => n6071, A2 => n5382, B1 => n5383, B2 => 
                           n5945, C1 => n5433, C2 => n5386, ZN => n1445);
   U2920 : NOR2_X1 port map( A1 => n5940, A2 => n6082, ZN => n6081);
   U2921 : NAND2_X1 port map( A1 => n6081, A2 => n1445, ZN => n4231);
   U2922 : NOR2_X1 port map( A1 => n5923, A2 => n4231, ZN => n4230);
   U2923 : INV_X1 port map( A => datapath_i_alu_output_val_i_14_port, ZN => 
                           n6072);
   U2924 : OAI222_X1 port map( A1 => n6072, A2 => n5389, B1 => n5386, B2 => 
                           n5431, C1 => n5906, C2 => n5383, ZN => n1443);
   U2925 : NAND2_X1 port map( A1 => n4230, A2 => n1443, ZN => n4228);
   U2926 : INV_X1 port map( A => datapath_i_alu_output_val_i_16_port, ZN => 
                           n6073);
   U2927 : OAI222_X1 port map( A1 => n6073, A2 => n5389, B1 => n5386, B2 => 
                           n5444, C1 => n5908, C2 => n5383, ZN => n1441);
   U2928 : INV_X1 port map( A => datapath_i_alu_output_val_i_18_port, ZN => 
                           n6074);
   U2929 : OAI222_X1 port map( A1 => n6074, A2 => n5389, B1 => n5386, B2 => 
                           n5442, C1 => n5907, C2 => n5383, ZN => n1439);
   U2930 : OAI211_X1 port map( C1 => n6081, C2 => n1445, A => n5408, B => n4231
                           , ZN => n4155);
   U2931 : INV_X1 port map( A => datapath_i_alu_output_val_i_20_port, ZN => 
                           n6075);
   U2932 : OAI222_X1 port map( A1 => n6075, A2 => n5389, B1 => n5386, B2 => 
                           n5429, C1 => n5905, C2 => n5383, ZN => n1437);
   U2933 : INV_X1 port map( A => datapath_i_alu_output_val_i_22_port, ZN => 
                           n6076);
   U2934 : OAI222_X1 port map( A1 => n6076, A2 => n5389, B1 => n5386, B2 => 
                           n5426, C1 => n5904, C2 => n5383, ZN => n1435);
   U2935 : INV_X1 port map( A => datapath_i_alu_output_val_i_24_port, ZN => 
                           n6077);
   U2936 : OAI222_X1 port map( A1 => n6077, A2 => n5389, B1 => n5386, B2 => 
                           n5418, C1 => n5903, C2 => n5383, ZN => n1433);
   U2937 : INV_X1 port map( A => datapath_i_alu_output_val_i_26_port, ZN => 
                           n6078);
   U2938 : OAI222_X1 port map( A1 => n6078, A2 => n5389, B1 => n5386, B2 => 
                           n5416, C1 => n5902, C2 => n5383, ZN => n1431);
   U2939 : INV_X1 port map( A => datapath_i_alu_output_val_i_28_port, ZN => 
                           n6079);
   U2940 : OAI222_X1 port map( A1 => n6079, A2 => n5389, B1 => n5386, B2 => 
                           n5414, C1 => n5901, C2 => n5383, ZN => n1429);
   U2941 : INV_X1 port map( A => datapath_i_alu_output_val_i_30_port, ZN => 
                           n6080);
   U2942 : OAI222_X1 port map( A1 => n6080, A2 => n5389, B1 => n5386, B2 => 
                           n5412, C1 => n5900, C2 => n5383, ZN => n1427);
   U2943 : INV_X1 port map( A => n5920, ZN => n6109);
   U2944 : AOI22_X1 port map( A1 => n5335, A2 => n6221, B1 => n5095, B2 => 
                           n6109, ZN => n4193);
   U2945 : AOI211_X1 port map( C1 => n5940, C2 => n6082, A => n5385, B => n6081
                           , ZN => n6083);
   U2946 : NOR2_X1 port map( A1 => n4984, A2 => n6083, ZN => n4128);
   U2947 : MUX2_X1 port map( A => n5010, B => n5151, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U2948 : AOI22_X1 port map( A1 => n5278, A2 => n5409, B1 => n5392, B2 => 
                           n5938, ZN => n6084);
   U2949 : OAI21_X1 port map( B1 => n5098, B2 => n5290, A => n6084, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U2950 : AOI22_X1 port map( A1 => n5097, A2 => n6085, B1 => n5387, B2 => 
                           n5280, ZN => n6086);
   U2951 : OAI21_X1 port map( B1 => n5098, B2 => n5412, A => n6086, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U2952 : AOI22_X1 port map( A1 => n5387, A2 => n5276, B1 => n5392, B2 => 
                           n6087, ZN => n6088);
   U2953 : OAI21_X1 port map( B1 => n5098, B2 => n5414, A => n6088, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U2954 : AOI22_X1 port map( A1 => n5097, A2 => n6089, B1 => n5387, B2 => 
                           n5272, ZN => n6090);
   U2955 : OAI21_X1 port map( B1 => n5098, B2 => n5416, A => n6090, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U2956 : AOI22_X1 port map( A1 => n5097, A2 => n5934, B1 => n5409, B2 => 
                           n5270, ZN => n6091);
   U2957 : OAI21_X1 port map( B1 => n5098, B2 => n5296, A => n6091, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U2958 : AOI22_X1 port map( A1 => n5097, A2 => n6092, B1 => n5409, B2 => 
                           n5268, ZN => n6093);
   U2959 : OAI21_X1 port map( B1 => n5098, B2 => n5418, A => n6093, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U2960 : AOI22_X1 port map( A1 => n5097, A2 => n6094, B1 => n5387, B2 => 
                           n5256, ZN => n6095);
   U2961 : OAI21_X1 port map( B1 => n5098, B2 => n5442, A => n6095, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U2962 : AOI22_X1 port map( A1 => n5869, A2 => n5237, B1 => n3241, B2 => 
                           n6096, ZN => n6097);
   U2963 : OAI21_X1 port map( B1 => n5332, B2 => n3261, A => n6097, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);
   U2964 : AOI22_X1 port map( A1 => n5869, A2 => n5238, B1 => n3241, B2 => 
                           n5502, ZN => n6098);
   U2965 : OAI21_X1 port map( B1 => n5517, B2 => n3261, A => n6098, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U2966 : AOI22_X1 port map( A1 => n5869, A2 => n5240, B1 => n3241, B2 => 
                           n5501, ZN => n4268);
   U2967 : AOI22_X1 port map( A1 => n5097, A2 => n6099, B1 => n5409, B2 => 
                           n5252, ZN => n6100);
   U2968 : OAI21_X1 port map( B1 => n5098, B2 => n5444, A => n6100, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U2969 : AOI22_X1 port map( A1 => n5244, A2 => n5409, B1 => n5392, B2 => 
                           n6101, ZN => n6102);
   U2970 : OAI21_X1 port map( B1 => n5433, B2 => n5098, A => n6102, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U2971 : AOI22_X1 port map( A1 => n5241, A2 => n5869, B1 => n3241, B2 => 
                           n6103, ZN => n4280);
   U2972 : NOR2_X1 port map( A1 => n5539, A2 => n6224, ZN => n6141);
   U2973 : INV_X1 port map( A => n6141, ZN => n6143);
   U2974 : NOR2_X1 port map( A1 => n6143, A2 => n6225, ZN => n6142);
   U2975 : NOR2_X1 port map( A1 => n6142, A2 => n5540, ZN => n6104);
   U2976 : AOI211_X1 port map( C1 => n6142, C2 => n5540, A => n5117, B => n6104
                           , ZN => cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U2978 : AOI22_X1 port map( A1 => n5869, A2 => n5239, B1 => n3241, B2 => 
                           n6105, ZN => n6106);
   U2979 : OAI21_X1 port map( B1 => n5424, B2 => n3261, A => n6106, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U2980 : INV_X1 port map( A => n5919, ZN => n6107);
   U2981 : AOI22_X1 port map( A1 => n5869, A2 => n5232, B1 => n3241, B2 => 
                           n6107, ZN => n6108);
   U2982 : OAI21_X1 port map( B1 => n5356, B2 => n3261, A => n6108, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U2983 : AOI22_X1 port map( A1 => n5869, A2 => n5236, B1 => n3241, B2 => 
                           n6109, ZN => n6110);
   U2984 : OAI21_X1 port map( B1 => n5503, B2 => n3261, A => n6110, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U2985 : AOI22_X1 port map( A1 => n5387, A2 => n5260, B1 => n5392, B2 => 
                           n6111, ZN => n6112);
   U2986 : OAI21_X1 port map( B1 => n5098, B2 => n5429, A => n6112, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U2987 : MUX2_X1 port map( A => n5014, B => n5139, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U2988 : AOI22_X1 port map( A1 => n5869, A2 => n5235, B1 => n3241, B2 => 
                           n6113, ZN => n6114);
   U2989 : OAI21_X1 port map( B1 => n5329, B2 => n3261, A => n6114, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U2990 : AOI22_X1 port map( A1 => n3555, A2 => cu_i_cmd_word_6_port, B1 => 
                           n5074, B2 => n5874, ZN => n6117);
   U2991 : AOI22_X1 port map( A1 => n3555, A2 => n4187, B1 => n5323, B2 => 
                           n5874, ZN => n6115);
   U2992 : NAND2_X1 port map( A1 => n5084, A2 => n6115, ZN => n6116);
   U2993 : OAI22_X1 port map( A1 => n6117, A2 => n6116, B1 => n5084, B2 => 
                           n6115, ZN => n5870);
   U2994 : NOR2_X1 port map( A1 => n5870, A2 => n5462, ZN => n3257);
   U2995 : NAND2_X1 port map( A1 => n5087, A2 => n4052, ZN => n3252);
   U2996 : NOR2_X1 port map( A1 => n6118, A2 => n5865, ZN => n6152);
   U2997 : NAND2_X1 port map( A1 => n6152, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n6151);
   U2998 : NOR2_X1 port map( A1 => n5943, A2 => n6151, ZN => n6154);
   U2999 : NAND2_X1 port map( A1 => n6154, A2 => n1453, ZN => n6153);
   U3000 : NOR2_X1 port map( A1 => n5941, A2 => n6153, ZN => n6156);
   U3001 : AOI211_X1 port map( C1 => n5941, C2 => n6153, A => n6156, B => n5946
                           , ZN => n3148);
   U3002 : AOI211_X1 port map( C1 => n5943, C2 => n6151, A => n6154, B => n5946
                           , ZN => n3147);
   U3003 : NAND2_X1 port map( A1 => n6156, A2 => n1449, ZN => n6155);
   U3004 : NOR2_X1 port map( A1 => n5942, A2 => n6155, ZN => n6158);
   U3005 : AOI211_X1 port map( C1 => n5942, C2 => n6155, A => n6158, B => n5946
                           , ZN => n3146);
   U3006 : NAND2_X1 port map( A1 => n6158, A2 => n1447, ZN => n6157);
   U3007 : NOR2_X1 port map( A1 => n5940, A2 => n6157, ZN => n6159);
   U3008 : AOI211_X1 port map( C1 => n5940, C2 => n6157, A => n6159, B => n5946
                           , ZN => n3145);
   U3009 : NAND2_X1 port map( A1 => n6159, A2 => n1445, ZN => n4341);
   U3010 : NOR2_X1 port map( A1 => n5923, A2 => n4341, ZN => n4344);
   U3011 : AOI211_X1 port map( C1 => n5091, C2 => n5370, A => n5090, B => n5408
                           , ZN => n3144);
   U3012 : NAND2_X1 port map( A1 => n5090, A2 => n5341, ZN => n6160);
   U3013 : NOR2_X1 port map( A1 => n5372, A2 => n6160, ZN => n6162);
   U3014 : AOI211_X1 port map( C1 => n5372, C2 => n6160, A => n6162, B => n5408
                           , ZN => n3143);
   U3015 : NAND2_X1 port map( A1 => n5342, A2 => n6162, ZN => n6161);
   U3016 : NOR2_X1 port map( A1 => n5368, A2 => n6161, ZN => n6164);
   U3017 : AOI211_X1 port map( C1 => n5368, C2 => n6161, A => n6164, B => n5408
                           , ZN => n3142);
   U3018 : NAND2_X1 port map( A1 => n5343, A2 => n6164, ZN => n6163);
   U3019 : NOR2_X1 port map( A1 => n5366, A2 => n6163, ZN => n6166);
   U3020 : AOI211_X1 port map( C1 => n5366, C2 => n6163, A => n6166, B => n5408
                           , ZN => n3141);
   U3021 : NAND2_X1 port map( A1 => n5344, A2 => n6166, ZN => n6165);
   U3022 : NOR2_X1 port map( A1 => n5364, A2 => n6165, ZN => n6168);
   U3023 : AOI211_X1 port map( C1 => n5364, C2 => n6165, A => n6168, B => n5408
                           , ZN => n3140);
   U3024 : NAND2_X1 port map( A1 => n5345, A2 => n6168, ZN => n6167);
   U3025 : NOR2_X1 port map( A1 => n5374, A2 => n6167, ZN => n6170);
   U3026 : AOI211_X1 port map( C1 => n5374, C2 => n6167, A => n6170, B => n5408
                           , ZN => n3139);
   U3027 : NAND2_X1 port map( A1 => n5346, A2 => n6170, ZN => n6169);
   U3028 : NOR2_X1 port map( A1 => n5376, A2 => n6169, ZN => n6172);
   U3029 : AOI211_X1 port map( C1 => n5376, C2 => n6169, A => n6172, B => n5408
                           , ZN => n3138);
   U3030 : NAND2_X1 port map( A1 => n5347, A2 => n6172, ZN => n6171);
   U3031 : NOR2_X1 port map( A1 => n5378, A2 => n6171, ZN => n6174);
   U3032 : AOI211_X1 port map( C1 => n5378, C2 => n6171, A => n6174, B => n5408
                           , ZN => n3137);
   U3033 : NAND2_X1 port map( A1 => n5348, A2 => n6174, ZN => n6173);
   U3034 : NOR2_X1 port map( A1 => n5380, A2 => n6173, ZN => n6175);
   U3035 : AOI211_X1 port map( C1 => n5380, C2 => n6173, A => n6175, B => n5408
                           , ZN => n3136);
   U3036 : AOI22_X1 port map( A1 => n3555, A2 => n301, B1 => n5428, B2 => n5874
                           , ZN => n3135);
   U3037 : INV_X1 port map( A => datapath_i_alu_output_val_i_31_port, ZN => 
                           n6119);
   U3038 : OAI222_X1 port map( A1 => n5899, A2 => n5383, B1 => n6119, B2 => 
                           n5382, C1 => n5386, C2 => n5410, ZN => n3692);
   U3039 : NOR2_X1 port map( A1 => n5076, A2 => n4995, ZN => n6120);
   U3040 : NAND2_X1 port map( A1 => n5449, A2 => n6120, ZN => n6121);
   U3041 : NOR2_X1 port map( A1 => n5077, A2 => n6121, ZN => n6136);
   U3042 : NOR2_X1 port map( A1 => n5509, A2 => n5078, ZN => n6133);
   U3043 : NAND2_X1 port map( A1 => n5088, A2 => n6227, ZN => n6128);
   U3044 : INV_X1 port map( A => n6121, ZN => n6122);
   U3045 : NAND3_X1 port map( A1 => n5077, A2 => n5532, A3 => n6122, ZN => 
                           n6140);
   U3046 : INV_X1 port map( A => n6136, ZN => n6123);
   U3047 : OAI211_X1 port map( C1 => n5532, C2 => n6128, A => n6140, B => n6123
                           , ZN => n6124);
   U3048 : AOI22_X1 port map( A1 => n6136, A2 => n5089, B1 => n6133, B2 => 
                           n6124, ZN => n6127);
   U3049 : NAND3_X1 port map( A1 => n5454, A2 => n5534, A3 => n6226, ZN => 
                           n6126);
   U3050 : NAND2_X1 port map( A1 => n5448, A2 => n5075, ZN => n6125);
   U3051 : NAND4_X1 port map( A1 => n4954, A2 => n6127, A3 => n6126, A4 => 
                           n6125, ZN => cu_i_N264);
   U3052 : NOR2_X1 port map( A1 => n6128, A2 => n5449, ZN => n6129);
   U3053 : AOI21_X1 port map( B1 => n6129, B2 => n6133, A => n5075, ZN => n6138
                           );
   U3054 : NOR3_X1 port map( A1 => n5340, A2 => n5457, A3 => n6140, ZN => n6132
                           );
   U3055 : NAND3_X1 port map( A1 => n5454, A2 => n5504, A3 => n5537, ZN => 
                           n6130);
   U3056 : NAND2_X1 port map( A1 => n6130, A2 => n5115, ZN => n6131);
   U3057 : AOI211_X1 port map( C1 => n5534, C2 => n5511, A => n6132, B => n6131
                           , ZN => n6135);
   U3058 : NAND3_X1 port map( A1 => n5532, A2 => n6136, A3 => n6133, ZN => 
                           n6134);
   U3059 : NAND3_X1 port map( A1 => n6138, A2 => n6135, A3 => n6134, ZN => 
                           cu_i_N265);
   U3060 : OAI221_X1 port map( B1 => n5089, B2 => n5532, C1 => n5089, C2 => 
                           n5078, A => n6136, ZN => n6139);
   U3061 : OAI221_X1 port map( B1 => n5504, B2 => n5448, C1 => n5504, C2 => 
                           n5538, A => n5511, ZN => n6137);
   U3062 : OAI211_X1 port map( C1 => n5509, C2 => n6139, A => n6138, B => n6137
                           , ZN => cu_i_N266);
   U3063 : OAI221_X1 port map( B1 => n6140, B2 => n5340, C1 => n6140, C2 => 
                           n5509, A => n5541, ZN => cu_i_N267);
   U3064 : NAND2_X1 port map( A1 => n5388, A2 => n5117, ZN => cu_i_N274);
   U3065 : AOI211_X1 port map( C1 => n5539, C2 => n6224, A => n5117, B => n6141
                           , ZN => cu_i_N275);
   U3066 : NOR2_X1 port map( A1 => n5117, A2 => n5131, ZN => cu_i_N273);
   U3067 : AOI211_X1 port map( C1 => n6143, C2 => n6225, A => n5117, B => n6142
                           , ZN => cu_i_N276);
   U3068 : AOI211_X1 port map( C1 => n5388, C2 => n5073, A => n5117, B => n5324
                           , ZN => cu_i_N279);
   U3069 : NOR2_X1 port map( A1 => n3238, A2 => n3236, ZN => n492);
   U3070 : NAND4_X1 port map( A1 => n6212, A2 => n6144, A3 => n5322, A4 => 
                           n6213, ZN => n6147);
   U3071 : INV_X1 port map( A => n5879, ZN => n6145);
   U3072 : NAND4_X1 port map( A1 => n6145, A2 => n3248, A3 => n492, A4 => n5891
                           , ZN => n6146);
   U3073 : OAI22_X1 port map( A1 => n6148, A2 => n6147, B1 => n6146, B2 => 
                           n5881, ZN => cu_i_cmd_word_8_port);
   U3074 : MUX2_X1 port map( A => n4973, B => cu_i_cmd_word_8_port, S => n3555,
                           Z => alu_cin_i);
   U3075 : MUX2_X1 port map( A => n5125, B => n5053, S => n3555, Z => n3211);
   U3076 : MUX2_X1 port map( A => n5126, B => n5052, S => n3555, Z => n3210);
   U3077 : MUX2_X1 port map( A => n4952, B => n5051, S => n3555, Z => n3209);
   U3078 : MUX2_X1 port map( A => IRAM_DATA(25), B => n5049, S => n5127, Z => 
                           n3207);
   U3079 : MUX2_X1 port map( A => IRAM_DATA(24), B => n5048, S => n5127, Z => 
                           n3206);
   U3080 : MUX2_X1 port map( A => IRAM_DATA(21), B => n5046, S => n5388, Z => 
                           n3203);
   U3081 : MUX2_X1 port map( A => IRAM_DATA(10), B => n5045, S => n5127, Z => 
                           n3202);
   U3082 : MUX2_X1 port map( A => IRAM_DATA(9), B => n5044, S => n5127, Z => 
                           n3201);
   U3083 : MUX2_X1 port map( A => IRAM_DATA(8), B => n5043, S => n5127, Z => 
                           n3200);
   U3084 : MUX2_X1 port map( A => IRAM_DATA(7), B => n5042, S => n5127, Z => 
                           n3199);
   U3085 : MUX2_X1 port map( A => IRAM_DATA(6), B => n5041, S => n5127, Z => 
                           n3198);
   U3086 : NOR2_X1 port map( A1 => n5921, A2 => n5865, ZN => n6150);
   U3087 : INV_X1 port map( A => n6152, ZN => n6149);
   U3088 : OAI211_X1 port map( C1 => n6150, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n5947, B => n6149, ZN => n3133);
   U3089 : OAI211_X1 port map( C1 => n6152, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n5947, B => n6151, ZN => n3132);
   U3090 : OAI211_X1 port map( C1 => n6154, C2 => n1453, A => n5947, B => n6153
                           , ZN => n3131);
   U3091 : OAI211_X1 port map( C1 => n6156, C2 => n1449, A => n5947, B => n6155
                           , ZN => n3130);
   U3092 : OAI211_X1 port map( C1 => n6158, C2 => n1447, A => n5947, B => n6157
                           , ZN => n3129);
   U3093 : OAI211_X1 port map( C1 => n6159, C2 => n1445, A => n5947, B => n4341
                           , ZN => n3128);
   U3094 : OAI211_X1 port map( C1 => n5090, C2 => IRAM_ADDRESS_14_port, A => 
                           n5385, B => n6160, ZN => n3127);
   U3095 : OAI211_X1 port map( C1 => n6162, C2 => IRAM_ADDRESS_16_port, A => 
                           n5385, B => n6161, ZN => n3126);
   U3096 : OAI211_X1 port map( C1 => n6164, C2 => IRAM_ADDRESS_18_port, A => 
                           n5385, B => n6163, ZN => n3125);
   U3097 : OAI211_X1 port map( C1 => n6166, C2 => IRAM_ADDRESS_20_port, A => 
                           n5385, B => n6165, ZN => n3124);
   U3098 : OAI211_X1 port map( C1 => n6168, C2 => IRAM_ADDRESS_22_port, A => 
                           n5385, B => n6167, ZN => n3123);
   U3099 : OAI211_X1 port map( C1 => n6170, C2 => IRAM_ADDRESS_24_port, A => 
                           n5385, B => n6169, ZN => n3122);
   U3100 : OAI211_X1 port map( C1 => n6172, C2 => IRAM_ADDRESS_26_port, A => 
                           n5385, B => n6171, ZN => n3121);
   U3101 : OAI211_X1 port map( C1 => n6174, C2 => IRAM_ADDRESS_28_port, A => 
                           n5385, B => n6173, ZN => n3120);
   U3102 : NAND2_X1 port map( A1 => n5349, A2 => n6175, ZN => n6176);
   U3103 : OAI211_X1 port map( C1 => n6175, C2 => IRAM_ADDRESS_30_port, A => 
                           n5385, B => n6176, ZN => n3119);
   U3104 : XOR2_X1 port map( A => n5465, B => n6176, Z => n3243);
   U3105 : AND2_X1 port map( A1 => n5428, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U3106 : OAI21_X1 port map( B1 => n6177, B2 => n5885, A => n6180, ZN => 
                           read_rf_p2_i);
   U3107 : OAI221_X1 port map( B1 => n6182, B2 => n6181, C1 => n6180, C2 => 
                           n6179, A => n6178, ZN => n3112);
   U3108 : OAI21_X1 port map( B1 => n5353, B2 => n6183, A => n5716, ZN => 
                           datapath_i_decode_stage_dp_n44);
   U3109 : OAI21_X1 port map( B1 => n5356, B2 => n6183, A => n5713, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U3110 : OAI21_X1 port map( B1 => n5362, B2 => n6183, A => n5712, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U3111 : OAI21_X1 port map( B1 => n5338, B2 => n6183, A => n5711, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U3112 : OAI21_X1 port map( B1 => n5329, B2 => n6183, A => n5710, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U3113 : OAI21_X1 port map( B1 => n6183, B2 => n5326, A => n5709, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U3114 : OAI21_X1 port map( B1 => n5332, B2 => n6183, A => n5708, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U3115 : OAI21_X1 port map( B1 => n6183, B2 => n5111, A => n5707, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U3116 : OAI21_X1 port map( B1 => n5424, B2 => n6183, A => n5706, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U3117 : OAI21_X1 port map( B1 => n5081, B2 => n5113, A => n5705, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U3118 : OAI21_X1 port map( B1 => n5081, B2 => n5421, A => n5704, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U3119 : OAI21_X1 port map( B1 => n6183, B2 => n5100, A => n5703, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U3120 : OAI21_X1 port map( B1 => n6183, B2 => n5434, A => n5702, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U3121 : OAI21_X1 port map( B1 => n5081, B2 => n5102, A => n5701, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U3122 : OAI21_X1 port map( B1 => n5081, B2 => n5432, A => n5700, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U3123 : OAI21_X1 port map( B1 => n6183, B2 => n5103, A => n5699, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U3124 : OAI21_X1 port map( B1 => n6183, B2 => n5445, A => n5698, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U3125 : OAI21_X1 port map( B1 => n5081, B2 => n5104, A => n5697, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U3126 : OAI21_X1 port map( B1 => n5081, B2 => n5443, A => n5696, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U3127 : OAI21_X1 port map( B1 => n6183, B2 => n5105, A => n5695, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U3128 : OAI21_X1 port map( B1 => n6183, B2 => n5430, A => n5694, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U3129 : OAI21_X1 port map( B1 => n5081, B2 => n5106, A => n5693, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U3130 : OAI21_X1 port map( B1 => n5081, B2 => n5427, A => n5692, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U3131 : OAI21_X1 port map( B1 => n6183, B2 => n5107, A => n5691, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U3132 : OAI21_X1 port map( B1 => n6183, B2 => n5419, A => n5690, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U3133 : OAI21_X1 port map( B1 => n5081, B2 => n5108, A => n5689, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U3134 : OAI21_X1 port map( B1 => n5081, B2 => n5417, A => n5688, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U3135 : OAI21_X1 port map( B1 => n6183, B2 => n5109, A => n5687, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U3136 : OAI21_X1 port map( B1 => n6183, B2 => n5415, A => n5686, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U3137 : OAI21_X1 port map( B1 => n5081, B2 => n5110, A => n5685, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U3138 : OAI21_X1 port map( B1 => n5081, B2 => n5413, A => n5684, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U3139 : OAI21_X1 port map( B1 => n6183, B2 => n5411, A => n5683, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U3140 : NOR4_X1 port map( A1 => n1641, A2 => n1643, A3 => n1645, A4 => n1647
                           , ZN => n6187);
   U3141 : NOR4_X1 port map( A1 => n1649, A2 => n1651, A3 => n1653, A4 => n1655
                           , ZN => n6186);
   U3142 : NOR4_X1 port map( A1 => n1625, A2 => n1627, A3 => n1629, A4 => n1631
                           , ZN => n6185);
   U3143 : NOR4_X1 port map( A1 => n1633, A2 => n1635, A3 => n1637, A4 => n1639
                           , ZN => n6184);
   U3144 : NAND4_X1 port map( A1 => n6187, A2 => n6186, A3 => n6185, A4 => 
                           n6184, ZN => n6193);
   U3145 : NOR4_X1 port map( A1 => n1663, A2 => n1617, A3 => n1619, A4 => n1621
                           , ZN => n6191);
   U3146 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1661
                           , ZN => n6190);
   U3147 : NOR4_X1 port map( A1 => n1667, A2 => n1669, A3 => n1657, A4 => n1659
                           , ZN => n6189);
   U3148 : NOR4_X1 port map( A1 => n1623, A2 => n1671, A3 => n1673, A4 => n1665
                           , ZN => n6188);
   U3149 : NAND4_X1 port map( A1 => n6191, A2 => n6190, A3 => n6189, A4 => 
                           n6188, ZN => n6192);
   U3150 : NOR2_X1 port map( A1 => n6193, A2 => n6192, ZN => n3242);
   U3151 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n5462, Z => n3197);
   U3152 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n5462, Z => n3196);
   U3153 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n5462, Z => n3195);
   U3154 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n5462, Z => n3194);
   U3155 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n5440, Z => n3193);
   U3156 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n5440, Z => n3192);
   U3157 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n5440, Z => n3191);
   U3158 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n5440, Z => n3190);
   U3159 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, S 
                           => n5440, Z => n3189);
   U3160 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, S 
                           => n5440, Z => n3188);
   U3161 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, S 
                           => n5440, Z => n3187);
   U3162 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, S 
                           => n5440, Z => n3186);
   U3163 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, S 
                           => n5440, Z => n3185);
   U3164 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, S 
                           => n5440, Z => n3184);
   U3165 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, S 
                           => n5462, Z => n3183);
   U3166 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, S 
                           => n5462, Z => n3182);
   U3167 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, S 
                           => n5462, Z => n3181);
   U3168 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, S 
                           => n5462, Z => n3180);
   U3169 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, S 
                           => n5462, Z => n3179);
   U3170 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, S 
                           => n5462, Z => n3178);
   U3171 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n5440, Z => n3177);
   U3172 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, S 
                           => n5440, Z => n3176);
   U3173 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, S 
                           => n5440, Z => n3175);
   U3174 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, S 
                           => n5440, Z => n3174);
   U3175 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, S 
                           => n5440, Z => n3173);
   U3176 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, S 
                           => n5440, Z => n3172);
   U3177 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n5440, Z => n3171);
   U3178 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n5440, Z => n3170);
   U3179 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n5440, Z => n3169);
   U3180 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n5440, Z => n3168);
   U3181 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n5440, Z => n3167);
   U3182 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n5462, Z => n3166);
   U3183 : MUX2_X1 port map( A => n5040, B => n5157, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U3184 : MUX2_X1 port map( A => n5039, B => n5160, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U3185 : MUX2_X1 port map( A => n5038, B => n5163, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U3186 : MUX2_X1 port map( A => n5037, B => n5166, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U3187 : MUX2_X1 port map( A => n5036, B => n5169, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U3188 : MUX2_X1 port map( A => n5035, B => n5172, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U3189 : MUX2_X1 port map( A => n5034, B => n5175, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U3190 : MUX2_X1 port map( A => n5033, B => n5178, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U3191 : MUX2_X1 port map( A => n5032, B => n5181, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U3192 : MUX2_X1 port map( A => n5031, B => n5184, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U3193 : MUX2_X1 port map( A => n5030, B => n5187, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U3194 : MUX2_X1 port map( A => n5029, B => n5190, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U3195 : MUX2_X1 port map( A => n5028, B => n5193, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U3196 : MUX2_X1 port map( A => n5027, B => n5196, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U3197 : MUX2_X1 port map( A => n5026, B => n5199, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U3198 : MUX2_X1 port map( A => n5025, B => n5202, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U3199 : MUX2_X1 port map( A => n5024, B => n5205, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U3200 : MUX2_X1 port map( A => n5023, B => n5208, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U3201 : MUX2_X1 port map( A => n5022, B => n5211, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U3202 : MUX2_X1 port map( A => n5021, B => n5214, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U3203 : MUX2_X1 port map( A => n5019, B => n5217, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U3204 : MUX2_X1 port map( A => n5018, B => n5220, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U3205 : MUX2_X1 port map( A => n5017, B => n5223, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U3206 : MUX2_X1 port map( A => n5016, B => n5226, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U3207 : MUX2_X1 port map( A => n5015, B => n5229, S => n5463, Z => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U3208 : MUX2_X1 port map( A => n5009, B => n5154, S => n4974, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U3209 : AOI22_X1 port map( A1 => n5097, A2 => n5922, B1 => n5387, B2 => 
                           n5246, ZN => n6194);
   U3210 : OAI21_X1 port map( B1 => n5098, B2 => n5314, A => n6194, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U3211 : AOI22_X1 port map( A1 => n5392, A2 => n5926, B1 => n5409, B2 => 
                           n5254, ZN => n6195);
   U3212 : OAI21_X1 port map( B1 => n5098, B2 => n5308, A => n6195, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U3213 : AOI22_X1 port map( A1 => n5097, A2 => n5930, B1 => n5387, B2 => 
                           n5262, ZN => n6196);
   U3214 : OAI21_X1 port map( B1 => n5098, B2 => n5302, A => n6196, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U3215 : AOI22_X1 port map( A1 => n5097, A2 => n6197, B1 => n5387, B2 => 
                           n5264, ZN => n6198);
   U3216 : OAI21_X1 port map( B1 => n5098, B2 => n5426, A => n6198, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U3217 : AOI22_X1 port map( A1 => n5392, A2 => n5932, B1 => n5409, B2 => 
                           n5266, ZN => n6199);
   U3218 : OAI21_X1 port map( B1 => n5098, B2 => n5299, A => n6199, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U3219 : INV_X1 port map( A => n5918, ZN => n6200);
   U3220 : AOI22_X1 port map( A1 => n5869, A2 => n5231, B1 => n3241, B2 => 
                           n6200, ZN => n6201);
   U3221 : OAI21_X1 port map( B1 => n5353, B2 => n3261, A => n6201, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U3222 : AOI22_X1 port map( A1 => n5097, A2 => n5936, B1 => n5387, B2 => 
                           n5274, ZN => n6202);
   U3223 : OAI21_X1 port map( B1 => n5098, B2 => n5293, A => n6202, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U3224 : AOI22_X1 port map( A1 => n6203, A2 => n5097, B1 => n5387, B2 => 
                           n5282, ZN => n6204);
   U3225 : OAI21_X1 port map( B1 => n5410, B2 => n5098, A => n6204, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U3226 : INV_X1 port map( A => n5865, ZN => n6206);
   U3227 : AOI22_X1 port map( A1 => n5921, A2 => n6206, B1 => n5865, B2 => 
                           n6205, ZN => n3161);
   U3228 : AOI22_X1 port map( A1 => n5869, A2 => n5233, B1 => n3241, B2 => 
                           n6207, ZN => n6208);
   U3229 : OAI21_X1 port map( B1 => n5362, B2 => n3261, A => n6208, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U3230 : AOI22_X1 port map( A1 => n5869, A2 => n5234, B1 => n3241, B2 => 
                           n6209, ZN => n6210);
   U3231 : OAI21_X1 port map( B1 => n5338, B2 => n3261, A => n6210, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U3232 : MUX2_X1 port map( A => n5051, B => n5006, S => n3555, Z => n3160);
   U3233 : AND4_X1 port map( A1 => n5436, A2 => n5438, A3 => n4953, A4 => n5435
                           , ZN => n6211);
   U3234 : NAND2_X1 port map( A1 => n5437, A2 => n6211, ZN => n3596);
   U3235 : OAI211_X1 port map( C1 => n5892, C2 => n5887, A => n6212, B => n6213
                           , ZN => n3239);
   U3236 : NAND2_X1 port map( A1 => n6213, A2 => n5887, ZN => n2299);
   U3237 : NOR2_X1 port map( A1 => n5870, A2 => n6217, ZN => n5505);
   U3238 : NOR2_X1 port map( A1 => n5087, A2 => n4052, ZN => n5513);
   U3239 : AOI222_X1 port map( A1 => n5938, A2 => n6215, B1 => n5286, B2 => 
                           datapath_i_alu_output_val_i_29_port, C1 => n5288, C2
                           => n5334, ZN => n5939);
   U3240 : AOI222_X1 port map( A1 => n5936, A2 => n6215, B1 => n5286, B2 => 
                           datapath_i_alu_output_val_i_27_port, C1 => n5291, C2
                           => n5334, ZN => n5937);
   U3241 : AOI222_X1 port map( A1 => n5934, A2 => n6215, B1 => n5286, B2 => 
                           datapath_i_alu_output_val_i_25_port, C1 => n5294, C2
                           => n5334, ZN => n5935);
   U3242 : AOI222_X1 port map( A1 => n5932, A2 => n6215, B1 => n5286, B2 => 
                           datapath_i_alu_output_val_i_23_port, C1 => n5297, C2
                           => n5334, ZN => n5933);
   U3243 : AOI222_X1 port map( A1 => n5930, A2 => n6215, B1 => n5334, B2 => 
                           n5300, C1 => datapath_i_alu_output_val_i_21_port, C2
                           => n5286, ZN => n5931);
   U3244 : AOI222_X1 port map( A1 => n5928, A2 => n6215, B1 => n5334, B2 => 
                           n5303, C1 => datapath_i_alu_output_val_i_19_port, C2
                           => n5286, ZN => n5929);
   U3245 : AOI222_X1 port map( A1 => n5926, A2 => n6215, B1 => n5334, B2 => 
                           n5306, C1 => datapath_i_alu_output_val_i_17_port, C2
                           => n5286, ZN => n5927);
   U3246 : AOI222_X1 port map( A1 => n5924, A2 => n6215, B1 => n5334, B2 => 
                           n5309, C1 => datapath_i_alu_output_val_i_15_port, C2
                           => n5286, ZN => n5925);
   U3247 : AOI22_X1 port map( A1 => n3555, A2 => n5050, B1 => n5122, B2 => 
                           n5874, ZN => n5875);
   U3248 : MUX2_X1 port map( A => n5351, B => n5285, S => n3555, Z => n5868);

end SYN_dlx_rtl;
