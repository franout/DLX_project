
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal DATA2_I_30_port, DATA2_I_28_port, DATA2_I_27_port, DATA2_I_26_port, 
      DATA2_I_25_port, DATA2_I_24_port, DATA2_I_23_port, DATA2_I_22_port, 
      DATA2_I_21_port, DATA2_I_20_port, DATA2_I_19_port, DATA2_I_18_port, 
      DATA2_I_17_port, DATA2_I_16_port, DATA2_I_15_port, DATA2_I_14_port, 
      DATA2_I_13_port, DATA2_I_12_port, DATA2_I_11_port, DATA2_I_10_port, 
      DATA2_I_9_port, DATA2_I_8_port, DATA2_I_7_port, DATA2_I_6_port, 
      DATA2_I_5_port, DATA2_I_4_port, DATA2_I_3_port, DATA2_I_2_port, 
      DATA2_I_1_port, DATA2_I_0_port, data1_mul_15_port, data1_mul_0_port, 
      data2_mul_2_port, data2_mul_1_port, N2517, N2518, N2519, N2520, N2521, 
      N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n554, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1429, 
      n2808, n3020, n3026, n3027, n3028, n3029, n3030, n3036, n3940, n3957, 
      n3958, n3973, n3974, n3990, n3991, n3992, n3993, n3994, n3995, n4007, 
      n4008, n4009, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4293, 
      n4295, n4302, n4395, n7769, n7822, n8626, n8732, n8733, n8734, n8735, 
      n8736, n8737, n8738, n8739, n8740, n8748, n8749, n8751, n8752, n8753, 
      n8754, n8755, n8764, n8847, n8928, n8978, n9045, n9048, n9051, n9054, 
      n9057, n9060, n9063, n9066, n9069, n9072, n9075, n9078, n9081, n9084, 
      n11449, n11966, n12313, n12526, n13151, n13848, n13854, n13855, n13856, 
      n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13867, n13868, 
      n13873, n13878, n13884, n13896, n13897, n13898, n13899, n13900, n13901, 
      n13902, n13903, n13904, n13906, n13907, n13908, n13910, n13912, n13913, 
      n13914, n13915, n13916, n13917, n13918, n13919, n13922, n13924, n13927, 
      n13928, n13929, n13930, n13931, n13932, n13933, n13935, n13936, n13938, 
      n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13949, 
      n13950, n13953, n13954, n13955, n13956, n13963, n13964, n13965, n13966, 
      n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13976, 
      n13977, n13978, n13980, n13984, n13985, n13987, n13988, n13989, n13990, 
      n13992, n13997, n13999, n14000, n14003, n14004, n14009, n14011, n14013, 
      n14015, n14017, n14019, n14022, n14023, n14026, n14029, n14032, n14035, 
      n14038, n14041, n14044, n14047, n14050, n14053, n14056, n14057, n14058, 
      n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, 
      n14068, n14070, n14074, n14075, n14076, n14077, n14078, n14080, n14085, 
      n14086, n14087, n14088, n14093, n14094, n14095, n14100, n14101, n14102, 
      n14103, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, 
      n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14132, n14140, 
      n14141, n14142, n14143, n14144, n14145, n14146, n14149, n14150, n14151, 
      n14152, n14154, n14155, n14157, n14158, n14159, n14160, n14161, n14163, 
      n14164, n14165, n14168, n14170, n14176, n14182, n14184, n14234, n14235, 
      n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, 
      n14245, n14246, n14247, n14248, n14249, n14251, n14252, n14253, n14259, 
      n14261, n14262, n14263, n14264, n14265, n14266, n14268, n14269, n14271, 
      n14272, n14273, n14278, n14281, n14285, n14286, n14287, n14288, n14290, 
      n14292, n14407, n14416, n14431, n14432, n14452, n1809, n1871, n1894, 
      n1896, n16695, n16696, n16698, n16700, n16702, n16705, n16706, n16709, 
      n16713, n16766, n16770, n16771, n16782, n16783, n16797, n16807, n16808, 
      n16831, n16857, n16909, n17011, n17012, n17016, n17017, n17018, n17019, 
      n17020, n17068, n17089, n17140, n17160, n17254, n17269, n17270, n17359, 
      n17360, n17388, n17471, n17479, n17503, n17504, n17505, n17506, n17527, 
      n17537, n17728, n17733, n17734, n17735, n17932, n17965, n17966, n17968, 
      n18051, n18133, n18195, n18199, n18839, n18840, n18841, n18842, n18843, 
      n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, 
      n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, 
      n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, 
      n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, 
      n18880, n18881, n18882, n18884, n18885, n18886, n18887, n18888, n18889, 
      n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, 
      n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18907, n18908, 
      n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, 
      n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, 
      n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, 
      n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, 
      n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, 
      n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, 
      n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, 
      n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, 
      n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, 
      n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, 
      n18999, n19000, n19001, n19003, n19004, n19005, n19006, n19007, n19008, 
      n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, 
      n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, 
      n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, 
      n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, 
      n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, 
      n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, 
      n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, 
      n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, 
      n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, 
      n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, 
      n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, 
      n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, 
      n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, 
      n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, 
      n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, 
      n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, 
      n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, 
      n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, 
      n19171, n19172, n19174, n19175, n19176, n19177, n19178, n19179, n19180, 
      n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, 
      n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, 
      n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, 
      n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, 
      n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, 
      n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, 
      n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, 
      n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, 
      n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, 
      n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, 
      n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, 
      n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, 
      n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19297, n19298, 
      n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, 
      n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, 
      n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, 
      n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, 
      n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, 
      n19344, n19345, n19346, n19347, n19348, n19349, n19352, n19353, n19354, 
      n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, 
      n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, 
      n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, 
      n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, 
      n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, 
      n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, 
      n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, 
      n19418, n19419, n19420, n19421, n19422, n19423, n19425, n19426, n19427, 
      n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, 
      n19437, n19439, n19440, n19441, n19442, n19443, n19444, n19446, n21157, 
      n21158, n21159, n21160, n21161, n21162, n21163, n21165, n21166, n21167, 
      n21168, n21169, n21170, n21171, n21172, n21174, n21175, n21176, n21177, 
      n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, 
      n21187, n21188, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
      n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1843, n1844, n1845, n1846, n1847, 
      n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, 
      n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, 
      n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, 
      n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, 
      n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, 
      n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, 
      n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, 
      n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, 
      n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, 
      n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, 
      n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, 
      n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, 
      n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, 
      n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, 
      n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, 
      n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, 
      n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, 
      n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, 
      n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, 
      n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, 
      n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, 
      n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, 
      n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, 
      n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, 
      n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, 
      n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, 
      n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, 
      n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, 
      n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, 
      n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, 
      n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, 
      n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, 
      n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, 
      n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, 
      n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, 
      n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, 
      n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, 
      n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, 
      n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, 
      n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, 
      n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, 
      n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, 
      n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, 
      n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, 
      n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, 
      n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, 
      n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, 
      n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, 
      n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, 
      n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, 
      n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, 
      n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, 
      n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, 
      n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, 
      n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, 
      n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, 
      n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, 
      n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, 
      n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, 
      n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, 
      n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, 
      n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, 
      n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, 
      n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, 
      n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, 
      n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, 
      n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, 
      n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, 
      n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, 
      n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, 
      n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, 
      n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, 
      n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, 
      n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, 
      n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, 
      n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, 
      n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, 
      n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, 
      n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, 
      n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, 
      n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, 
      n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, 
      n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, 
      n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, 
      n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, 
      n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, 
      n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, 
      n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, 
      n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, 
      n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, 
      n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, 
      n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, 
      n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, 
      n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, 
      n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, 
      n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, 
      n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, 
      n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, 
      n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, 
      n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, 
      n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, 
      n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, 
      n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, 
      n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, 
      n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, 
      n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, 
      n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, 
      n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, 
      n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, 
      n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, 
      n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, 
      n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, 
      n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, 
      n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, 
      n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, 
      n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, 
      n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, 
      n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, 
      n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, 
      n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, 
      n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, 
      n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, 
      n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, 
      n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, 
      n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, 
      n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, 
      n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, 
      n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, 
      n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, 
      n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, 
      n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, 
      n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, 
      n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, 
      n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, 
      n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, 
      n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, 
      n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, 
      n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, 
      n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, 
      n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, 
      n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, 
      n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, 
      n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, 
      n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, 
      n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, 
      n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, 
      n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, 
      n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, 
      n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, 
      n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, 
      n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, 
      n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, 
      n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, 
      n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, 
      n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, 
      n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, 
      n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, 
      n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, 
      n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, 
      n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, 
      n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, 
      n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, 
      n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, 
      n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, 
      n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, 
      n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, 
      n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, 
      n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, 
      n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, 
      n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, 
      n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, 
      n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, 
      n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, 
      n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, 
      n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, 
      n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, 
      n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, 
      n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, 
      n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, 
      n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, 
      n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, 
      n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, 
      n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, 
      n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, 
      n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, 
      n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, 
      n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, 
      n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, 
      n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, 
      n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, 
      n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, 
      n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, 
      n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, 
      n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, 
      n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, 
      n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, 
      n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, 
      n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, 
      n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, 
      n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, 
      n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, 
      n22998, n22999, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578 : std_logic;

begin
   
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n554, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n554, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n22999, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n554, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n554, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n22999, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n554, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n554, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n554, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n554, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n554, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n554, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n554, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n554, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n554, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n554, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n22999, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n554, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n554, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n554, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n554, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n22999, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n554, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n554, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n22999, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n554, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n554, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n7822, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n7822, Q => 
                           n9045);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n7822, Q => 
                           n9048);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n7822, Q => 
                           n9051);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n7822, Q => 
                           n9054);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n7822, Q => 
                           n9057);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n7822, Q => 
                           n9060);
   data1_mul_reg_8_inst : DLL_X1 port map( D => n19446, GN => n7822, Q => n9063
                           );
   data1_mul_reg_7_inst : DLL_X1 port map( D => n19444, GN => n7822, Q => n9066
                           );
   data1_mul_reg_6_inst : DLL_X1 port map( D => n19298, GN => n7822, Q => n9069
                           );
   data1_mul_reg_5_inst : DLL_X1 port map( D => n19299, GN => n7822, Q => n9072
                           );
   data1_mul_reg_4_inst : DLL_X1 port map( D => n19300, GN => n7822, Q => n9075
                           );
   data1_mul_reg_3_inst : DLL_X1 port map( D => n19443, GN => n7822, Q => n9078
                           );
   data1_mul_reg_2_inst : DLL_X1 port map( D => n19442, GN => n7822, Q => n9081
                           );
   data1_mul_reg_1_inst : DLL_X1 port map( D => n19302, GN => n7822, Q => n9084
                           );
   data1_mul_reg_0_inst : DLL_X1 port map( D => n19303, GN => n7822, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n7822, Q => 
                           n18199);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n7822, Q => 
                           n14292);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n7822, Q => 
                           n14290);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n7822, Q => 
                           n14288);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n7822, Q => 
                           n14287);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n7822, Q => 
                           n14286);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n7822, Q => 
                           n4302);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n7822, Q => 
                           n8978);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n7822, Q => 
                           n7769);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n7822, Q => 
                           n4295);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n7822, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n7822, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n554, Q => n4293);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1795, B => n1796, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1794, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1793, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1792, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1790, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1789, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1788, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1787, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1786, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1785, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1784, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1783, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1782, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1781, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1780, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3036,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => n14123);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => n14122);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => n14121);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => n14120);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => n14119);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => n14118);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => n14117);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => n14116);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => n14115);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => n14114);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => n14113);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => n14112);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => n14111);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => n14110);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1004, S => n14109);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => n19134, 
                           CI => n3026, CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => n14103);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => n19133, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => n19132, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => n19131, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => n19130, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => n19129,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => n19128,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => n19127,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => n19126,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => n19125,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => n19124,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => n19123,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => n19122,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => n19121,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => n14102);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => n19121,
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => n14101, S => n14100);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n18847, B => n19120, CI => n19114, CO => n_1005, S 
                           => boothmul_pipelined_i_sum_B_in_3_22_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3030,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => n14095);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => n4018);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => n4017);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => n4016);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => n4015);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => n4014);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => n4013);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => n4012);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => n8764);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => n14094, S => n14093);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n14145, B => n14102, CI => n14094, CO => n4009, S =>
                           n4008);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n19163, B => n19113, CI => n19106, CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n19162, B => boothmul_pipelined_i_sum_B_in_3_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n19161, B => boothmul_pipelined_i_sum_B_in_3_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n18846, B => boothmul_pipelined_i_sum_B_in_3_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1006, S => n4007);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => n4018, 
                           CI => n3029, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => n14088);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => n4017, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => n4016, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => n8755);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => n4015, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => n8754);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => n4014, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => n8753);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => n4013, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => n8752);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => n4012, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => n8751, S => n14087);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n8928, B => n8764, CI => n8751, CO => n14086, S => 
                           n14085);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n18899, B => n19107, CI => n19098, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => n3995);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n18898, B => n19105, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => n3994);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n18897, B => boothmul_pipelined_i_sum_B_in_4_19_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => n3993);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n18896, B => boothmul_pipelined_i_sum_B_in_4_20_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => n3992);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n18895, B => boothmul_pipelined_i_sum_B_in_4_21_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => n3991, S => n3990);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n18894, B => n4007, CI => n3991, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n18893, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => n8749);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n18852, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1007, S => n8748);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => n8755, 
                           CI => n3028, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => n14080);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => n8754, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => n8753, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => n14078);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => n8752, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => n14077, S => n14076);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           n19158, B => n19099, CI => n19090, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => n8740);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n19157, B => n19097, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => n8739);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n19156, B => n3995, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => n8738);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n19155, B => n3994, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => n8737);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n19154, B => n3993, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => n8736);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n19153, B => n3992, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => n8735);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n19152, B => n3990, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => n8734);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n19151, B => boothmul_pipelined_i_sum_B_in_5_22_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => n8733, S => n8732);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n19150, B => n8749, CI => n8733, CO => n3974, S => 
                           n3973);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n19149, B => n8748, CI => n3974, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n19148, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => n14075);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n18845, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1008, S => n14074);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           n18851, B => n19091, CI => n19193, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => n14070);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           n19247, B => n19089, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           n19246, B => n8740, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => n14068);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n19245, B => n8739, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => n14067);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n19244, B => n8738, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => n14066);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n19243, B => n8737, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => n14065);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n19242, B => n8736, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => n14064);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n19241, B => n8735, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => n14063);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n19240, B => n8734, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => n14062);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n19239, B => n8732, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => n14061);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n19238, B => n3973, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => n14060);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n19237, B => boothmul_pipelined_i_sum_B_in_6_24_port
                           , CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => n14059, S => n14058);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n19236, B => n14075, CI => n14059, CO => n3958, S =>
                           n3957);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n19235, B => n14074, CI => n3958, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n18892, B => n14074, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => n14057);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n18850, B => n14074, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1009, S => n14056);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => n14068,
                           CI => n3020, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => n14053);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => n14067,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => n14050);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => n14066,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => n14047);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => n14065,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => n14044);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => n14064,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => n14041);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => n14063,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => n14038);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => n14062,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => n14035);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => n14061,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => n14032);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => n14060,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => n14029);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => n14058,
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => n14026);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => n3957, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => n14023);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => n14022, S => n14019);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n19234, B => n19084, CI => n19037, CO => n3940, S =>
                           n14017);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n19233, B => n19083, CI => n3940, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => n14015);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           n19232, B => n19083, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => n14013);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           n19231, B => n19083, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => n14011);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           n19231, B => n19083, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1010, S => n14009);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n7822, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n554, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n554, Q => n4395);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n554, Q => 
                           DATA2_I_28_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port);
   clk_r_REG10887_S3 : DFFR_X1 port map( D => DATA1(8), CK => clk, RN => 
                           rst_BAR, Q => n19446, QN => n22969);
   clk_r_REG10319_S6 : DFFR_X1 port map( D => DATA1(7), CK => clk, RN => n21194
                           , Q => n19444, QN => n21165);
   clk_r_REG11582_S3 : DFFS_X1 port map( D => n1832, CK => clk, SN => n21195, Q
                           => n_1011, QN => n19443);
   clk_r_REG11724_S3 : DFFS_X1 port map( D => n1833, CK => clk, SN => n21202, Q
                           => n_1012, QN => n19442);
   clk_r_REG13375_S1 : DFFR_X1 port map( D => cin, CK => clk, RN => n21189, Q 
                           => n19441, QN => n22966);
   clk_r_REG13214_S5 : DFFS_X1 port map( D => n1796, CK => clk, SN => n21207, Q
                           => n19440, QN => n_1013);
   clk_r_REG11283_S5 : DFFS_X1 port map( D => n1791, CK => clk, SN => n21201, Q
                           => n19439, QN => n_1014);
   clk_r_REG11121_S16 : DFFS_X1 port map( D => n1780, CK => clk, SN => n21206, 
                           Q => n_1015, QN => n21181);
   clk_r_REG11223_S4 : DFFS_X1 port map( D => n18195, CK => clk, SN => n21207, 
                           Q => n_1016, QN => n19437);
   clk_r_REG13369_S3 : DFFR_X1 port map( D => n1815, CK => clk, RN => n21189, Q
                           => n19436, QN => n_1017);
   clk_r_REG10494_S5 : DFFR_X1 port map( D => n1779, CK => clk, RN => n21189, Q
                           => n19435, QN => n_1018);
   clk_r_REG10539_S11 : DFFR_X1 port map( D => n1811, CK => clk, RN => n21209, 
                           Q => n19434, QN => n_1019);
   clk_r_REG10587_S11 : DFFR_X1 port map( D => n1812, CK => clk, RN => n21190, 
                           Q => n19433, QN => n_1020);
   clk_r_REG12704_S4 : DFFS_X1 port map( D => n1825, CK => clk, SN => n21208, Q
                           => n19432, QN => n_1021);
   clk_r_REG12002_S4 : DFFS_X1 port map( D => n22998, CK => clk, SN => n21203, 
                           Q => n19431, QN => n_1022);
   clk_r_REG11867_S3 : DFFR_X1 port map( D => DATA1(1), CK => clk, RN => n21189
                           , Q => n_1023, QN => n19430);
   clk_r_REG13212_S3 : DFFR_X1 port map( D => DATA1(0), CK => clk, RN => 
                           rst_BAR, Q => n_1024, QN => n19429);
   clk_r_REG11278_S3 : DFFR_X1 port map( D => DATA1(4), CK => clk, RN => 
                           rst_BAR, Q => n_1025, QN => n19428);
   clk_r_REG11363_S6 : DFFR_X1 port map( D => DATA1(6), CK => clk, RN => n21189
                           , Q => n_1026, QN => n19427);
   clk_r_REG11358_S6 : DFFR_X1 port map( D => DATA1(5), CK => clk, RN => 
                           rst_BAR, Q => n22986, QN => n19426);
   clk_r_REG11239_S4 : DFFR_X1 port map( D => n22997, CK => clk, RN => n21195, 
                           Q => n19425, QN => n_1027);
   clk_r_REG10997_S15 : DFFR_X1 port map( D => n1822, CK => clk, RN => n21198, 
                           Q => n22977, QN => n21169);
   clk_r_REG11235_S4 : DFFS_X1 port map( D => n13151, CK => clk, SN => n21205, 
                           Q => n_1028, QN => n19423);
   clk_r_REG11228_S4 : DFFS_X1 port map( D => n1896, CK => clk, SN => n21196, Q
                           => n_1029, QN => n19422);
   clk_r_REG11232_S4 : DFFS_X1 port map( D => n1894, CK => clk, SN => n21195, Q
                           => n_1030, QN => n19421);
   clk_r_REG11212_S4 : DFFS_X1 port map( D => n17728, CK => clk, SN => n21207, 
                           Q => n_1031, QN => n19420);
   clk_r_REG10982_S15 : DFFS_X1 port map( D => n1820, CK => clk, SN => n21198, 
                           Q => n19419, QN => n_1032);
   clk_r_REG10507_S4 : DFFS_X1 port map( D => n1829, CK => clk, SN => n21211, Q
                           => n19418, QN => n_1033);
   clk_r_REG10498_S4 : DFFR_X1 port map( D => n1827, CK => clk, RN => n21209, Q
                           => n19417, QN => n_1034);
   clk_r_REG10497_S4 : DFFR_X1 port map( D => n1818, CK => clk, RN => n21210, Q
                           => n19416, QN => n_1035);
   clk_r_REG10757_S4 : DFFS_X1 port map( D => n1804, CK => clk, SN => n21203, Q
                           => n19414, QN => n_1036);
   clk_r_REG11209_S4 : DFFS_X1 port map( D => n21157, CK => clk, SN => n21204, 
                           Q => n19412, QN => n_1037);
   clk_r_REG11442_S5 : DFFS_X1 port map( D => n1799, CK => clk, SN => n21198, Q
                           => n19411, QN => n_1038);
   clk_r_REG11206_S4 : DFFS_X1 port map( D => n21171, CK => clk, SN => n21197, 
                           Q => n19409, QN => n22982);
   clk_r_REG11240_S4 : DFFS_X1 port map( D => n22997, CK => clk, SN => n21200, 
                           Q => n19408, QN => n_1039);
   clk_r_REG11186_S4 : DFFS_X1 port map( D => n21172, CK => clk, SN => n21204, 
                           Q => n19407, QN => n_1040);
   clk_r_REG10863_S4 : DFFR_X1 port map( D => n1808, CK => clk, RN => n21196, Q
                           => n19406, QN => n_1041);
   clk_r_REG11166_S4 : DFFR_X1 port map( D => n21174, CK => clk, RN => n21207, 
                           Q => n19405, QN => n22974);
   clk_r_REG11185_S4 : DFFR_X1 port map( D => n21172, CK => clk, RN => n21209, 
                           Q => n19404, QN => n22978);
   clk_r_REG10518_S4 : DFFR_X1 port map( D => n1819, CK => clk, RN => n21212, Q
                           => n19403, QN => n_1042);
   clk_r_REG10679_S4 : DFFS_X1 port map( D => n1805, CK => clk, SN => n21203, Q
                           => n19402, QN => n_1043);
   clk_r_REG10413_S4 : DFFR_X1 port map( D => n1816, CK => clk, RN => n21202, Q
                           => n19401, QN => n_1044);
   clk_r_REG11013_S4 : DFFS_X1 port map( D => n1821, CK => clk, SN => n21202, Q
                           => n19400, QN => n_1045);
   clk_r_REG12195_S4 : DFFR_X1 port map( D => n1817, CK => clk, RN => n21193, Q
                           => n19399, QN => n_1046);
   clk_r_REG10995_S15 : DFFS_X1 port map( D => n1824, CK => clk, SN => n21202, 
                           Q => n19398, QN => n_1047);
   clk_r_REG11192_S4 : DFFR_X1 port map( D => n1838, CK => clk, RN => n21196, Q
                           => n19397, QN => n22989);
   clk_r_REG11201_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => n21200, Q
                           => n19396, QN => n_1048);
   clk_r_REG11247_S4 : DFFR_X1 port map( D => n1847, CK => clk, RN => n21198, Q
                           => n19395, QN => n_1049);
   clk_r_REG11273_S4 : DFFS_X1 port map( D => n1846, CK => clk, SN => n21207, Q
                           => n19394, QN => n22985);
   clk_r_REG11179_S4 : DFFR_X1 port map( D => n21160, CK => clk, RN => n21195, 
                           Q => n19393, QN => n_1050);
   clk_r_REG11180_S4 : DFFS_X1 port map( D => n21160, CK => clk, SN => n21196, 
                           Q => n19392, QN => n22972);
   clk_r_REG11176_S4 : DFFS_X1 port map( D => n21170, CK => clk, SN => n21195, 
                           Q => n19391, QN => n_1051);
   clk_r_REG11253_S4 : DFFS_X1 port map( D => n21178, CK => clk, SN => n21203, 
                           Q => n19390, QN => n_1052);
   clk_r_REG11275_S4 : DFFS_X1 port map( D => n21180, CK => clk, SN => n21206, 
                           Q => n19389, QN => n_1053);
   clk_r_REG10515_S4 : DFFS_X1 port map( D => n1823, CK => clk, SN => n21201, Q
                           => n19388, QN => n_1054);
   clk_r_REG10884_S5 : DFFS_X1 port map( D => n1798, CK => clk, SN => n21200, Q
                           => n19387, QN => n_1055);
   clk_r_REG11236_S4 : DFFS_X1 port map( D => n13151, CK => clk, SN => n21208, 
                           Q => n19386, QN => n_1056);
   clk_r_REG11222_S4 : DFFS_X1 port map( D => n1841, CK => clk, SN => n21195, Q
                           => n19385, QN => n22979);
   clk_r_REG12640_S5 : DFFS_X1 port map( D => n1800, CK => clk, SN => n21200, Q
                           => n19384, QN => n_1057);
   clk_r_REG10672_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_102_port, CK => clk,
                           RN => n21195, Q => n19383, QN => n_1058);
   clk_r_REG10668_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_103_port, CK => clk,
                           RN => n21207, Q => n19382, QN => n_1059);
   clk_r_REG10749_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_104_port, CK => clk,
                           RN => n21189, Q => n19381, QN => n_1060);
   clk_r_REG10748_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_105_port, CK => clk,
                           RN => n21200, Q => n19380, QN => n_1061);
   clk_r_REG10745_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_106_port, CK => clk,
                           RN => n21212, Q => n19379, QN => n_1062);
   clk_r_REG10785_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_107_port, CK => clk,
                           RN => n21189, Q => n19378, QN => n_1063);
   clk_r_REG10852_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_108_port, CK => clk,
                           RN => n21204, Q => n19377, QN => n_1064);
   clk_r_REG10889_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_109_port, CK => clk,
                           RN => n21203, Q => n19376, QN => n_1065);
   clk_r_REG11287_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_110_port, CK => clk,
                           RN => n21209, Q => n19375, QN => n_1066);
   clk_r_REG11286_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_111_port, CK => clk,
                           RN => n21205, Q => n19374, QN => n_1067);
   clk_r_REG11285_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_112_port, CK => clk,
                           RN => n21190, Q => n19373, QN => n_1068);
   clk_r_REG11284_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_113_port, CK => clk,
                           RN => n21204, Q => n19372, QN => n_1069);
   clk_r_REG11584_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_114_port, CK => clk,
                           RN => n21205, Q => n19371, QN => n_1070);
   clk_r_REG11726_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_115_port, CK => clk,
                           RN => n21204, Q => n19370, QN => n_1071);
   clk_r_REG11871_S5 : DFFR_X1 port map( D => n21214, CK => clk, RN => n21189, 
                           Q => n19369, QN => n_1072);
   clk_r_REG11193_S4 : DFFR_X1 port map( D => n1840, CK => clk, RN => n21203, Q
                           => n19368, QN => n_1073);
   clk_r_REG11194_S4 : DFFS_X1 port map( D => n1840, CK => clk, SN => n21200, Q
                           => n19367, QN => n_1074);
   clk_r_REG11255_S4 : DFFS_X1 port map( D => n21177, CK => clk, SN => n21194, 
                           Q => n19366, QN => n22993);
   clk_r_REG10798_S5 : DFFS_X1 port map( D => n21183, CK => clk, SN => n21207, 
                           Q => n19365, QN => n_1075);
   clk_r_REG11196_S4 : DFFS_X1 port map( D => n21179, CK => clk, SN => n21200, 
                           Q => n19364, QN => n22973);
   clk_r_REG11213_S4 : DFFS_X1 port map( D => n17728, CK => clk, SN => n21201, 
                           Q => n19363, QN => n_1076);
   clk_r_REG11257_S4 : DFFS_X1 port map( D => n21175, CK => clk, SN => n21198, 
                           Q => n19362, QN => n_1077);
   clk_r_REG11250_S4 : DFFR_X1 port map( D => n1845, CK => clk, RN => n21190, Q
                           => n19361, QN => n22990);
   clk_r_REG11249_S4 : DFFS_X1 port map( D => n1845, CK => clk, SN => n21200, Q
                           => n19360, QN => n22994);
   clk_r_REG11259_S4 : DFFR_X1 port map( D => n21176, CK => clk, RN => n21191, 
                           Q => n19359, QN => n_1078);
   clk_r_REG10422_S5 : DFFS_X1 port map( D => n21186, CK => clk, SN => n21200, 
                           Q => n19358, QN => n_1079);
   clk_r_REG10847_S5 : DFFS_X1 port map( D => n21163, CK => clk, SN => n21204, 
                           Q => n19357, QN => n_1080);
   clk_r_REG11234_S4 : DFFS_X1 port map( D => n1837, CK => clk, SN => n21196, Q
                           => n19356, QN => n_1081);
   clk_r_REG11267_S4 : DFFS_X1 port map( D => n1813, CK => clk, SN => n21195, Q
                           => n19355, QN => n_1082);
   clk_r_REG11263_S4 : DFFS_X1 port map( D => n1814, CK => clk, SN => n21206, Q
                           => n19354, QN => n_1083);
   clk_r_REG13370_S3 : DFFS_X1 port map( D => n17537, CK => clk, SN => n21197, 
                           Q => n19353, QN => n_1084);
   clk_r_REG10673_S5 : DFFR_X1 port map( D => n18051, CK => clk, RN => n21207, 
                           Q => n19352, QN => n_1085);
   clk_r_REG10728_S5 : DFFS_X1 port map( D => n1797, CK => clk, SN => n21205, Q
                           => n_1086, QN => n21161);
   clk_r_REG10547_S6 : DFFS_X1 port map( D => n21158, CK => clk, SN => n21206, 
                           Q => n_1087, QN => n21159);
   clk_r_REG11872_S5 : DFFR_X1 port map( D => n9084, CK => clk, RN => n21199, Q
                           => n19349, QN => n_1088);
   clk_r_REG11727_S5 : DFFR_X1 port map( D => n9081, CK => clk, RN => n21199, Q
                           => n19348, QN => n_1089);
   clk_r_REG11585_S5 : DFFR_X1 port map( D => n9078, CK => clk, RN => n21190, Q
                           => n19347, QN => n_1090);
   clk_r_REG11288_S5 : DFFR_X1 port map( D => n9075, CK => clk, RN => n21194, Q
                           => n19346, QN => n_1091);
   clk_r_REG11360_S8 : DFFR_X1 port map( D => n9072, CK => clk, RN => n21206, Q
                           => n19345, QN => n_1092);
   clk_r_REG11366_S8 : DFFR_X1 port map( D => n9069, CK => clk, RN => n21212, Q
                           => n19344, QN => n_1093);
   clk_r_REG13282_S8 : DFFR_X1 port map( D => n9066, CK => clk, RN => n21209, Q
                           => n19343, QN => n_1094);
   clk_r_REG10890_S5 : DFFR_X1 port map( D => n9063, CK => clk, RN => n21200, Q
                           => n19342, QN => n_1095);
   clk_r_REG10853_S5 : DFFR_X1 port map( D => n9060, CK => clk, RN => n21192, Q
                           => n19341, QN => n_1096);
   clk_r_REG10786_S5 : DFFR_X1 port map( D => n9057, CK => clk, RN => n21211, Q
                           => n19340, QN => n_1097);
   clk_r_REG10750_S5 : DFFR_X1 port map( D => n9054, CK => clk, RN => n21210, Q
                           => n19339, QN => n_1098);
   clk_r_REG11139_S15 : DFFR_X1 port map( D => n9051, CK => clk, RN => n21196, 
                           Q => n19338, QN => n_1099);
   clk_r_REG11128_S15 : DFFR_X1 port map( D => n9048, CK => clk, RN => n21191, 
                           Q => n19337, QN => n_1100);
   clk_r_REG10674_S5 : DFFR_X1 port map( D => n9045, CK => clk, RN => n21194, Q
                           => n19336, QN => n_1101);
   clk_r_REG11868_S3 : DFFR_X1 port map( D => DATA1(1), CK => clk, RN => n21192
                           , Q => n19335, QN => n_1102);
   clk_r_REG11224_S4 : DFFS_X1 port map( D => n18195, CK => clk, SN => n21196, 
                           Q => n19334, QN => n_1103);
   clk_r_REG11202_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => n21205, Q
                           => n19333, QN => n22981);
   clk_r_REG11175_S4 : DFFS_X1 port map( D => n21170, CK => clk, SN => n21200, 
                           Q => n19332, QN => n_1104);
   clk_r_REG11181_S4 : DFFS_X1 port map( D => n21160, CK => clk, SN => n21206, 
                           Q => n19331, QN => n_1105);
   clk_r_REG11210_S4 : DFFS_X1 port map( D => n21157, CK => clk, SN => n21195, 
                           Q => n19330, QN => n_1106);
   clk_r_REG11203_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => n21204, Q
                           => n19329, QN => n_1107);
   clk_r_REG11272_S4 : DFFR_X1 port map( D => n1846, CK => clk, RN => n21212, Q
                           => n19328, QN => n22995);
   clk_r_REG11271_S4 : DFFS_X1 port map( D => n1846, CK => clk, SN => n21199, Q
                           => n19327, QN => n_1108);
   clk_r_REG11268_S4 : DFFS_X1 port map( D => n1813, CK => clk, SN => n21203, Q
                           => n19326, QN => n_1109);
   clk_r_REG11204_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => n21206, Q
                           => n19325, QN => n_1110);
   clk_r_REG11197_S4 : DFFS_X1 port map( D => n21179, CK => clk, SN => n21201, 
                           Q => n19324, QN => n_1111);
   clk_r_REG11252_S4 : DFFS_X1 port map( D => n21178, CK => clk, SN => n21198, 
                           Q => n19323, QN => n_1112);
   clk_r_REG11174_S4 : DFFR_X1 port map( D => n21170, CK => clk, RN => n21210, 
                           Q => n19322, QN => n_1113);
   clk_r_REG11246_S4 : DFFR_X1 port map( D => n1847, CK => clk, RN => n21193, Q
                           => n19321, QN => n22992);
   clk_r_REG11191_S4 : DFFR_X1 port map( D => n1838, CK => clk, RN => n21191, Q
                           => n19320, QN => n_1114);
   clk_r_REG11184_S4 : DFFS_X1 port map( D => n21172, CK => clk, SN => n21204, 
                           Q => n19319, QN => n_1115);
   clk_r_REG10500_S4 : DFFS_X1 port map( D => n1826, CK => clk, SN => n21199, Q
                           => n19318, QN => n_1116);
   clk_r_REG11167_S4 : DFFR_X1 port map( D => n21174, CK => clk, RN => n21199, 
                           Q => n19317, QN => n_1117);
   clk_r_REG11264_S4 : DFFS_X1 port map( D => n1814, CK => clk, SN => n21190, Q
                           => n19316, QN => n_1118);
   clk_r_REG11208_S4 : DFFS_X1 port map( D => n21157, CK => clk, SN => n21199, 
                           Q => n19315, QN => n_1119);
   clk_r_REG11233_S4 : DFFS_X1 port map( D => n1894, CK => clk, SN => n21208, Q
                           => n19314, QN => n_1120);
   clk_r_REG11237_S4 : DFFR_X1 port map( D => n1836, CK => clk, RN => n21194, Q
                           => n19313, QN => n_1121);
   clk_r_REG11364_S6 : DFFR_X1 port map( D => DATA1(6), CK => clk, RN => n21190
                           , Q => n19312, QN => n_1122);
   clk_r_REG11583_S3 : DFFS_X1 port map( D => n1832, CK => clk, SN => n21206, Q
                           => n19311, QN => n_1123);
   clk_r_REG10384_S5 : DFFR_X1 port map( D => n1801, CK => clk, RN => n21211, Q
                           => n19310, QN => n_1124);
   clk_r_REG11725_S3 : DFFS_X1 port map( D => n1833, CK => clk, SN => n21206, Q
                           => n19309, QN => n_1125);
   clk_r_REG11229_S4 : DFFS_X1 port map( D => n1896, CK => clk, SN => n21206, Q
                           => n19308, QN => n_1126);
   clk_r_REG11226_S4 : DFFS_X1 port map( D => n18195, CK => clk, SN => n21204, 
                           Q => n19307, QN => n_1127);
   clk_r_REG11243_S4 : DFFR_X1 port map( D => n1834, CK => clk, RN => n21191, Q
                           => n19306, QN => n_1128);
   clk_r_REG11244_S4 : DFFS_X1 port map( D => n1834, CK => clk, SN => n21205, Q
                           => n19305, QN => n_1129);
   clk_r_REG11242_S4 : DFFS_X1 port map( D => n1839, CK => clk, SN => n21198, Q
                           => n19304, QN => n22991);
   clk_r_REG13213_S3 : DFFR_X1 port map( D => DATA1(0), CK => clk, RN => 
                           rst_BAR, Q => n19303, QN => n22987);
   clk_r_REG11869_S3 : DFFR_X1 port map( D => DATA1(1), CK => clk, RN => n21192
                           , Q => n19302, QN => n_1130);
   clk_r_REG11870_S4 : DFFS_X1 port map( D => n19302, CK => clk, SN => n21205, 
                           Q => n19301, QN => n_1131);
   clk_r_REG11279_S3 : DFFR_X1 port map( D => DATA1(4), CK => clk, RN => n21189
                           , Q => n19300, QN => n_1132);
   clk_r_REG11359_S6 : DFFR_X1 port map( D => DATA1(5), CK => clk, RN => n21189
                           , Q => n19299, QN => n_1133);
   clk_r_REG11365_S6 : DFFR_X1 port map( D => DATA1(6), CK => clk, RN => n21194
                           , Q => n19298, QN => n22970);
   clk_r_REG10624_S5 : DFFR_X1 port map( D => n18199, CK => clk, RN => n21212, 
                           Q => n19297, QN => n_1134);
   clk_r_REG10625_S6 : DFFR_X1 port map( D => n19297, CK => clk, RN => n21194, 
                           Q => n22975, QN => n21166);
   clk_r_REG10640_S5 : DFFR_X1 port map( D => n14292, CK => clk, RN => n21210, 
                           Q => n19295, QN => n_1135);
   clk_r_REG10641_S6 : DFFR_X1 port map( D => n19295, CK => clk, RN => n21201, 
                           Q => n19294, QN => n_1136);
   clk_r_REG10546_S5 : DFFR_X1 port map( D => n14290, CK => clk, RN => n21212, 
                           Q => n19293, QN => n21158);
   clk_r_REG10527_S5 : DFFR_X1 port map( D => n14288, CK => clk, RN => n21205, 
                           Q => n19292, QN => n_1137);
   clk_r_REG11157_S5 : DFFR_X1 port map( D => n21188, CK => clk, RN => n21202, 
                           Q => n_1138, QN => n19290);
   clk_r_REG11199_S4 : DFFR_X1 port map( D => n1834, CK => clk, RN => n21193, Q
                           => n_1139, QN => n19289);
   clk_r_REG11198_S4 : DFFS_X1 port map( D => n1834, CK => clk, SN => n21194, Q
                           => n_1140, QN => n19288);
   clk_r_REG11241_S4 : DFFS_X1 port map( D => n1839, CK => clk, SN => n21197, Q
                           => n22962, QN => n19287);
   clk_r_REG11270_S4 : DFFR_X1 port map( D => n1846, CK => clk, RN => n21204, Q
                           => n_1141, QN => n19286);
   clk_r_REG11269_S4 : DFFS_X1 port map( D => n1846, CK => clk, SN => n21206, Q
                           => n_1142, QN => n19285);
   clk_r_REG11101_S5 : DFFS_X1 port map( D => n1809, CK => clk, SN => n21195, Q
                           => n19284, QN => n_1143);
   clk_r_REG10468_S5 : DFFS_X1 port map( D => n13929, CK => clk, SN => n21203, 
                           Q => n19283, QN => n_1144);
   clk_r_REG11265_S4 : DFFS_X1 port map( D => n1813, CK => clk, SN => n21208, Q
                           => n22983, QN => n19282);
   clk_r_REG11262_S4 : DFFS_X1 port map( D => n1814, CK => clk, SN => n21197, Q
                           => n_1145, QN => n19281);
   clk_r_REG11440_S5 : DFFS_X1 port map( D => n1799, CK => clk, SN => n21204, Q
                           => n_1146, QN => n19279);
   clk_r_REG11441_S5 : DFFS_X1 port map( D => n14281, CK => clk, SN => n21208, 
                           Q => n19278, QN => n_1147);
   clk_r_REG10630_S5 : DFFR_X1 port map( D => n14278, CK => clk, RN => n21194, 
                           Q => n19277, QN => n_1148);
   clk_r_REG10871_S6 : DFFR_X1 port map( D => n14176, CK => clk, RN => n21211, 
                           Q => n19276, QN => n_1149);
   clk_r_REG10872_S7 : DFFR_X1 port map( D => n19276, CK => clk, RN => n21190, 
                           Q => n19275, QN => n_1150);
   clk_r_REG10873_S8 : DFFR_X1 port map( D => n19275, CK => clk, RN => n21211, 
                           Q => n19274, QN => n_1151);
   clk_r_REG10874_S9 : DFFR_X1 port map( D => n19274, CK => clk, RN => n21210, 
                           Q => n19273, QN => n_1152);
   clk_r_REG10875_S10 : DFFR_X1 port map( D => n19273, CK => clk, RN => n21189,
                           Q => n19272, QN => n_1153);
   clk_r_REG11266_S4 : DFFS_X1 port map( D => n14273, CK => clk, SN => n21208, 
                           Q => n19271, QN => n_1154);
   clk_r_REG11170_S5 : DFFS_X1 port map( D => n14272, CK => clk, SN => n21199, 
                           Q => n19270, QN => n_1155);
   clk_r_REG11580_S5 : DFFS_X1 port map( D => n14271, CK => clk, SN => n21194, 
                           Q => n19269, QN => n_1156);
   clk_r_REG10383_S5 : DFFS_X1 port map( D => n17140, CK => clk, SN => n21196, 
                           Q => n19268, QN => n_1157);
   clk_r_REG11050_S4 : DFFS_X1 port map( D => n14268, CK => clk, SN => n21204, 
                           Q => n19267, QN => n_1158);
   clk_r_REG11042_S5 : DFFS_X1 port map( D => n14266, CK => clk, SN => n21202, 
                           Q => n19266, QN => n_1159);
   clk_r_REG10433_S11 : DFFS_X1 port map( D => n14265, CK => clk, SN => n21199,
                           Q => n19265, QN => n_1160);
   clk_r_REG10598_S11 : DFFR_X1 port map( D => n17388, CK => clk, RN => n21196,
                           Q => n19264, QN => n_1161);
   clk_r_REG10736_S5 : DFFS_X1 port map( D => n17503, CK => clk, SN => n21199, 
                           Q => n19263, QN => n_1162);
   clk_r_REG11225_S4 : DFFS_X1 port map( D => n17471, CK => clk, SN => n21208, 
                           Q => n19262, QN => n_1163);
   clk_r_REG11190_S4 : DFFR_X1 port map( D => n17506, CK => clk, RN => n21197, 
                           Q => n19261, QN => n_1164);
   clk_r_REG11260_S4 : DFFS_X1 port map( D => n8626, CK => clk, SN => n21208, Q
                           => n19260, QN => n_1165);
   clk_r_REG11261_S4 : DFFS_X1 port map( D => n14259, CK => clk, SN => n21199, 
                           Q => n19259, QN => n_1166);
   clk_r_REG10327_S5 : DFFR_X1 port map( D => n14253, CK => clk, RN => n21191, 
                           Q => n19258, QN => n_1167);
   clk_r_REG10328_S6 : DFFR_X1 port map( D => n19258, CK => clk, RN => n21191, 
                           Q => n19257, QN => n_1168);
   clk_r_REG10329_S7 : DFFR_X1 port map( D => n19257, CK => clk, RN => n21212, 
                           Q => n19256, QN => n_1169);
   clk_r_REG10330_S8 : DFFR_X1 port map( D => n19256, CK => clk, RN => n21195, 
                           Q => n19255, QN => n_1170);
   clk_r_REG10331_S9 : DFFR_X1 port map( D => n19255, CK => clk, RN => n21199, 
                           Q => n19254, QN => n_1171);
   clk_r_REG10332_S10 : DFFR_X1 port map( D => n19254, CK => clk, RN => n21192,
                           Q => n19253, QN => n_1172);
   clk_r_REG10811_S5 : DFFS_X1 port map( D => n14252, CK => clk, SN => n21207, 
                           Q => n19252, QN => n_1173);
   clk_r_REG10729_S5 : DFFS_X1 port map( D => n21185, CK => clk, SN => n21206, 
                           Q => n_1174, QN => n19249);
   clk_r_REG10727_S5 : DFFS_X1 port map( D => n17966, CK => clk, SN => n21199, 
                           Q => n19248, QN => n_1175);
   clk_r_REG10732_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_14_port, CK => clk, 
                           RN => n21196, Q => n19247, QN => n_1176);
   clk_r_REG10612_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_15_port, CK => clk, 
                           RN => n21204, Q => n19246, QN => n_1177);
   clk_r_REG10611_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_16_port, CK => clk, 
                           RN => n21208, Q => n19245, QN => n_1178);
   clk_r_REG10605_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_17_port, CK => clk, 
                           RN => n21212, Q => n19244, QN => n_1179);
   clk_r_REG10599_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_18_port, CK => clk, 
                           RN => n21207, Q => n19243, QN => n_1180);
   clk_r_REG10593_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_19_port, CK => clk, 
                           RN => n21203, Q => n19242, QN => n_1181);
   clk_r_REG10588_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_20_port, CK => clk, 
                           RN => n21197, Q => n19241, QN => n_1182);
   clk_r_REG10582_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_21_port, CK => clk, 
                           RN => n21192, Q => n19240, QN => n_1183);
   clk_r_REG10581_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_22_port, CK => clk, 
                           RN => n21189, Q => n19239, QN => n_1184);
   clk_r_REG10580_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_23_port, CK => clk, 
                           RN => n21203, Q => n19238, QN => n_1185);
   clk_r_REG10579_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_24_port, CK => clk, 
                           RN => n21211, Q => n19237, QN => n_1186);
   clk_r_REG10574_S6 : DFFR_X1 port map( D => n14239, CK => clk, RN => n21211, 
                           Q => n19236, QN => n_1187);
   clk_r_REG10568_S6 : DFFR_X1 port map( D => n14238, CK => clk, RN => n21192, 
                           Q => n19235, QN => n_1188);
   clk_r_REG10629_S7 : DFFR_X1 port map( D => n14237, CK => clk, RN => n21189, 
                           Q => n19234, QN => n_1189);
   clk_r_REG10628_S7 : DFFR_X1 port map( D => n14236, CK => clk, RN => n21204, 
                           Q => n19233, QN => n_1190);
   clk_r_REG10627_S7 : DFFR_X1 port map( D => n14235, CK => clk, RN => n21195, 
                           Q => n19232, QN => n_1191);
   clk_r_REG10626_S7 : DFFR_X1 port map( D => n14234, CK => clk, RN => n21190, 
                           Q => n19231, QN => n_1192);
   clk_r_REG11188_S4 : DFFR_X1 port map( D => n1840, CK => clk, RN => n21203, Q
                           => n22971, QN => n19230);
   clk_r_REG11187_S4 : DFFS_X1 port map( D => n1840, CK => clk, SN => n21204, Q
                           => n_1193, QN => n19229);
   clk_r_REG11251_S4 : DFFS_X1 port map( D => n21178, CK => clk, SN => n21198, 
                           Q => n_1194, QN => n19228);
   clk_r_REG11178_S4 : DFFR_X1 port map( D => n21160, CK => clk, RN => n21202, 
                           Q => n_1195, QN => n19227);
   clk_r_REG11177_S4 : DFFS_X1 port map( D => n21160, CK => clk, SN => n21195, 
                           Q => n_1196, QN => n19226);
   clk_r_REG11173_S4 : DFFR_X1 port map( D => n21170, CK => clk, RN => n21211, 
                           Q => n22984, QN => n19225);
   clk_r_REG11172_S4 : DFFS_X1 port map( D => n21170, CK => clk, SN => n21198, 
                           Q => n_1197, QN => n19224);
   clk_r_REG11258_S4 : DFFR_X1 port map( D => n21176, CK => clk, RN => n21202, 
                           Q => n22967, QN => n19223);
   clk_r_REG11207_S4 : DFFS_X1 port map( D => n21157, CK => clk, SN => n21196, 
                           Q => n22963, QN => n19222);
   clk_r_REG11254_S4 : DFFS_X1 port map( D => n21177, CK => clk, SN => n21202, 
                           Q => n_1198, QN => n19221);
   clk_r_REG11256_S4 : DFFS_X1 port map( D => n21175, CK => clk, SN => n21198, 
                           Q => n22964, QN => n19220);
   clk_r_REG10844_S5 : DFFR_X1 port map( D => n21187, CK => clk, RN => n21208, 
                           Q => n_1199, QN => n19218);
   clk_r_REG11238_S4 : DFFS_X1 port map( D => n22997, CK => clk, SN => n21200, 
                           Q => n_1200, QN => n19216);
   clk_r_REG10883_S5 : DFFS_X1 port map( D => n1798, CK => clk, SN => n21206, Q
                           => n_1201, QN => n19214);
   clk_r_REG11156_S5 : DFFS_X1 port map( D => n14132, CK => clk, SN => n21204, 
                           Q => n19213, QN => n_1202);
   clk_r_REG11274_S4 : DFFS_X1 port map( D => n21180, CK => clk, SN => n21196, 
                           Q => n22965, QN => n19212);
   clk_r_REG11195_S4 : DFFS_X1 port map( D => n21179, CK => clk, SN => n21201, 
                           Q => n22960, QN => n19211);
   clk_r_REG11221_S4 : DFFS_X1 port map( D => n1841, CK => clk, SN => n21203, Q
                           => n_1203, QN => n19210);
   clk_r_REG11168_S5 : DFFS_X1 port map( D => n1429, CK => clk, SN => n21199, Q
                           => n19209, QN => n_1204);
   clk_r_REG10363_S5 : DFFS_X1 port map( D => n8847, CK => clk, SN => n21202, Q
                           => n19208, QN => n_1205);
   clk_r_REG10788_S4 : DFFS_X1 port map( D => n14146, CK => clk, SN => n21203, 
                           Q => n19207, QN => n_1206);
   clk_r_REG11230_S4 : DFFR_X1 port map( D => n1836, CK => clk, RN => n21201, Q
                           => n_1207, QN => n19206);
   clk_r_REG11227_S4 : DFFS_X1 port map( D => n1835, CK => clk, SN => n21207, Q
                           => n_1208, QN => n19205);
   clk_r_REG11231_S4 : DFFS_X1 port map( D => n1837, CK => clk, SN => n21204, Q
                           => n_1209, QN => n19204);
   clk_r_REG11211_S4 : DFFS_X1 port map( D => n1843, CK => clk, SN => n21197, Q
                           => n_1210, QN => n19203);
   clk_r_REG11032_S15 : DFFR_X1 port map( D => n14184, CK => clk, RN => n21212,
                           Q => n19202, QN => n_1211);
   clk_r_REG11155_S5 : DFFS_X1 port map( D => n2808, CK => clk, SN => n21199, Q
                           => n19201, QN => n_1212);
   clk_r_REG10781_S5 : DFFS_X1 port map( D => n17932, CK => clk, SN => n21203, 
                           Q => n19199, QN => n_1213);
   clk_r_REG10769_S6 : DFFR_X1 port map( D => n13873, CK => clk, RN => n21198, 
                           Q => n19198, QN => n_1214);
   clk_r_REG10770_S7 : DFFR_X1 port map( D => n19198, CK => clk, RN => n21204, 
                           Q => n19197, QN => n_1215);
   clk_r_REG10771_S8 : DFFR_X1 port map( D => n19197, CK => clk, RN => n21211, 
                           Q => n19196, QN => n_1216);
   clk_r_REG10772_S9 : DFFR_X1 port map( D => n19196, CK => clk, RN => n21197, 
                           Q => n19195, QN => n_1217);
   clk_r_REG10773_S10 : DFFR_X1 port map( D => n19195, CK => clk, RN => n21201,
                           Q => n19194, QN => n_1218);
   clk_r_REG10534_S6 : DFFR_X1 port map( D => n3027, CK => clk, RN => n21193, Q
                           => n19193, QN => n_1219);
   clk_r_REG11716_S5 : DFFR_X1 port map( D => n14170, CK => clk, RN => n21190, 
                           Q => n19192, QN => n_1220);
   clk_r_REG11717_S6 : DFFR_X1 port map( D => n19192, CK => clk, RN => n21203, 
                           Q => n19191, QN => n_1221);
   clk_r_REG11718_S7 : DFFR_X1 port map( D => n19191, CK => clk, RN => n21190, 
                           Q => n19190, QN => n_1222);
   clk_r_REG11719_S8 : DFFR_X1 port map( D => n19190, CK => clk, RN => n21204, 
                           Q => n19189, QN => n_1223);
   clk_r_REG11720_S9 : DFFR_X1 port map( D => n19189, CK => clk, RN => n21195, 
                           Q => n19188, QN => n_1224);
   clk_r_REG11721_S10 : DFFR_X1 port map( D => n19188, CK => clk, RN => n21192,
                           Q => n19187, QN => n_1225);
   clk_r_REG10860_S4 : DFFS_X1 port map( D => n14168, CK => clk, SN => n21208, 
                           Q => n19186, QN => n_1226);
   clk_r_REG10837_S11 : DFFS_X1 port map( D => n16797, CK => clk, SN => n21202,
                           Q => n19185, QN => n_1227);
   clk_r_REG10823_S11 : DFFS_X1 port map( D => n13976, CK => clk, SN => n21205,
                           Q => n19184, QN => n_1228);
   clk_r_REG11033_S15 : DFFR_X1 port map( D => n13942, CK => clk, RN => n21211,
                           Q => n19183, QN => n_1229);
   clk_r_REG10382_S5 : DFFR_X1 port map( D => n14269, CK => clk, RN => n21210, 
                           Q => n19182, QN => n_1230);
   clk_r_REG10364_S5 : DFFR_X1 port map( D => n14164, CK => clk, RN => n21201, 
                           Q => n19181, QN => n_1231);
   clk_r_REG11214_S4 : DFFS_X1 port map( D => n14161, CK => clk, SN => n21200, 
                           Q => n19180, QN => n_1232);
   clk_r_REG10447_S5 : DFFS_X1 port map( D => n17254, CK => clk, SN => n21196, 
                           Q => n19179, QN => n_1233);
   clk_r_REG10446_S5 : DFFS_X1 port map( D => n14160, CK => clk, SN => n21195, 
                           Q => n19178, QN => n_1234);
   clk_r_REG10445_S4 : DFFR_X1 port map( D => n17270, CK => clk, RN => n21198, 
                           Q => n19177, QN => n_1235);
   clk_r_REG10409_S4 : DFFS_X1 port map( D => n14159, CK => clk, SN => n21201, 
                           Q => n19176, QN => n_1236);
   clk_r_REG10395_S5 : DFFR_X1 port map( D => n14158, CK => clk, RN => n21190, 
                           Q => n19175, QN => n_1237);
   clk_r_REG11030_S4 : DFFR_X1 port map( D => n14157, CK => clk, RN => n21210, 
                           Q => n19174, QN => n_1238);
   clk_r_REG10388_S4 : DFFS_X1 port map( D => n12313, CK => clk, SN => n21199, 
                           Q => n_1239, QN => n21182);
   clk_r_REG10486_S5 : DFFS_X1 port map( D => n14263, CK => clk, SN => n21199, 
                           Q => n19172, QN => n_1240);
   clk_r_REG11219_S4 : DFFR_X1 port map( D => n14155, CK => clk, RN => n21210, 
                           Q => n19171, QN => n_1241);
   clk_r_REG11220_S4 : DFFS_X1 port map( D => n14154, CK => clk, SN => n21204, 
                           Q => n19170, QN => n_1242);
   clk_r_REG11114_S4 : DFFS_X1 port map( D => n14152, CK => clk, SN => n21196, 
                           Q => n19169, QN => n_1243);
   clk_r_REG10646_S5 : DFFR_X1 port map( D => n14150, CK => clk, RN => n21193, 
                           Q => n19168, QN => n_1244);
   clk_r_REG10739_S5 : DFFR_X1 port map( D => n14149, CK => clk, RN => n21193, 
                           Q => n19167, QN => n_1245);
   clk_r_REG10751_S4 : DFFS_X1 port map( D => n17479, CK => clk, SN => n21202, 
                           Q => n19166, QN => n_1246);
   clk_r_REG10734_S5 : DFFR_X1 port map( D => n17504, CK => clk, RN => n21195, 
                           Q => n19165, QN => n_1247);
   clk_r_REG10774_S11 : DFFS_X1 port map( D => n17527, CK => clk, SN => n21195,
                           Q => n19164, QN => n_1248);
   clk_r_REG10747_S5 : DFFR_X1 port map( D => n14144, CK => clk, RN => n21210, 
                           Q => n19163, QN => n_1249);
   clk_r_REG10662_S5 : DFFR_X1 port map( D => n14143, CK => clk, RN => n21189, 
                           Q => n19162, QN => n_1250);
   clk_r_REG10667_S5 : DFFR_X1 port map( D => n14142, CK => clk, RN => n21189, 
                           Q => n19161, QN => n_1251);
   clk_r_REG10717_S6 : DFFR_X1 port map( D => n14249, CK => clk, RN => n21191, 
                           Q => n19158, QN => n_1252);
   clk_r_REG10718_S6 : DFFR_X1 port map( D => n14248, CK => clk, RN => n21194, 
                           Q => n19157, QN => n_1253);
   clk_r_REG10719_S6 : DFFR_X1 port map( D => n14247, CK => clk, RN => n21201, 
                           Q => n19156, QN => n_1254);
   clk_r_REG10720_S6 : DFFR_X1 port map( D => n14246, CK => clk, RN => n21211, 
                           Q => n19155, QN => n_1255);
   clk_r_REG10721_S6 : DFFR_X1 port map( D => n14245, CK => clk, RN => n21191, 
                           Q => n19154, QN => n_1256);
   clk_r_REG10722_S6 : DFFR_X1 port map( D => n14244, CK => clk, RN => n21198, 
                           Q => n19153, QN => n_1257);
   clk_r_REG10723_S6 : DFFR_X1 port map( D => n14243, CK => clk, RN => n21194, 
                           Q => n19152, QN => n_1258);
   clk_r_REG10724_S6 : DFFR_X1 port map( D => n14242, CK => clk, RN => n21191, 
                           Q => n19151, QN => n_1259);
   clk_r_REG10725_S6 : DFFR_X1 port map( D => n14241, CK => clk, RN => n21208, 
                           Q => n19150, QN => n_1260);
   clk_r_REG10649_S5 : DFFR_X1 port map( D => n14240, CK => clk, RN => n21203, 
                           Q => n19149, QN => n_1261);
   clk_r_REG10666_S5 : DFFR_X1 port map( D => n13897, CK => clk, RN => n21210, 
                           Q => n19148, QN => n_1262);
   clk_r_REG11579_S5 : DFFR_X1 port map( D => n14140, CK => clk, RN => n21197, 
                           Q => n19147, QN => n_1263);
   clk_r_REG11165_S4 : DFFR_X1 port map( D => n21174, CK => clk, RN => n21211, 
                           Q => n22961, QN => n19146);
   clk_r_REG10797_S5 : DFFS_X1 port map( D => n21183, CK => clk, SN => n21205, 
                           Q => n_1264, QN => n19145);
   clk_r_REG11248_S4 : DFFR_X1 port map( D => n1845, CK => clk, RN => n21197, Q
                           => n_1265, QN => n19144);
   clk_r_REG11245_S4 : DFFR_X1 port map( D => n1847, CK => clk, RN => n21190, Q
                           => n22988, QN => n19143);
   clk_r_REG11189_S4 : DFFR_X1 port map( D => n1838, CK => clk, RN => n21190, Q
                           => n22976, QN => n19142);
   clk_r_REG11200_S4 : DFFS_X1 port map( D => n1844, CK => clk, SN => n21205, Q
                           => n22959, QN => n19141);
   clk_r_REG11570_S5 : DFFR_X1 port map( D => n14123, CK => clk, RN => n21203, 
                           Q => n19140, QN => n_1266);
   clk_r_REG11571_S6 : DFFR_X1 port map( D => n19140, CK => clk, RN => n21205, 
                           Q => n19139, QN => n_1267);
   clk_r_REG11572_S7 : DFFR_X1 port map( D => n19139, CK => clk, RN => n21211, 
                           Q => n19138, QN => n_1268);
   clk_r_REG11573_S8 : DFFR_X1 port map( D => n19138, CK => clk, RN => n21211, 
                           Q => n19137, QN => n_1269);
   clk_r_REG11574_S9 : DFFR_X1 port map( D => n19137, CK => clk, RN => n21205, 
                           Q => n19136, QN => n_1270);
   clk_r_REG11575_S10 : DFFR_X1 port map( D => n19136, CK => clk, RN => n21192,
                           Q => n19135, QN => n_1271);
   clk_r_REG11281_S5 : DFFR_X1 port map( D => n14122, CK => clk, RN => n21204, 
                           Q => n19134, QN => n_1272);
   clk_r_REG11282_S5 : DFFR_X1 port map( D => n14121, CK => clk, RN => n21198, 
                           Q => n19133, QN => n_1273);
   clk_r_REG11280_S5 : DFFR_X1 port map( D => n14120, CK => clk, RN => n21192, 
                           Q => n19132, QN => n_1274);
   clk_r_REG10888_S5 : DFFR_X1 port map( D => n14119, CK => clk, RN => n21208, 
                           Q => n19131, QN => n_1275);
   clk_r_REG10851_S5 : DFFR_X1 port map( D => n14118, CK => clk, RN => n21209, 
                           Q => n19130, QN => n_1276);
   clk_r_REG10768_S5 : DFFR_X1 port map( D => n14117, CK => clk, RN => n21205, 
                           Q => n19129, QN => n_1277);
   clk_r_REG10703_S5 : DFFR_X1 port map( D => n14116, CK => clk, RN => n21209, 
                           Q => n19128, QN => n_1278);
   clk_r_REG10702_S5 : DFFR_X1 port map( D => n14115, CK => clk, RN => n21193, 
                           Q => n19127, QN => n_1279);
   clk_r_REG10700_S5 : DFFR_X1 port map( D => n14114, CK => clk, RN => n21204, 
                           Q => n19126, QN => n_1280);
   clk_r_REG10663_S5 : DFFR_X1 port map( D => n14113, CK => clk, RN => n21201, 
                           Q => n19125, QN => n_1281);
   clk_r_REG10659_S5 : DFFR_X1 port map( D => n14112, CK => clk, RN => n21209, 
                           Q => n19124, QN => n_1282);
   clk_r_REG10334_S5 : DFFR_X1 port map( D => n14111, CK => clk, RN => n21203, 
                           Q => n19123, QN => n_1283);
   clk_r_REG10655_S5 : DFFR_X1 port map( D => n14110, CK => clk, RN => n21206, 
                           Q => n19122, QN => n_1284);
   clk_r_REG10657_S5 : DFFR_X1 port map( D => n14109, CK => clk, RN => n21196, 
                           Q => n19121, QN => n_1285);
   clk_r_REG10658_S6 : DFFR_X1 port map( D => n19121, CK => clk, RN => n21206, 
                           Q => n19120, QN => n_1286);
   clk_r_REG10799_S6 : DFFR_X1 port map( D => n14103, CK => clk, RN => n21193, 
                           Q => n19119, QN => n_1287);
   clk_r_REG10800_S7 : DFFR_X1 port map( D => n19119, CK => clk, RN => n21190, 
                           Q => n19118, QN => n_1288);
   clk_r_REG10801_S8 : DFFR_X1 port map( D => n19118, CK => clk, RN => n21195, 
                           Q => n19117, QN => n_1289);
   clk_r_REG10802_S9 : DFFR_X1 port map( D => n19117, CK => clk, RN => n21205, 
                           Q => n19116, QN => n_1290);
   clk_r_REG10803_S10 : DFFR_X1 port map( D => n19116, CK => clk, RN => n21189,
                           Q => n19115, QN => n_1291);
   clk_r_REG10653_S5 : DFFR_X1 port map( D => n14101, CK => clk, RN => n21200, 
                           Q => n19114, QN => n_1292);
   clk_r_REG10654_S5 : DFFR_X1 port map( D => n14100, CK => clk, RN => n21205, 
                           Q => n19113, QN => n_1293);
   clk_r_REG10818_S6 : DFFR_X1 port map( D => n14095, CK => clk, RN => n21210, 
                           Q => n19112, QN => n_1294);
   clk_r_REG10819_S7 : DFFR_X1 port map( D => n19112, CK => clk, RN => n21196, 
                           Q => n19111, QN => n_1295);
   clk_r_REG10820_S8 : DFFR_X1 port map( D => n19111, CK => clk, RN => n21207, 
                           Q => n19110, QN => n_1296);
   clk_r_REG10821_S9 : DFFR_X1 port map( D => n19110, CK => clk, RN => n21193, 
                           Q => n19109, QN => n_1297);
   clk_r_REG10822_S10 : DFFR_X1 port map( D => n19109, CK => clk, RN => n21211,
                           Q => n19108, QN => n_1298);
   clk_r_REG10656_S6 : DFFR_X1 port map( D => n14093, CK => clk, RN => n21204, 
                           Q => n19107, QN => n_1299);
   clk_r_REG10651_S5 : DFFR_X1 port map( D => n4009, CK => clk, RN => n21192, Q
                           => n19106, QN => n_1300);
   clk_r_REG10652_S5 : DFFR_X1 port map( D => n4008, CK => clk, RN => n21207, Q
                           => n19105, QN => n_1301);
   clk_r_REG10832_S6 : DFFR_X1 port map( D => n14088, CK => clk, RN => n21194, 
                           Q => n19104, QN => n_1302);
   clk_r_REG10833_S7 : DFFR_X1 port map( D => n19104, CK => clk, RN => n21201, 
                           Q => n19103, QN => n_1303);
   clk_r_REG10834_S8 : DFFR_X1 port map( D => n19103, CK => clk, RN => n21190, 
                           Q => n19102, QN => n_1304);
   clk_r_REG10835_S9 : DFFR_X1 port map( D => n19102, CK => clk, RN => n21203, 
                           Q => n19101, QN => n_1305);
   clk_r_REG10836_S10 : DFFR_X1 port map( D => n19101, CK => clk, RN => n21202,
                           Q => n19100, QN => n_1306);
   clk_r_REG10660_S6 : DFFR_X1 port map( D => n14087, CK => clk, RN => n21195, 
                           Q => n19099, QN => n_1307);
   clk_r_REG10335_S6 : DFFR_X1 port map( D => n14086, CK => clk, RN => n21208, 
                           Q => n19098, QN => n_1308);
   clk_r_REG10336_S6 : DFFR_X1 port map( D => n14085, CK => clk, RN => n21196, 
                           Q => n19097, QN => n_1309);
   clk_r_REG10704_S6 : DFFR_X1 port map( D => n14080, CK => clk, RN => n21194, 
                           Q => n19096, QN => n_1310);
   clk_r_REG10705_S7 : DFFR_X1 port map( D => n19096, CK => clk, RN => n21197, 
                           Q => n19095, QN => n_1311);
   clk_r_REG10706_S8 : DFFR_X1 port map( D => n19095, CK => clk, RN => n21197, 
                           Q => n19094, QN => n_1312);
   clk_r_REG10707_S9 : DFFR_X1 port map( D => n19094, CK => clk, RN => n21192, 
                           Q => n19093, QN => n_1313);
   clk_r_REG10708_S10 : DFFR_X1 port map( D => n19093, CK => clk, RN => n21190,
                           Q => n19092, QN => n_1314);
   clk_r_REG10701_S6 : DFFR_X1 port map( D => n14078, CK => clk, RN => n21209, 
                           Q => n19091, QN => n_1315);
   clk_r_REG10664_S6 : DFFR_X1 port map( D => n14077, CK => clk, RN => n21205, 
                           Q => n19090, QN => n_1316);
   clk_r_REG10665_S6 : DFFR_X1 port map( D => n14076, CK => clk, RN => n21209, 
                           Q => n19089, QN => n_1317);
   clk_r_REG10535_S7 : DFFR_X1 port map( D => n14070, CK => clk, RN => n21191, 
                           Q => n19088, QN => n_1318);
   clk_r_REG10536_S8 : DFFR_X1 port map( D => n19088, CK => clk, RN => n21202, 
                           Q => n19087, QN => n_1319);
   clk_r_REG10537_S9 : DFFR_X1 port map( D => n19087, CK => clk, RN => n21196, 
                           Q => n19086, QN => n_1320);
   clk_r_REG10538_S10 : DFFR_X1 port map( D => n19086, CK => clk, RN => n21209,
                           Q => n19085, QN => n_1321);
   clk_r_REG10564_S7 : DFFR_X1 port map( D => n14057, CK => clk, RN => n21202, 
                           Q => n19084, QN => n_1322);
   clk_r_REG10549_S7 : DFFR_X1 port map( D => n14056, CK => clk, RN => n21192, 
                           Q => n19083, QN => n_1323);
   clk_r_REG10613_S7 : DFFR_X1 port map( D => n14053, CK => clk, RN => n21209, 
                           Q => n19082, QN => n_1324);
   clk_r_REG10614_S8 : DFFR_X1 port map( D => n19082, CK => clk, RN => n21210, 
                           Q => n19081, QN => n_1325);
   clk_r_REG10615_S9 : DFFR_X1 port map( D => n19081, CK => clk, RN => n21191, 
                           Q => n19080, QN => n_1326);
   clk_r_REG10616_S10 : DFFR_X1 port map( D => n19080, CK => clk, RN => n21210,
                           Q => n19079, QN => n_1327);
   clk_r_REG10337_S7 : DFFR_X1 port map( D => n14050, CK => clk, RN => n21192, 
                           Q => n19078, QN => n_1328);
   clk_r_REG10338_S8 : DFFR_X1 port map( D => n19078, CK => clk, RN => n21210, 
                           Q => n19077, QN => n_1329);
   clk_r_REG10339_S9 : DFFR_X1 port map( D => n19077, CK => clk, RN => n21212, 
                           Q => n19076, QN => n_1330);
   clk_r_REG10340_S10 : DFFR_X1 port map( D => n19076, CK => clk, RN => n21210,
                           Q => n19075, QN => n_1331);
   clk_r_REG10606_S7 : DFFR_X1 port map( D => n14047, CK => clk, RN => n21209, 
                           Q => n19074, QN => n_1332);
   clk_r_REG10607_S8 : DFFR_X1 port map( D => n19074, CK => clk, RN => n21212, 
                           Q => n19073, QN => n_1333);
   clk_r_REG10608_S9 : DFFR_X1 port map( D => n19073, CK => clk, RN => n21209, 
                           Q => n19072, QN => n_1334);
   clk_r_REG10609_S10 : DFFR_X1 port map( D => n19072, CK => clk, RN => n21201,
                           Q => n19071, QN => n_1335);
   clk_r_REG10600_S7 : DFFR_X1 port map( D => n14044, CK => clk, RN => n21193, 
                           Q => n19070, QN => n_1336);
   clk_r_REG10601_S8 : DFFR_X1 port map( D => n19070, CK => clk, RN => n21208, 
                           Q => n19069, QN => n_1337);
   clk_r_REG10602_S9 : DFFR_X1 port map( D => n19069, CK => clk, RN => n21195, 
                           Q => n19068, QN => n_1338);
   clk_r_REG10603_S10 : DFFR_X1 port map( D => n19068, CK => clk, RN => n21193,
                           Q => n19067, QN => n_1339);
   clk_r_REG10594_S7 : DFFR_X1 port map( D => n14041, CK => clk, RN => n21199, 
                           Q => n19066, QN => n_1340);
   clk_r_REG10595_S8 : DFFR_X1 port map( D => n19066, CK => clk, RN => n21212, 
                           Q => n19065, QN => n_1341);
   clk_r_REG10596_S9 : DFFR_X1 port map( D => n19065, CK => clk, RN => n21191, 
                           Q => n19064, QN => n_1342);
   clk_r_REG10597_S10 : DFFR_X1 port map( D => n19064, CK => clk, RN => n21209,
                           Q => n19063, QN => n_1343);
   clk_r_REG10589_S7 : DFFR_X1 port map( D => n14038, CK => clk, RN => n21194, 
                           Q => n19062, QN => n_1344);
   clk_r_REG10590_S8 : DFFR_X1 port map( D => n19062, CK => clk, RN => n21208, 
                           Q => n19061, QN => n_1345);
   clk_r_REG10591_S9 : DFFR_X1 port map( D => n19061, CK => clk, RN => n21201, 
                           Q => n19060, QN => n_1346);
   clk_r_REG10592_S10 : DFFR_X1 port map( D => n19060, CK => clk, RN => n21210,
                           Q => n19059, QN => n_1347);
   clk_r_REG10583_S7 : DFFR_X1 port map( D => n14035, CK => clk, RN => n21199, 
                           Q => n19058, QN => n_1348);
   clk_r_REG10584_S8 : DFFR_X1 port map( D => n19058, CK => clk, RN => n21199, 
                           Q => n19057, QN => n_1349);
   clk_r_REG10585_S9 : DFFR_X1 port map( D => n19057, CK => clk, RN => n21189, 
                           Q => n19056, QN => n_1350);
   clk_r_REG10586_S10 : DFFR_X1 port map( D => n19056, CK => clk, RN => n21193,
                           Q => n19055, QN => n_1351);
   clk_r_REG10424_S7 : DFFR_X1 port map( D => n14032, CK => clk, RN => n21192, 
                           Q => n19054, QN => n_1352);
   clk_r_REG10425_S8 : DFFR_X1 port map( D => n19054, CK => clk, RN => n21212, 
                           Q => n19053, QN => n_1353);
   clk_r_REG10426_S9 : DFFR_X1 port map( D => n19053, CK => clk, RN => n21193, 
                           Q => n19052, QN => n_1354);
   clk_r_REG10427_S10 : DFFR_X1 port map( D => n19052, CK => clk, RN => n21193,
                           Q => n19051, QN => n_1355);
   clk_r_REG10429_S7 : DFFR_X1 port map( D => n14029, CK => clk, RN => n21206, 
                           Q => n19050, QN => n_1356);
   clk_r_REG10430_S8 : DFFR_X1 port map( D => n19050, CK => clk, RN => n21189, 
                           Q => n19049, QN => n_1357);
   clk_r_REG10431_S9 : DFFR_X1 port map( D => n19049, CK => clk, RN => n21209, 
                           Q => n19048, QN => n_1358);
   clk_r_REG10432_S10 : DFFR_X1 port map( D => n19048, CK => clk, RN => n21211,
                           Q => n19047, QN => n_1359);
   clk_r_REG10434_S7 : DFFR_X1 port map( D => n14026, CK => clk, RN => n21192, 
                           Q => n19046, QN => n_1360);
   clk_r_REG10435_S8 : DFFR_X1 port map( D => n19046, CK => clk, RN => n21191, 
                           Q => n19045, QN => n_1361);
   clk_r_REG10436_S9 : DFFR_X1 port map( D => n19045, CK => clk, RN => n21198, 
                           Q => n19044, QN => n_1362);
   clk_r_REG10437_S10 : DFFR_X1 port map( D => n19044, CK => clk, RN => n21206,
                           Q => n19043, QN => n_1363);
   clk_r_REG10438_S11 : DFFR_X1 port map( D => n19043, CK => clk, RN => n21193,
                           Q => n19042, QN => n_1364);
   clk_r_REG10575_S7 : DFFR_X1 port map( D => n14023, CK => clk, RN => n21190, 
                           Q => n19041, QN => n_1365);
   clk_r_REG10576_S8 : DFFR_X1 port map( D => n19041, CK => clk, RN => n21208, 
                           Q => n19040, QN => n_1366);
   clk_r_REG10577_S9 : DFFR_X1 port map( D => n19040, CK => clk, RN => n21193, 
                           Q => n19039, QN => n_1367);
   clk_r_REG10578_S10 : DFFR_X1 port map( D => n19039, CK => clk, RN => n21197,
                           Q => n19038, QN => n_1368);
   clk_r_REG10569_S7 : DFFR_X1 port map( D => n14022, CK => clk, RN => n21205, 
                           Q => n19037, QN => n_1369);
   clk_r_REG10570_S7 : DFFR_X1 port map( D => n14019, CK => clk, RN => n21205, 
                           Q => n19036, QN => n_1370);
   clk_r_REG10571_S8 : DFFR_X1 port map( D => n19036, CK => clk, RN => n21194, 
                           Q => n19035, QN => n_1371);
   clk_r_REG10572_S9 : DFFR_X1 port map( D => n19035, CK => clk, RN => n21210, 
                           Q => n19034, QN => n_1372);
   clk_r_REG10573_S10 : DFFR_X1 port map( D => n19034, CK => clk, RN => n21194,
                           Q => n19033, QN => n_1373);
   clk_r_REG10565_S8 : DFFR_X1 port map( D => n14017, CK => clk, RN => n21202, 
                           Q => n19032, QN => n_1374);
   clk_r_REG10566_S9 : DFFR_X1 port map( D => n19032, CK => clk, RN => n21205, 
                           Q => n19031, QN => n_1375);
   clk_r_REG10567_S10 : DFFR_X1 port map( D => n19031, CK => clk, RN => n21192,
                           Q => n19030, QN => n_1376);
   clk_r_REG10550_S8 : DFFR_X1 port map( D => n14015, CK => clk, RN => n21206, 
                           Q => n19029, QN => n_1377);
   clk_r_REG10551_S9 : DFFR_X1 port map( D => n19029, CK => clk, RN => n21192, 
                           Q => n19028, QN => n_1378);
   clk_r_REG10552_S10 : DFFR_X1 port map( D => n19028, CK => clk, RN => n21208,
                           Q => n19027, QN => n_1379);
   clk_r_REG10553_S8 : DFFR_X1 port map( D => n14013, CK => clk, RN => n21193, 
                           Q => n19026, QN => n_1380);
   clk_r_REG10554_S9 : DFFR_X1 port map( D => n19026, CK => clk, RN => n21193, 
                           Q => n19025, QN => n_1381);
   clk_r_REG10555_S10 : DFFR_X1 port map( D => n19025, CK => clk, RN => n21191,
                           Q => n19024, QN => n_1382);
   clk_r_REG10557_S8 : DFFR_X1 port map( D => n14011, CK => clk, RN => n21212, 
                           Q => n19023, QN => n_1383);
   clk_r_REG10558_S9 : DFFR_X1 port map( D => n19023, CK => clk, RN => n21211, 
                           Q => n19022, QN => n_1384);
   clk_r_REG10559_S10 : DFFR_X1 port map( D => n19022, CK => clk, RN => n21211,
                           Q => n19021, QN => n_1385);
   clk_r_REG10560_S8 : DFFR_X1 port map( D => n14009, CK => clk, RN => n21199, 
                           Q => n19020, QN => n_1386);
   clk_r_REG10561_S9 : DFFR_X1 port map( D => n19020, CK => clk, RN => n21190, 
                           Q => n19019, QN => n_1387);
   clk_r_REG10562_S10 : DFFR_X1 port map( D => n19019, CK => clk, RN => n21200,
                           Q => n19018, QN => n_1388);
   clk_r_REG10632_S4 : DFFR_X1 port map( D => n22998, CK => clk, RN => n21193, 
                           Q => n19017, QN => n_1389);
   clk_r_REG10475_S5 : DFFR_X1 port map( D => n1778, CK => clk, RN => n21210, Q
                           => n_1390, QN => n19016);
   clk_r_REG11004_S4 : DFFS_X1 port map( D => n1810, CK => clk, SN => n21195, Q
                           => n_1391, QN => n19015);
   clk_r_REG10755_S4 : DFFS_X1 port map( D => n1803, CK => clk, SN => n21205, Q
                           => n_1392, QN => n19014);
   clk_r_REG10787_S4 : DFFS_X1 port map( D => n12526, CK => clk, SN => n21206, 
                           Q => n19013, QN => n_1393);
   clk_r_REG10994_S15 : DFFS_X1 port map( D => n1824, CK => clk, SN => n21203, 
                           Q => n_1394, QN => n19012);
   clk_r_REG10991_S4 : DFFS_X1 port map( D => n1828, CK => clk, SN => n21205, Q
                           => n_1395, QN => n19011);
   clk_r_REG11277_S3 : DFFR_X1 port map( D => n13984, CK => clk, RN => rst_BAR,
                           Q => n19010, QN => n_1396);
   clk_r_REG10753_S4 : DFFS_X1 port map( D => n1802, CK => clk, SN => n21208, Q
                           => n_1397, QN => n19009);
   clk_r_REG10996_S15 : DFFR_X1 port map( D => n1822, CK => clk, RN => n21211, 
                           Q => n_1398, QN => n19008);
   clk_r_REG10858_S4 : DFFR_X1 port map( D => n1806, CK => clk, RN => n21200, Q
                           => n_1399, QN => n19007);
   clk_r_REG10789_S4 : DFFS_X1 port map( D => n1807, CK => clk, SN => n21197, Q
                           => n_1400, QN => n19006);
   clk_r_REG10680_S4 : DFFS_X1 port map( D => n16696, CK => clk, SN => n21207, 
                           Q => n19005, QN => n_1401);
   clk_r_REG10689_S4 : DFFR_X1 port map( D => n16695, CK => clk, RN => n21200, 
                           Q => n19004, QN => n_1402);
   clk_r_REG10683_S4 : DFFR_X1 port map( D => n16700, CK => clk, RN => n21206, 
                           Q => n19003, QN => n_1403);
   clk_r_REG10676_S4 : DFFR_X1 port map( D => n16698, CK => clk, RN => n21195, 
                           Q => n_1404, QN => n21168);
   clk_r_REG10681_S4 : DFFR_X1 port map( D => n16702, CK => clk, RN => n21192, 
                           Q => n19001, QN => n_1405);
   clk_r_REG10691_S4 : DFFR_X1 port map( D => n16705, CK => clk, RN => n21196, 
                           Q => n19000, QN => n_1406);
   clk_r_REG10690_S4 : DFFR_X1 port map( D => n16706, CK => clk, RN => n21197, 
                           Q => n18999, QN => n_1407);
   clk_r_REG10508_S4 : DFFR_X1 port map( D => n16709, CK => clk, RN => n21189, 
                           Q => n18998, QN => n_1408);
   clk_r_REG10752_S4 : DFFS_X1 port map( D => n16713, CK => clk, SN => n21197, 
                           Q => n18997, QN => n_1409);
   clk_r_REG10985_S4 : DFFR_X1 port map( D => n14004, CK => clk, RN => n21194, 
                           Q => n18996, QN => n_1410);
   clk_r_REG10987_S4 : DFFS_X1 port map( D => n14000, CK => clk, SN => n21202, 
                           Q => n18995, QN => n_1411);
   clk_r_REG10980_S15 : DFFR_X1 port map( D => n14003, CK => clk, RN => n21190,
                           Q => n18994, QN => n_1412);
   clk_r_REG10983_S15 : DFFS_X1 port map( D => n13999, CK => clk, SN => n21205,
                           Q => n18993, QN => n_1413);
   clk_r_REG10988_S15 : DFFS_X1 port map( D => n11449, CK => clk, SN => n21209,
                           Q => n18992, QN => n_1414);
   clk_r_REG10990_S15 : DFFR_X1 port map( D => n13997, CK => clk, RN => n21192,
                           Q => n18991, QN => n_1415);
   clk_r_REG10989_S15 : DFFR_X1 port map( D => n13992, CK => clk, RN => n21197,
                           Q => n18990, QN => n_1416);
   clk_r_REG10992_S4 : DFFS_X1 port map( D => n13990, CK => clk, SN => n21201, 
                           Q => n18989, QN => n_1417);
   clk_r_REG10984_S15 : DFFS_X1 port map( D => n13989, CK => clk, SN => n21195,
                           Q => n18988, QN => n_1418);
   clk_r_REG11003_S4 : DFFR_X1 port map( D => n13988, CK => clk, RN => n21193, 
                           Q => n18987, QN => n_1419);
   clk_r_REG11002_S4 : DFFR_X1 port map( D => n13987, CK => clk, RN => n21211, 
                           Q => n18986, QN => n_1420);
   clk_r_REG11014_S4 : DFFS_X1 port map( D => n16766, CK => clk, SN => n21205, 
                           Q => n18985, QN => n_1421);
   clk_r_REG10414_S4 : DFFS_X1 port map( D => n16770, CK => clk, SN => n21207, 
                           Q => n18984, QN => n_1422);
   clk_r_REG10520_S4 : DFFR_X1 port map( D => n16771, CK => clk, RN => n21203, 
                           Q => n18983, QN => n_1423);
   clk_r_REG10981_S15 : DFFS_X1 port map( D => n16783, CK => clk, SN => n21203,
                           Q => n18982, QN => n_1424);
   clk_r_REG10986_S4 : DFFS_X1 port map( D => n16782, CK => clk, SN => n21207, 
                           Q => n18981, QN => n_1425);
   clk_r_REG10876_S11 : DFFS_X1 port map( D => n13980, CK => clk, SN => n21202,
                           Q => n18980, QN => n_1426);
   clk_r_REG10885_S5 : DFFS_X1 port map( D => n13978, CK => clk, SN => n21204, 
                           Q => n18979, QN => n_1427);
   clk_r_REG10999_S4 : DFFR_X1 port map( D => n16808, CK => clk, RN => n21201, 
                           Q => n18978, QN => n_1428);
   clk_r_REG10993_S4 : DFFS_X1 port map( D => n16807, CK => clk, SN => n21198, 
                           Q => n18977, QN => n_1429);
   clk_r_REG11171_S4 : DFFS_X1 port map( D => n13977, CK => clk, SN => n21196, 
                           Q => n18976, QN => n_1430);
   clk_r_REG10998_S4 : DFFR_X1 port map( D => n16831, CK => clk, RN => n21191, 
                           Q => n18975, QN => n_1431);
   clk_r_REG11215_S4 : DFFS_X1 port map( D => n13974, CK => clk, SN => n21198, 
                           Q => n18974, QN => n_1432);
   clk_r_REG10804_S11 : DFFS_X1 port map( D => n13973, CK => clk, SN => n21198,
                           Q => n18973, QN => n_1433);
   clk_r_REG11169_S5 : DFFS_X1 port map( D => n13972, CK => clk, SN => n21197, 
                           Q => n18972, QN => n_1434);
   clk_r_REG11000_S4 : DFFS_X1 port map( D => n13971, CK => clk, SN => n21197, 
                           Q => n18971, QN => n_1435);
   clk_r_REG10693_S4 : DFFR_X1 port map( D => n16857, CK => clk, RN => n21198, 
                           Q => n18970, QN => n_1436);
   clk_r_REG11578_S5 : DFFS_X1 port map( D => n13970, CK => clk, SN => n21198, 
                           Q => n18969, QN => n_1437);
   clk_r_REG11164_S11 : DFFS_X1 port map( D => n13969, CK => clk, SN => n21197,
                           Q => n18968, QN => n_1438);
   clk_r_REG11577_S5 : DFFR_X1 port map( D => n13968, CK => clk, RN => n21196, 
                           Q => n18967, QN => n_1439);
   clk_r_REG11005_S4 : DFFS_X1 port map( D => n13967, CK => clk, SN => n21198, 
                           Q => n18966, QN => n_1440);
   clk_r_REG11216_S4 : DFFS_X1 port map( D => n13966, CK => clk, SN => n21198, 
                           Q => n18965, QN => n_1441);
   clk_r_REG11576_S4 : DFFS_X1 port map( D => n13965, CK => clk, SN => n21197, 
                           Q => n18964, QN => n_1442);
   clk_r_REG10857_S4 : DFFR_X1 port map( D => n13964, CK => clk, RN => n21212, 
                           Q => n18963, QN => n_1443);
   clk_r_REG10862_S4 : DFFR_X1 port map( D => n16909, CK => clk, RN => n21209, 
                           Q => n18962, QN => n_1444);
   clk_r_REG10509_S4 : DFFR_X1 port map( D => n11966, CK => clk, RN => n21201, 
                           Q => n18961, QN => n_1445);
   clk_r_REG10512_S4 : DFFS_X1 port map( D => n13956, CK => clk, SN => n21197, 
                           Q => n18960, QN => n_1446);
   clk_r_REG10511_S4 : DFFS_X1 port map( D => n13955, CK => clk, SN => n21208, 
                           Q => n18959, QN => n_1447);
   clk_r_REG10513_S4 : DFFS_X1 port map( D => n13954, CK => clk, SN => n21199, 
                           Q => n18958, QN => n_1448);
   clk_r_REG10510_S4 : DFFS_X1 port map( D => n13953, CK => clk, SN => n21208, 
                           Q => n18957, QN => n_1449);
   clk_r_REG10685_S4 : DFFS_X1 port map( D => n13963, CK => clk, SN => n21208, 
                           Q => n18956, QN => n_1450);
   clk_r_REG10684_S4 : DFFR_X1 port map( D => n13950, CK => clk, RN => n21198, 
                           Q => n18955, QN => n_1451);
   clk_r_REG11015_S4 : DFFS_X1 port map( D => n13949, CK => clk, SN => n21200, 
                           Q => n18954, QN => n_1452);
   clk_r_REG10677_S4 : DFFS_X1 port map( D => n1805, CK => clk, SN => n21200, Q
                           => n_1453, QN => n18953);
   clk_r_REG10678_S4 : DFFS_X1 port map( D => n13947, CK => clk, SN => n21208, 
                           Q => n18952, QN => n_1454);
   clk_r_REG10686_S4 : DFFR_X1 port map( D => n13946, CK => clk, RN => n21209, 
                           Q => n18951, QN => n_1455);
   clk_r_REG10688_S4 : DFFR_X1 port map( D => n13945, CK => clk, RN => n21207, 
                           Q => n18950, QN => n_1456);
   clk_r_REG10687_S4 : DFFR_X1 port map( D => n13944, CK => clk, RN => n21210, 
                           Q => n18949, QN => n_1457);
   clk_r_REG10756_S4 : DFFR_X1 port map( D => n13943, CK => clk, RN => n21191, 
                           Q => n18948, QN => n_1458);
   clk_r_REG10517_S4 : DFFR_X1 port map( D => n13941, CK => clk, RN => n21189, 
                           Q => n18947, QN => n_1459);
   clk_r_REG11031_S4 : DFFS_X1 port map( D => n13940, CK => clk, SN => n21202, 
                           Q => n18946, QN => n_1460);
   clk_r_REG10365_S5 : DFFS_X1 port map( D => n14165, CK => clk, SN => n21208, 
                           Q => n18945, QN => n_1461);
   clk_r_REG10505_S4 : DFFR_X1 port map( D => n17012, CK => clk, RN => n21191, 
                           Q => n18944, QN => n_1462);
   clk_r_REG10682_S4 : DFFR_X1 port map( D => n17011, CK => clk, RN => n21207, 
                           Q => n18943, QN => n_1463);
   clk_r_REG10501_S4 : DFFS_X1 port map( D => n17016, CK => clk, SN => n21196, 
                           Q => n18942, QN => n_1464);
   clk_r_REG10504_S4 : DFFR_X1 port map( D => n17018, CK => clk, RN => n21200, 
                           Q => n18941, QN => n_1465);
   clk_r_REG10499_S4 : DFFS_X1 port map( D => n17017, CK => clk, SN => n21200, 
                           Q => n18940, QN => n_1466);
   clk_r_REG10506_S4 : DFFR_X1 port map( D => n17020, CK => clk, RN => n21197, 
                           Q => n18939, QN => n_1467);
   clk_r_REG10503_S4 : DFFR_X1 port map( D => n17019, CK => clk, RN => n21200, 
                           Q => n18938, QN => n_1468);
   clk_r_REG10514_S4 : DFFR_X1 port map( D => n17068, CK => clk, RN => n21190, 
                           Q => n18937, QN => n_1469);
   clk_r_REG10516_S4 : DFFR_X1 port map( D => n17089, CK => clk, RN => n21195, 
                           Q => n18936, QN => n_1470);
   clk_r_REG10375_S4 : DFFR_X1 port map( D => n13938, CK => clk, RN => n21193, 
                           Q => n18935, QN => n_1471);
   clk_r_REG11217_S4 : DFFS_X1 port map( D => n13936, CK => clk, SN => n21197, 
                           Q => n18934, QN => n_1472);
   clk_r_REG11722_S11 : DFFS_X1 port map( D => n13935, CK => clk, SN => n21202,
                           Q => n18933, QN => n_1473);
   clk_r_REG10761_S4 : DFFR_X1 port map( D => n13933, CK => clk, RN => n21212, 
                           Q => n18932, QN => n_1474);
   clk_r_REG10859_S4 : DFFR_X1 port map( D => n17160, CK => clk, RN => n21190, 
                           Q => n18931, QN => n_1475);
   clk_r_REG10556_S11 : DFFS_X1 port map( D => n13932, CK => clk, SN => n21201,
                           Q => n18930, QN => n_1476);
   clk_r_REG11076_S4 : DFFS_X1 port map( D => n13931, CK => clk, SN => n21203, 
                           Q => n18929, QN => n_1477);
   clk_r_REG10356_S5 : DFFR_X1 port map( D => n13930, CK => clk, RN => n21211, 
                           Q => n18928, QN => n_1478);
   clk_r_REG10476_S4 : DFFS_X1 port map( D => n14163, CK => clk, SN => n21195, 
                           Q => n18927, QN => n_1479);
   clk_r_REG10461_S5 : DFFS_X1 port map( D => n13928, CK => clk, SN => n21196, 
                           Q => n18926, QN => n_1480);
   clk_r_REG10454_S5 : DFFS_X1 port map( D => n13927, CK => clk, SN => n21200, 
                           Q => n18925, QN => n_1481);
   clk_r_REG11041_S4 : DFFR_X1 port map( D => n17269, CK => clk, RN => n21210, 
                           Q => n18924, QN => n_1482);
   clk_r_REG10402_S5 : DFFR_X1 port map( D => n14264, CK => clk, RN => n21208, 
                           Q => n18923, QN => n_1483);
   clk_r_REG10428_S11 : DFFS_X1 port map( D => n13924, CK => clk, SN => n21205,
                           Q => n18922, QN => n_1484);
   clk_r_REG10387_S4 : DFFS_X1 port map( D => n13985, CK => clk, SN => n21207, 
                           Q => n18921, QN => n_1485);
   clk_r_REG11864_S11 : DFFS_X1 port map( D => n13922, CK => clk, SN => n21204,
                           Q => n18920, QN => n_1486);
   clk_r_REG10856_S4 : DFFR_X1 port map( D => n17360, CK => clk, RN => n21198, 
                           Q => n18919, QN => n_1487);
   clk_r_REG10760_S4 : DFFR_X1 port map( D => n17359, CK => clk, RN => n21193, 
                           Q => n18918, QN => n_1488);
   clk_r_REG10306_S5 : DFFR_X1 port map( D => n13919, CK => clk, RN => n21192, 
                           Q => n18917, QN => n_1489);
   clk_r_REG10604_S11 : DFFS_X1 port map( D => n14262, CK => clk, SN => n21207,
                           Q => n18916, QN => n_1490);
   clk_r_REG10610_S11 : DFFS_X1 port map( D => n13918, CK => clk, SN => n21207,
                           Q => n18915, QN => n_1491);
   clk_r_REG10348_S5 : DFFR_X1 port map( D => n13917, CK => clk, RN => n21193, 
                           Q => n18914, QN => n_1492);
   clk_r_REG10355_S5 : DFFR_X1 port map( D => n13916, CK => clk, RN => n21194, 
                           Q => n18913, QN => n_1493);
   clk_r_REG10341_S11 : DFFS_X1 port map( D => n13915, CK => clk, SN => n21202,
                           Q => n18912, QN => n_1494);
   clk_r_REG10631_S5 : DFFS_X1 port map( D => n14151, CK => clk, SN => n21195, 
                           Q => n18911, QN => n_1495);
   clk_r_REG10617_S11 : DFFS_X1 port map( D => n13914, CK => clk, SN => n21196,
                           Q => n18910, QN => n_1496);
   clk_r_REG10633_S4 : DFFR_X1 port map( D => n13913, CK => clk, RN => n21212, 
                           Q => n18909, QN => n_1497);
   clk_r_REG10738_S5 : DFFS_X1 port map( D => n13912, CK => clk, SN => n21205, 
                           Q => n18908, QN => n_1498);
   clk_r_REG11129_S4 : DFFS_X1 port map( D => n14261, CK => clk, SN => n21205, 
                           Q => n18907, QN => n_1499);
   clk_r_REG10709_S11 : DFFS_X1 port map( D => n13910, CK => clk, SN => n21194,
                           Q => n_1500, QN => n22996);
   clk_r_REG10758_S4 : DFFS_X1 port map( D => n17505, CK => clk, SN => n21202, 
                           Q => n18905, QN => n_1501);
   clk_r_REG10333_S11 : DFFS_X1 port map( D => n13908, CK => clk, SN => n21203,
                           Q => n18904, QN => n_1502);
   clk_r_REG10372_S4 : DFFR_X1 port map( D => n13907, CK => clk, RN => n21194, 
                           Q => n18903, QN => n_1503);
   clk_r_REG10854_S4 : DFFS_X1 port map( D => n17735, CK => clk, SN => n21198, 
                           Q => n18902, QN => n_1504);
   clk_r_REG10855_S4 : DFFR_X1 port map( D => n17734, CK => clk, RN => n21203, 
                           Q => n18901, QN => n_1505);
   clk_r_REG10759_S4 : DFFR_X1 port map( D => n17733, CK => clk, RN => n21193, 
                           Q => n18900, QN => n_1506);
   clk_r_REG10831_S6 : DFFR_X1 port map( D => n13904, CK => clk, RN => n21190, 
                           Q => n18899, QN => n_1507);
   clk_r_REG10784_S5 : DFFR_X1 port map( D => n13903, CK => clk, RN => n21209, 
                           Q => n18898, QN => n_1508);
   clk_r_REG10743_S5 : DFFR_X1 port map( D => n13902, CK => clk, RN => n21209, 
                           Q => n18897, QN => n_1509);
   clk_r_REG10744_S5 : DFFR_X1 port map( D => n13901, CK => clk, RN => n21189, 
                           Q => n18896, QN => n_1510);
   clk_r_REG10746_S5 : DFFR_X1 port map( D => n13900, CK => clk, RN => n21198, 
                           Q => n18895, QN => n_1511);
   clk_r_REG10650_S5 : DFFR_X1 port map( D => n13899, CK => clk, RN => n21210, 
                           Q => n18894, QN => n_1512);
   clk_r_REG10661_S5 : DFFR_X1 port map( D => n13898, CK => clk, RN => n21191, 
                           Q => n18893, QN => n_1513);
   clk_r_REG10563_S6 : DFFR_X1 port map( D => n13896, CK => clk, RN => n21209, 
                           Q => n18892, QN => n_1514);
   clk_r_REG11183_S4 : DFFR_X1 port map( D => n21172, CK => clk, RN => n21191, 
                           Q => n_1515, QN => n18891);
   clk_r_REG11182_S4 : DFFS_X1 port map( D => n21172, CK => clk, SN => n21201, 
                           Q => n_1516, QN => n18890);
   clk_r_REG11205_S4 : DFFS_X1 port map( D => n21171, CK => clk, SN => n21199, 
                           Q => n22968, QN => n18889);
   clk_r_REG10692_S4 : DFFR_X1 port map( D => n1830, CK => clk, RN => n21206, Q
                           => n_1517, QN => n18888);
   clk_r_REG10675_S4 : DFFS_X1 port map( D => n1831, CK => clk, SN => n21207, Q
                           => n_1518, QN => n18887);
   clk_r_REG10502_S4 : DFFS_X1 port map( D => n14407, CK => clk, SN => n21196, 
                           Q => n18886, QN => n_1519);
   clk_r_REG10519_S4 : DFFR_X1 port map( D => n1817, CK => clk, RN => n21200, Q
                           => n_1520, QN => n18885);
   clk_r_REG10412_S4 : DFFR_X1 port map( D => n1816, CK => clk, RN => n21192, Q
                           => n_1521, QN => n18884);
   clk_r_REG10479_S4 : DFFS_X1 port map( D => n1871, CK => clk, SN => n21203, Q
                           => n22980, QN => n21167);
   clk_r_REG10817_S4 : DFFS_X1 port map( D => n18133, CK => clk, SN => n21199, 
                           Q => n18882, QN => n_1522);
   clk_r_REG11001_S4 : DFFS_X1 port map( D => n14432, CK => clk, SN => n21197, 
                           Q => n18881, QN => n_1523);
   clk_r_REG10861_S4 : DFFR_X1 port map( D => n1808, CK => clk, RN => n21207, Q
                           => n_1524, QN => n18880);
   clk_r_REG10790_S4 : DFFR_X1 port map( D => n14431, CK => clk, RN => n21208, 
                           Q => n18879, QN => n_1525);
   clk_r_REG10737_S5 : DFFS_X1 port map( D => n14416, CK => clk, SN => n21203, 
                           Q => n18878, QN => n_1526);
   clk_r_REG10493_S5 : DFFS_X1 port map( D => n14452, CK => clk, SN => n21207, 
                           Q => n18877, QN => n_1527);
   clk_r_REG11159_S6 : DFFR_X1 port map( D => n13884, CK => clk, RN => n21194, 
                           Q => n18876, QN => n_1528);
   clk_r_REG11160_S7 : DFFR_X1 port map( D => n18876, CK => clk, RN => n21198, 
                           Q => n18875, QN => n_1529);
   clk_r_REG11161_S8 : DFFR_X1 port map( D => n18875, CK => clk, RN => n21192, 
                           Q => n18874, QN => n_1530);
   clk_r_REG11162_S9 : DFFR_X1 port map( D => n18874, CK => clk, RN => n21196, 
                           Q => n18873, QN => n_1531);
   clk_r_REG11163_S10 : DFFR_X1 port map( D => n18873, CK => clk, RN => n21207,
                           Q => n18872, QN => n_1532);
   clk_r_REG10812_S6 : DFFR_X1 port map( D => n13878, CK => clk, RN => n21194, 
                           Q => n18871, QN => n_1533);
   clk_r_REG10813_S7 : DFFR_X1 port map( D => n18871, CK => clk, RN => n21189, 
                           Q => n18870, QN => n_1534);
   clk_r_REG10814_S8 : DFFR_X1 port map( D => n18870, CK => clk, RN => n21200, 
                           Q => n18869, QN => n_1535);
   clk_r_REG10815_S9 : DFFR_X1 port map( D => n18869, CK => clk, RN => n21191, 
                           Q => n18868, QN => n_1536);
   clk_r_REG10816_S10 : DFFR_X1 port map( D => n18868, CK => clk, RN => n21207,
                           Q => n18867, QN => n_1537);
   clk_r_REG10528_S6 : DFFR_X1 port map( D => n13868, CK => clk, RN => n21212, 
                           Q => n18866, QN => n_1538);
   clk_r_REG10529_S7 : DFFR_X1 port map( D => n18866, CK => clk, RN => n21191, 
                           Q => n18865, QN => n_1539);
   clk_r_REG10530_S8 : DFFR_X1 port map( D => n18865, CK => clk, RN => n21197, 
                           Q => n18864, QN => n_1540);
   clk_r_REG10531_S9 : DFFR_X1 port map( D => n18864, CK => clk, RN => n21207, 
                           Q => n18863, QN => n_1541);
   clk_r_REG10532_S10 : DFFR_X1 port map( D => n18863, CK => clk, RN => n21199,
                           Q => n18862, QN => n_1542);
   clk_r_REG10533_S11 : DFFS_X1 port map( D => n18862, CK => clk, SN => n21201,
                           Q => n18861, QN => n_1543);
   clk_r_REG11865_S5 : DFFS_X1 port map( D => n13867, CK => clk, SN => n21201, 
                           Q => n18860, QN => n_1544);
   clk_r_REG10642_S7 : DFFR_X1 port map( D => n13864, CK => clk, RN => n21206, 
                           Q => n18859, QN => n_1545);
   clk_r_REG10643_S8 : DFFR_X1 port map( D => n18859, CK => clk, RN => n21212, 
                           Q => n18858, QN => n_1546);
   clk_r_REG10644_S9 : DFFR_X1 port map( D => n18858, CK => clk, RN => n21201, 
                           Q => n18857, QN => n_1547);
   clk_r_REG10645_S10 : DFFR_X1 port map( D => n18857, CK => clk, RN => n21194,
                           Q => n18856, QN => n_1548);
   clk_r_REG10740_S5 : DFFS_X1 port map( D => n13863, CK => clk, SN => n21206, 
                           Q => n18855, QN => n_1549);
   clk_r_REG10735_S5 : DFFR_X1 port map( D => n13862, CK => clk, RN => n21199, 
                           Q => n18854, QN => n_1550);
   clk_r_REG10320_S7 : DFFS_X1 port map( D => n13906, CK => clk, SN => n21206, 
                           Q => n18853, QN => n_1551);
   clk_r_REG10669_S5 : DFFR_X1 port map( D => n13861, CK => clk, RN => n21202, 
                           Q => n18852, QN => n_1552);
   clk_r_REG10733_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_13_port, CK => clk, 
                           RN => n21208, Q => n18851, QN => n_1553);
   clk_r_REG10548_S6 : DFFR_X1 port map( D => n13859, CK => clk, RN => n21206, 
                           Q => n18850, QN => n_1554);
   clk_r_REG10754_S4 : DFFR_X1 port map( D => n13858, CK => clk, RN => n21192, 
                           Q => n18849, QN => n_1555);
   clk_r_REG11218_S4 : DFFS_X1 port map( D => n13856, CK => clk, SN => n21201, 
                           Q => n18848, QN => n_1556);
   clk_r_REG10671_S5 : DFFR_X1 port map( D => n13855, CK => clk, RN => n21209, 
                           Q => n18847, QN => n_1557);
   clk_r_REG10423_S6 : DFFR_X1 port map( D => n13854, CK => clk, RN => n21199, 
                           Q => n18846, QN => n_1558);
   clk_r_REG10670_S5 : DFFR_X1 port map( D => n13860, CK => clk, RN => n21191, 
                           Q => n18845, QN => n_1559);
   clk_r_REG11858_S5 : DFFR_X1 port map( D => n13848, CK => clk, RN => n21206, 
                           Q => n18844, QN => n_1560);
   clk_r_REG11859_S6 : DFFR_X1 port map( D => n18844, CK => clk, RN => n21199, 
                           Q => n18843, QN => n_1561);
   clk_r_REG11860_S7 : DFFR_X1 port map( D => n18843, CK => clk, RN => n21212, 
                           Q => n18842, QN => n_1562);
   clk_r_REG11861_S8 : DFFR_X1 port map( D => n18842, CK => clk, RN => n21206, 
                           Q => n18841, QN => n_1563);
   clk_r_REG11862_S9 : DFFR_X1 port map( D => n18841, CK => clk, RN => n21204, 
                           Q => n18840, QN => n_1564);
   clk_r_REG11863_S10 : DFFR_X1 port map( D => n18840, CK => clk, RN => n21200,
                           Q => n18839, QN => n_1565);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n554, Q => 
                           DATA2_I_27_port);
   clk_r_REG10730_S5 : DFFS_X1 port map( D => n21185, CK => clk, SN => n21201, 
                           Q => n19415, QN => n_1566);
   clk_r_REG10845_S5 : DFFR_X1 port map( D => n21187, CK => clk, RN => n21212, 
                           Q => n19410, QN => n_1567);
   clk_r_REG10726_S5 : DFFR_X1 port map( D => n17965, CK => clk, RN => n21209, 
                           Q => n19291, QN => n_1568);
   clk_r_REG10830_S5 : DFFS_X1 port map( D => n14141, CK => clk, SN => n21201, 
                           Q => n19160, QN => n_1569);
   clk_r_REG10731_S5 : DFFR_X1 port map( D => n21162, CK => clk, RN => n21202, 
                           Q => n_1570, QN => n19159);
   clk_r_REG10716_S5 : DFFS_X1 port map( D => n17968, CK => clk, SN => n21190, 
                           Q => n19250, QN => n_1571);
   clk_r_REG10848_S5 : DFFR_X1 port map( D => n14285, CK => clk, RN => n21202, 
                           Q => n19280, QN => n_1572);
   clk_r_REG10846_S5 : DFFS_X1 port map( D => n21163, CK => clk, SN => n21195, 
                           Q => n_1573, QN => n19219);
   clk_r_REG11158_S5 : DFFR_X1 port map( D => n21188, CK => clk, RN => n21191, 
                           Q => n19413, QN => n_1574);
   clk_r_REG10870_S5 : DFFR_X1 port map( D => n14182, CK => clk, RN => n21191, 
                           Q => n19200, QN => n_1575);
   clk_r_REG11443_S5 : DFFR_X1 port map( D => n21184, CK => clk, RN => n21190, 
                           Q => n_1576, QN => n19215);
   clk_r_REG11439_S5 : DFFS_X1 port map( D => n14251, CK => clk, SN => n21197, 
                           Q => n19251, QN => n_1577);
   clk_r_REG10421_S5 : DFFS_X1 port map( D => n21186, CK => clk, SN => n21204, 
                           Q => n_1578, QN => n19217);
   U3 : CLKBUF_X1 port map( A => rst_BAR, Z => n21189);
   U4 : CLKBUF_X1 port map( A => rst_BAR, Z => n21190);
   U5 : CLKBUF_X1 port map( A => n21196, Z => n21191);
   U6 : CLKBUF_X1 port map( A => n21200, Z => n21192);
   U7 : CLKBUF_X1 port map( A => n21201, Z => n21193);
   U8 : CLKBUF_X1 port map( A => n21202, Z => n21194);
   U9 : CLKBUF_X1 port map( A => n21212, Z => n21195);
   U10 : CLKBUF_X1 port map( A => n21212, Z => n21196);
   U11 : CLKBUF_X1 port map( A => n21212, Z => n21197);
   U12 : CLKBUF_X1 port map( A => n21212, Z => n21198);
   U13 : CLKBUF_X1 port map( A => n21212, Z => n21199);
   U14 : CLKBUF_X1 port map( A => n21211, Z => n21200);
   U15 : CLKBUF_X1 port map( A => n21211, Z => n21201);
   U16 : CLKBUF_X1 port map( A => n21211, Z => n21202);
   U17 : CLKBUF_X1 port map( A => n21211, Z => n21203);
   U18 : CLKBUF_X1 port map( A => n21211, Z => n21204);
   U19 : CLKBUF_X1 port map( A => n21210, Z => n21205);
   U20 : CLKBUF_X1 port map( A => n21210, Z => n21206);
   U21 : CLKBUF_X1 port map( A => n21210, Z => n21207);
   U22 : CLKBUF_X1 port map( A => n21210, Z => n21208);
   U23 : CLKBUF_X1 port map( A => n21210, Z => n21209);
   U24 : CLKBUF_X1 port map( A => n21189, Z => n21210);
   U25 : CLKBUF_X1 port map( A => n21189, Z => n21211);
   U26 : CLKBUF_X1 port map( A => n21190, Z => n21212);
   U27 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n21213);
   U28 : INV_X1 port map( A => n21213, ZN => n21214);
   U29 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , A2 => n22602, ZN => n22631);
   U30 : NOR2_X2 port map( A1 => n21166, A2 => n22802, ZN => n22836);
   U31 : NOR2_X2 port map( A1 => n22765, A2 => n21158, ZN => n22797);
   U32 : NOR2_X2 port map( A1 => n22975, A2 => n22802, ZN => n22835);
   U33 : INV_X2 port map( A => n22092, ZN => n22874);
   U34 : NOR2_X2 port map( A1 => n19293, A2 => n22765, ZN => n22796);
   U35 : NOR2_X2 port map( A1 => n22602, A2 => n22635, ZN => n22637);
   U36 : NOR3_X4 port map( A1 => n21166, A2 => n21159, A3 => n19294, ZN => 
                           n22837);
   U37 : CLKBUF_X1 port map( A => n22083, Z => n22061);
   U38 : INV_X1 port map( A => n22086, ZN => n21982);
   U39 : INV_X1 port map( A => n22958, ZN => n22908);
   U40 : INV_X1 port map( A => n9078, ZN => n1793);
   U41 : INV_X1 port map( A => n22530, ZN => n22941);
   U42 : NAND2_X1 port map( A1 => n21281, A2 => n22874, ZN => n22530);
   U43 : INV_X1 port map( A => n554, ZN => n22568);
   U44 : CLKBUF_X1 port map( A => n22598, Z => n22592);
   U45 : NOR2_X1 port map( A1 => n22920, A2 => n21277, ZN => n1843);
   U46 : NAND2_X1 port map( A1 => n22596, A2 => n22913, ZN => n1834);
   U47 : INV_X1 port map( A => data1_mul_15_port, ZN => n1780);
   U48 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_2_4_port, ZN => 
                           n1791);
   U49 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4295, ZN => n21555);
   U50 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, B2 
                           => n4295, A => n21555, ZN => n1800);
   U51 : INV_X1 port map( A => n14287, ZN => n1797);
   U52 : NAND2_X1 port map( A1 => n4302, A2 => n14286, ZN => n22761);
   U53 : OAI21_X1 port map( B1 => n4302, B2 => n14286, A => n22761, ZN => 
                           n17932);
   U54 : OR2_X1 port map( A1 => n1797, A2 => n17932, ZN => n21185);
   U55 : NOR2_X1 port map( A1 => n7769, A2 => n1800, ZN => n21556);
   U56 : INV_X1 port map( A => n21556, ZN => n1799);
   U57 : XOR2_X1 port map( A => data1_mul_15_port, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => n22762);
   U58 : INV_X1 port map( A => n22762, ZN => n18051);
   U59 : INV_X1 port map( A => DATA2(5), ZN => n22596);
   U60 : INV_X1 port map( A => DATA2(4), ZN => n22913);
   U61 : NAND2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n22920);
   U62 : INV_X1 port map( A => n22920, ZN => n22930);
   U63 : INV_X1 port map( A => DATA2(2), ZN => n22934);
   U64 : INV_X1 port map( A => DATA2(3), ZN => n22933);
   U65 : INV_X1 port map( A => n1834, ZN => n22915);
   U66 : OAI21_X1 port map( B1 => n22934, B2 => n22933, A => n22915, ZN => 
                           n21526);
   U67 : OAI21_X1 port map( B1 => n22930, B2 => n1834, A => n21526, ZN => n1841
                           );
   U68 : INV_X1 port map( A => n1841, ZN => n18195);
   U69 : NOR2_X1 port map( A1 => n22913, A2 => n22933, ZN => n22929);
   U70 : NAND2_X1 port map( A1 => DATA2(2), A2 => n22929, ZN => n22918);
   U71 : NOR2_X1 port map( A1 => n22920, A2 => n22918, ZN => n22335);
   U72 : INV_X1 port map( A => FUNC(0), ZN => n22371);
   U73 : NAND4_X1 port map( A1 => FUNC(2), A2 => FUNC(1), A3 => n22371, A4 => 
                           n22596, ZN => n22336);
   U74 : NOR2_X1 port map( A1 => n22335, A2 => n22336, ZN => n21436);
   U75 : NAND2_X1 port map( A1 => FUNC(3), A2 => n21436, ZN => n1813);
   U76 : NOR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n22917);
   U77 : INV_X1 port map( A => n22929, ZN => n22931);
   U78 : AOI21_X1 port map( B1 => n22917, B2 => n22934, A => n22931, ZN => 
                           n1846);
   U79 : OR2_X1 port map( A1 => n1813, A2 => n1846, ZN => n14273);
   U80 : NAND2_X1 port map( A1 => DATA2(3), A2 => n1834, ZN => n1839);
   U81 : OAI21_X1 port map( B1 => n22934, B2 => n22913, A => n1839, ZN => n1840
                           );
   U82 : INV_X1 port map( A => n1839, ZN => n21215);
   U83 : INV_X1 port map( A => n22917, ZN => n22936);
   U84 : OAI21_X1 port map( B1 => n21215, B2 => n22936, A => n1840, ZN => n1838
                           );
   U85 : INV_X1 port map( A => n1813, ZN => n22126);
   U86 : AND2_X1 port map( A1 => n1838, A2 => n22126, ZN => n17506);
   U87 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n21260);
   U88 : INV_X1 port map( A => FUNC(2), ZN => n21245);
   U89 : NAND2_X1 port map( A1 => n21260, A2 => n21245, ZN => n554);
   U90 : INV_X1 port map( A => n22568, ZN => n22999);
   U91 : NAND2_X1 port map( A1 => n19300, A2 => DATA2_I_4_port, ZN => n21231);
   U92 : OAI21_X1 port map( B1 => n19300, B2 => DATA2_I_4_port, A => n21231, ZN
                           => n1429);
   U93 : NOR2_X1 port map( A1 => n19441, A2 => n22999, ZN => n17537);
   U94 : XNOR2_X1 port map( A => DATA2_I_6_port, B => n22970, ZN => n22880);
   U95 : NOR2_X1 port map( A1 => n22999, A2 => n22966, ZN => n22331);
   U96 : XOR2_X1 port map( A => n19426, B => DATA2_I_5_port, Z => n21674);
   U97 : NAND2_X1 port map( A1 => n19443, A2 => DATA2_I_3_port, ZN => n21221);
   U98 : INV_X1 port map( A => n21221, ZN => n21228);
   U99 : NAND2_X1 port map( A1 => n19442, A2 => DATA2_I_2_port, ZN => n21224);
   U100 : INV_X1 port map( A => n21224, ZN => n21217);
   U101 : NAND2_X1 port map( A1 => n19302, A2 => DATA2_I_1_port, ZN => n21225);
   U102 : INV_X1 port map( A => n21225, ZN => n21216);
   U103 : NOR2_X1 port map( A1 => n19303, A2 => DATA2_I_0_port, ZN => n22329);
   U104 : OAI21_X1 port map( B1 => n19302, B2 => DATA2_I_1_port, A => n21225, 
                           ZN => n22145);
   U105 : NOR2_X1 port map( A1 => n22329, A2 => n22145, ZN => n22141);
   U106 : NOR2_X1 port map( A1 => n21216, A2 => n22141, ZN => n21966);
   U107 : OAI21_X1 port map( B1 => n19442, B2 => DATA2_I_2_port, A => n21224, 
                           ZN => n21965);
   U108 : NOR2_X1 port map( A1 => n21966, A2 => n21965, ZN => n21964);
   U109 : NOR2_X1 port map( A1 => n21217, A2 => n21964, ZN => n21735);
   U110 : OAI21_X1 port map( B1 => n19443, B2 => DATA2_I_3_port, A => n21221, 
                           ZN => n22862);
   U111 : NOR2_X1 port map( A1 => n21735, A2 => n22862, ZN => n21734);
   U112 : NOR2_X1 port map( A1 => n21228, A2 => n21734, ZN => n21702);
   U113 : NOR2_X1 port map( A1 => n21702, A2 => n1429, ZN => n21226);
   U114 : INV_X1 port map( A => n21226, ZN => n21218);
   U115 : NAND2_X1 port map( A1 => n21231, A2 => n21218, ZN => n21670);
   U116 : INV_X1 port map( A => n21670, ZN => n21668);
   U117 : NAND2_X1 port map( A1 => n19299, A2 => DATA2_I_5_port, ZN => n21229);
   U118 : OAI21_X1 port map( B1 => n21674, B2 => n21668, A => n21229, ZN => 
                           n22877);
   U119 : INV_X1 port map( A => n22862, ZN => n21219);
   U120 : INV_X1 port map( A => n21965, ZN => n21969);
   U121 : NAND2_X1 port map( A1 => n19303, A2 => DATA2_I_0_port, ZN => n22146);
   U122 : OAI21_X1 port map( B1 => n22146, B2 => n22145, A => n21225, ZN => 
                           n21968);
   U123 : NAND2_X1 port map( A1 => n21969, A2 => n21968, ZN => n21967);
   U124 : NAND2_X1 port map( A1 => n21224, A2 => n21967, ZN => n22861);
   U125 : NAND2_X1 port map( A1 => n21219, A2 => n22861, ZN => n21220);
   U126 : AND2_X1 port map( A1 => n21221, A2 => n21220, ZN => n21701);
   U127 : OAI21_X1 port map( B1 => n1429, B2 => n21701, A => n21231, ZN => 
                           n21669);
   U128 : INV_X1 port map( A => n21669, ZN => n21667);
   U129 : OAI21_X1 port map( B1 => n21674, B2 => n21667, A => n21229, ZN => 
                           n22875);
   U130 : AOI22_X1 port map( A1 => n22331, A2 => n22877, B1 => n17537, B2 => 
                           n22875, ZN => n21222);
   U131 : OR2_X1 port map( A1 => n22880, A2 => n21222, ZN => n14272);
   U132 : XOR2_X1 port map( A => DATA1(21), B => DATA2_I_21_port, Z => n1809);
   U133 : INV_X1 port map( A => FUNC(3), ZN => n1815);
   U134 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n21243);
   U135 : INV_X1 port map( A => DATA1(20), ZN => n22127);
   U136 : XOR2_X1 port map( A => DATA2_I_20_port, B => n22127, Z => n21250);
   U137 : INV_X1 port map( A => n21250, ZN => n22132);
   U138 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n21242);
   U139 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n22213);
   U140 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n21239);
   U141 : OAI21_X1 port map( B1 => DATA1(17), B2 => DATA2_I_17_port, A => 
                           n21239, ZN => n22212);
   U142 : NOR2_X1 port map( A1 => n22213, A2 => n22212, ZN => n22211);
   U143 : AOI21_X1 port map( B1 => DATA2_I_17_port, B2 => DATA1(17), A => 
                           n22211, ZN => n22189);
   U144 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n21238);
   U145 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => 
                           n21238, ZN => n22194);
   U146 : NOR2_X1 port map( A1 => n22189, A2 => n22194, ZN => n22188);
   U147 : AOI21_X1 port map( B1 => DATA2_I_18_port, B2 => DATA1(18), A => 
                           n22188, ZN => n22175);
   U148 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n21249);
   U149 : OAI21_X1 port map( B1 => n21242, B2 => n22175, A => n21249, ZN => 
                           n22131);
   U150 : NAND2_X1 port map( A1 => n22132, A2 => n22131, ZN => n22130);
   U151 : NAND2_X1 port map( A1 => n21243, A2 => n22130, ZN => n22909);
   U152 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n21236);
   U153 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => 
                           n21236, ZN => n22240);
   U154 : INV_X1 port map( A => DATA1(14), ZN => n22458);
   U155 : XOR2_X1 port map( A => DATA2_I_14_port, B => n22458, Z => n22254);
   U156 : INV_X1 port map( A => n22254, ZN => n22263);
   U157 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n22251);
   U158 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => 
                           n22251, ZN => n22271);
   U159 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n22270);
   U160 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => 
                           n22270, ZN => n22902);
   U161 : NOR2_X1 port map( A1 => n22271, A2 => n22902, ZN => n22238);
   U162 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n21223);
   U163 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n22312
                           );
   U164 : XOR2_X1 port map( A => DATA1(9), B => DATA2_I_9_port, Z => n21598);
   U165 : NAND3_X1 port map( A1 => n19446, A2 => n21598, A3 => DATA2_I_8_port, 
                           ZN => n22309);
   U166 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n22232);
   U167 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n22232, ZN => n22314);
   U168 : AOI21_X1 port map( B1 => n22312, B2 => n22309, A => n22314, ZN => 
                           n22308);
   U169 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => DATA1(10), A => 
                           n22308, ZN => n22298);
   U170 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n22236);
   U171 : OAI21_X1 port map( B1 => n21223, B2 => n22298, A => n22236, ZN => 
                           n22285);
   U172 : NOR2_X1 port map( A1 => n22271, A2 => n22270, ZN => n22237);
   U173 : AOI21_X1 port map( B1 => n22238, B2 => n22285, A => n22237, ZN => 
                           n22253);
   U174 : NAND2_X1 port map( A1 => n22253, A2 => n22251, ZN => n22258);
   U175 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n22263, B2 => n22258, ZN => n22235);
   U176 : NOR2_X1 port map( A1 => n19446, A2 => DATA2_I_8_port, ZN => n21596);
   U177 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => n19446, A => n21596, 
                           ZN => n21635);
   U178 : INV_X1 port map( A => n21598, ZN => n21595);
   U179 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n22236, ZN => n22303);
   U180 : NOR4_X1 port map( A1 => n22314, A2 => n21595, A3 => n22254, A4 => 
                           n22303, ZN => n21235);
   U181 : NAND4_X1 port map( A1 => n21225, A2 => n22146, A3 => n21224, A4 => 
                           n22966, ZN => n21227);
   U182 : OAI21_X1 port map( B1 => n21228, B2 => n21227, A => n21226, ZN => 
                           n21230);
   U183 : OAI221_X1 port map( B1 => n21674, B2 => n21231, C1 => n21674, C2 => 
                           n21230, A => n21229, ZN => n21232);
   U184 : AND2_X1 port map( A1 => n19298, A2 => DATA2_I_6_port, ZN => n21646);
   U185 : AOI21_X1 port map( B1 => n22880, B2 => n21232, A => n21646, ZN => 
                           n21234);
   U186 : NAND2_X1 port map( A1 => DATA2_I_7_port, A2 => n19444, ZN => n21233);
   U187 : OAI21_X1 port map( B1 => DATA2_I_7_port, B2 => n19444, A => n21233, 
                           ZN => n21657);
   U188 : OAI21_X1 port map( B1 => n21234, B2 => n21657, A => n21233, ZN => 
                           n22268);
   U189 : NAND4_X1 port map( A1 => n22238, A2 => n21635, A3 => n21235, A4 => 
                           n22268, ZN => n21237);
   U190 : OAI221_X1 port map( B1 => n22240, B2 => n22235, C1 => n22240, C2 => 
                           n21237, A => n21236, ZN => n21251);
   U191 : NOR2_X1 port map( A1 => n22999, A2 => n21251, ZN => n22910);
   U192 : INV_X1 port map( A => n22910, ZN => n22210);
   U193 : NAND2_X1 port map( A1 => n22568, A2 => n21251, ZN => n22207);
   U194 : INV_X1 port map( A => n21238, ZN => n21241);
   U195 : INV_X1 port map( A => n21239, ZN => n21240);
   U196 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n22209);
   U197 : NOR2_X1 port map( A1 => n22209, A2 => n22212, ZN => n22208);
   U198 : NOR2_X1 port map( A1 => n21240, A2 => n22208, ZN => n22193);
   U199 : NOR2_X1 port map( A1 => n22193, A2 => n22194, ZN => n22192);
   U200 : NOR2_X1 port map( A1 => n21241, A2 => n22192, ZN => n22174);
   U201 : OAI21_X1 port map( B1 => n21242, B2 => n22174, A => n21249, ZN => 
                           n22129);
   U202 : NAND2_X1 port map( A1 => n22132, A2 => n22129, ZN => n22128);
   U203 : NAND2_X1 port map( A1 => n21243, A2 => n22128, ZN => n22911);
   U204 : OAI22_X1 port map( A1 => n22909, A2 => n22210, B1 => n22207, B2 => 
                           n22911, ZN => n21247);
   U205 : NAND2_X1 port map( A1 => FUNC(2), A2 => n21260, ZN => n21244);
   U206 : NOR2_X1 port map( A1 => n1815, A2 => n21244, ZN => n22881);
   U207 : INV_X1 port map( A => n22881, ZN => n22328);
   U208 : INV_X1 port map( A => DATA2(21), ZN => n22579);
   U209 : NAND3_X1 port map( A1 => FUNC(1), A2 => n21245, A3 => n22371, ZN => 
                           n22958);
   U210 : NOR2_X1 port map( A1 => FUNC(3), A2 => n22958, ZN => n22882);
   U211 : INV_X1 port map( A => n22882, ZN => n22221);
   U212 : OAI21_X1 port map( B1 => n22328, B2 => n22579, A => n22221, ZN => 
                           n21246);
   U213 : AOI22_X1 port map( A1 => n21247, A2 => n1809, B1 => n21246, B2 => 
                           DATA1(21), ZN => n21248);
   U214 : INV_X1 port map( A => n21248, ZN => n1779);
   U215 : INV_X1 port map( A => DATA1(2), ZN => n1833);
   U216 : INV_X1 port map( A => DATA1(3), ZN => n1832);
   U217 : INV_X1 port map( A => DATA1(23), ZN => n1825);
   U218 : XNOR2_X1 port map( A => DATA2_I_23_port, B => n1825, ZN => n22100);
   U219 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n22095);
   U220 : OAI21_X1 port map( B1 => DATA1(22), B2 => DATA2_I_22_port, A => 
                           n22095, ZN => n22112);
   U221 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, B1 => 
                           n1809, B2 => n22909, ZN => n22098);
   U222 : INV_X1 port map( A => n22212, ZN => n21253);
   U223 : OAI21_X1 port map( B1 => DATA1(16), B2 => DATA2_I_16_port, A => 
                           n22213, ZN => n21557);
   U224 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => 
                           n21249, ZN => n22179);
   U225 : NOR4_X1 port map( A1 => n22194, A2 => n21250, A3 => n21557, A4 => 
                           n22179, ZN => n21252);
   U226 : NAND4_X1 port map( A1 => n21253, A2 => n1809, A3 => n21252, A4 => 
                           n21251, ZN => n21254);
   U227 : OAI221_X1 port map( B1 => n22112, B2 => n22098, C1 => n22112, C2 => 
                           n21254, A => n22095, ZN => n21255);
   U228 : AOI22_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, B1 => 
                           n22100, B2 => n21255, ZN => n21257);
   U229 : NAND2_X1 port map( A1 => n22568, A2 => n21257, ZN => n22063);
   U230 : INV_X1 port map( A => n22063, ZN => n22079);
   U231 : INV_X1 port map( A => DATA1(27), ZN => n22032);
   U232 : XNOR2_X1 port map( A => DATA2_I_27_port, B => n22032, ZN => n22040);
   U233 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n22078);
   U234 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n21256);
   U235 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => 
                           n21256, ZN => n22068);
   U236 : NOR2_X1 port map( A1 => n22078, A2 => n22068, ZN => n22064);
   U237 : AOI21_X1 port map( B1 => DATA2_I_25_port, B2 => DATA1(25), A => 
                           n22064, ZN => n22052);
   U238 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n21258);
   U239 : OAI21_X1 port map( B1 => DATA1(26), B2 => DATA2_I_26_port, A => 
                           n21258, ZN => n22055);
   U240 : OAI21_X1 port map( B1 => n22052, B2 => n22055, A => n21258, ZN => 
                           n22031);
   U241 : AOI22_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, B1 => 
                           n22040, B2 => n22031, ZN => n21530);
   U242 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n22009);
   U243 : OAI21_X1 port map( B1 => DATA1(28), B2 => DATA2_I_28_port, A => 
                           n22009, ZN => n21529);
   U244 : NOR2_X1 port map( A1 => n21530, A2 => n21529, ZN => n21820);
   U245 : NOR2_X1 port map( A1 => n22999, A2 => n21257, ZN => n22081);
   U246 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n22080);
   U247 : NOR2_X1 port map( A1 => n22080, A2 => n22068, ZN => n22067);
   U248 : AOI21_X1 port map( B1 => DATA2_I_25_port, B2 => DATA1(25), A => 
                           n22067, ZN => n22051);
   U249 : OAI21_X1 port map( B1 => n22051, B2 => n22055, A => n21258, ZN => 
                           n22030);
   U250 : AOI22_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, B1 => 
                           n22040, B2 => n22030, ZN => n21528);
   U251 : NOR2_X1 port map( A1 => n21528, A2 => n21529, ZN => n21822);
   U252 : AOI22_X1 port map( A1 => n22079, A2 => n21820, B1 => n22081, B2 => 
                           n21822, ZN => n21259);
   U253 : INV_X1 port map( A => n21259, ZN => n13930);
   U254 : INV_X1 port map( A => data1_mul_0_port, ZN => n1796);
   U255 : OR4_X1 port map( A1 => DATA1(3), A2 => DATA1(5), A3 => DATA1(4), A4 
                           => DATA1(0), ZN => n13984);
   U256 : INV_X1 port map( A => n9045, ZN => n1781);
   U257 : INV_X1 port map( A => n9048, ZN => n1782);
   U258 : INV_X1 port map( A => n9075, ZN => n1792);
   U259 : INV_X1 port map( A => n9072, ZN => n1790);
   U260 : INV_X1 port map( A => n9069, ZN => n1789);
   U261 : INV_X1 port map( A => n9066, ZN => n1788);
   U262 : INV_X1 port map( A => n9063, ZN => n1787);
   U263 : INV_X1 port map( A => n9060, ZN => n1786);
   U264 : INV_X1 port map( A => n9057, ZN => n1785);
   U265 : INV_X1 port map( A => n9051, ZN => n1783);
   U266 : INV_X1 port map( A => n9054, ZN => n1784);
   U267 : NAND3_X1 port map( A1 => FUNC(2), A2 => n21260, A3 => n1815, ZN => 
                           n7822);
   U268 : NOR4_X1 port map( A1 => DATA2(13), A2 => DATA2(12), A3 => DATA2(11), 
                           A4 => DATA2(6), ZN => n21267);
   U269 : NOR2_X1 port map( A1 => n1834, A2 => DATA2(3), ZN => n21281);
   U270 : NAND2_X1 port map( A1 => n22934, A2 => n21281, ZN => n21440);
   U271 : INV_X1 port map( A => n21440, ZN => n22511);
   U272 : CLKBUF_X1 port map( A => n22511, Z => n21472);
   U273 : NAND2_X1 port map( A1 => n21472, A2 => n22917, ZN => n21981);
   U274 : INV_X1 port map( A => DATA2(15), ZN => n22585);
   U275 : INV_X1 port map( A => DATA2(14), ZN => n22586);
   U276 : INV_X1 port map( A => DATA2(10), ZN => n22589);
   U277 : INV_X1 port map( A => DATA2(8), ZN => n22591);
   U278 : NAND4_X1 port map( A1 => n22585, A2 => n22586, A3 => n22589, A4 => 
                           n22591, ZN => n21261);
   U279 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(7), A3 => n21981, A4 =>
                           n21261, ZN => n21266);
   U280 : OR4_X1 port map( A1 => n19444, A2 => DATA1(11), A3 => n19446, A4 => 
                           n19442, ZN => n21264);
   U281 : NOR4_X1 port map( A1 => DATA1(14), A2 => DATA1(13), A3 => DATA1(12), 
                           A4 => DATA1(9), ZN => n21262);
   U282 : INV_X1 port map( A => DATA1(15), ZN => n22399);
   U283 : INV_X1 port map( A => DATA1(10), ZN => n22451);
   U284 : NAND4_X1 port map( A1 => n19430, A2 => n21262, A3 => n22399, A4 => 
                           n22451, ZN => n21263);
   U285 : NOR4_X1 port map( A1 => n19312, A2 => n19010, A3 => n21264, A4 => 
                           n21263, ZN => n21265);
   U286 : AOI211_X1 port map( C1 => n21267, C2 => n21266, A => n21265, B => 
                           n7822, ZN => n22313);
   U287 : CLKBUF_X1 port map( A => n22313, Z => n22998);
   U288 : INV_X1 port map( A => DATA2(13), ZN => n22587);
   U289 : NOR2_X1 port map( A1 => n22587, A2 => DATA1(13), ZN => n22395);
   U290 : INV_X1 port map( A => n22395, ZN => n22453);
   U291 : NAND2_X1 port map( A1 => n22587, A2 => DATA1(13), ZN => n22457);
   U292 : NAND2_X1 port map( A1 => n22453, A2 => n22457, ZN => n21268);
   U293 : AOI22_X1 port map( A1 => n22998, A2 => n19085, B1 => n22908, B2 => 
                           n21268, ZN => n21269);
   U294 : INV_X1 port map( A => n21269, ZN => n1811);
   U295 : NAND2_X1 port map( A1 => DATA1(29), A2 => n4395, ZN => n21957);
   U296 : OAI21_X1 port map( B1 => DATA1(29), B2 => n4395, A => n21957, ZN => 
                           n8847);
   U297 : INV_X1 port map( A => DATA1(30), ZN => n22502);
   U298 : XOR2_X1 port map( A => DATA2_I_30_port, B => n22502, Z => n21827);
   U299 : INV_X1 port map( A => n21827, ZN => n1801);
   U300 : NAND3_X1 port map( A1 => DATA2(3), A2 => n22915, A3 => n22934, ZN => 
                           n21277);
   U301 : INV_X1 port map( A => n1843, ZN => n17728);
   U302 : INV_X1 port map( A => n21526, ZN => n21270);
   U303 : OAI21_X1 port map( B1 => n22933, B2 => n22920, A => n21270, ZN => 
                           n21533);
   U304 : CLKBUF_X1 port map( A => n21533, Z => n22997);
   U305 : AOI21_X1 port map( B1 => DATA2(1), B2 => DATA2(3), A => n21526, ZN =>
                           n21284);
   U306 : INV_X1 port map( A => n21284, ZN => n22939);
   U307 : NOR3_X1 port map( A1 => n22939, A2 => n21281, A3 => n22917, ZN => 
                           n21293);
   U308 : CLKBUF_X1 port map( A => n21293, Z => n22945);
   U309 : NOR2_X1 port map( A1 => n21440, A2 => n22920, ZN => n21275);
   U310 : INV_X1 port map( A => n21275, ZN => n22017);
   U311 : INV_X1 port map( A => DATA2(0), ZN => n22597);
   U312 : NOR2_X1 port map( A1 => DATA2(1), A2 => n22597, ZN => n22922);
   U313 : NAND2_X1 port map( A1 => n21472, A2 => n22922, ZN => n21802);
   U314 : INV_X1 port map( A => n21802, ZN => n22144);
   U315 : INV_X1 port map( A => DATA2(1), ZN => n22919);
   U316 : OR3_X1 port map( A1 => DATA2(0), A2 => n22919, A3 => n21440, ZN => 
                           n22016);
   U317 : NOR2_X1 port map( A1 => n21165, A2 => n22016, ZN => n21429);
   U318 : NOR2_X1 port map( A1 => n19426, A2 => n21472, ZN => n22150);
   U319 : AOI211_X1 port map( C1 => n22144, C2 => n19446, A => n21429, B => 
                           n22150, ZN => n21271);
   U320 : INV_X1 port map( A => n21981, ZN => n22514);
   U321 : CLKBUF_X1 port map( A => n22514, Z => n22002);
   U322 : NAND2_X1 port map( A1 => DATA1(9), A2 => n22002, ZN => n21396);
   U323 : OAI211_X1 port map( C1 => n22017, C2 => n22970, A => n21271, B => 
                           n21396, ZN => n21292);
   U324 : OAI21_X1 port map( B1 => n22934, B2 => n22919, A => n21281, ZN => 
                           n21274);
   U325 : CLKBUF_X1 port map( A => n21274, Z => n22516);
   U326 : INV_X1 port map( A => n22016, ZN => n21978);
   U327 : NOR2_X1 port map( A1 => n21165, A2 => n22017, ZN => n21708);
   U328 : NOR2_X1 port map( A1 => n19427, A2 => n21472, ZN => n21976);
   U329 : AOI211_X1 port map( C1 => n21978, C2 => n19446, A => n21708, B => 
                           n21976, ZN => n21272);
   U330 : NAND2_X1 port map( A1 => DATA1(9), A2 => n22144, ZN => n21385);
   U331 : OAI211_X1 port map( C1 => n21981, C2 => n22451, A => n21272, B => 
                           n21385, ZN => n21286);
   U332 : AND3_X1 port map( A1 => DATA2(2), A2 => n21281, A3 => n22922, ZN => 
                           n22518);
   U333 : INV_X1 port map( A => DATA1(11), ZN => n22294);
   U334 : NOR2_X1 port map( A1 => n22969, A2 => n22017, ZN => n21428);
   U335 : NOR2_X1 port map( A1 => n21165, A2 => n21472, ZN => n21738);
   U336 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(9), A => n21428, B => 
                           n21738, ZN => n21273);
   U337 : NAND2_X1 port map( A1 => DATA1(10), A2 => n22144, ZN => n21398);
   U338 : OAI211_X1 port map( C1 => n21981, C2 => n22294, A => n21273, B => 
                           n21398, ZN => n21279);
   U339 : INV_X1 port map( A => n21274, ZN => n22083);
   U340 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(0), ZN => n21527);
   U341 : NAND2_X1 port map( A1 => n22061, A2 => n21527, ZN => n22086);
   U342 : AOI222_X1 port map( A1 => n21292, A2 => n22516, B1 => n21286, B2 => 
                           n22518, C1 => n21279, C2 => n21982, ZN => n21791);
   U343 : INV_X1 port map( A => n21791, ZN => n21540);
   U344 : INV_X1 port map( A => DATA1(12), ZN => n22897);
   U345 : CLKBUF_X1 port map( A => n21275, Z => n22047);
   U346 : NOR2_X1 port map( A1 => n22294, A2 => n21802, ZN => n21392);
   U347 : NOR2_X1 port map( A1 => n21472, A2 => n22969, ZN => n21703);
   U348 : AOI211_X1 port map( C1 => n22047, C2 => DATA1(9), A => n21392, B => 
                           n21703, ZN => n21276);
   U349 : NAND2_X1 port map( A1 => DATA1(10), A2 => n21978, ZN => n21384);
   U350 : OAI211_X1 port map( C1 => n21981, C2 => n22897, A => n21276, B => 
                           n21384, ZN => n21283);
   U351 : AOI222_X1 port map( A1 => n21286, A2 => n22516, B1 => n21279, B2 => 
                           n22518, C1 => n21283, C2 => n21982, ZN => n21792);
   U352 : OR2_X1 port map( A1 => n22936, A2 => n21277, ZN => n22948);
   U353 : INV_X1 port map( A => DATA1(13), ZN => n21324);
   U354 : NOR2_X1 port map( A1 => n22897, A2 => n21802, ZN => n21410);
   U355 : NOR2_X1 port map( A1 => n22451, A2 => n22017, ZN => n21400);
   U356 : AOI211_X1 port map( C1 => DATA1(9), C2 => n21440, A => n21410, B => 
                           n21400, ZN => n21278);
   U357 : NAND2_X1 port map( A1 => DATA1(11), A2 => n21978, ZN => n21395);
   U358 : OAI211_X1 port map( C1 => n21981, C2 => n21324, A => n21278, B => 
                           n21395, ZN => n21302);
   U359 : AOI222_X1 port map( A1 => n21279, A2 => n22516, B1 => n21283, B2 => 
                           n22518, C1 => n21302, C2 => n21982, ZN => n21541);
   U360 : AOI21_X1 port map( B1 => n22597, B2 => n21281, A => n22061, ZN => 
                           n21280);
   U361 : INV_X1 port map( A => n21280, ZN => n22943);
   U362 : CLKBUF_X1 port map( A => n22943, Z => n22092);
   U363 : OAI22_X1 port map( A1 => n21792, A2 => n22948, B1 => n21541, B2 => 
                           n22530, ZN => n21289);
   U364 : NOR2_X1 port map( A1 => n21472, A2 => n22451, ZN => n21405);
   U365 : NOR2_X1 port map( A1 => n22294, A2 => n22017, ZN => n21382);
   U366 : AOI211_X1 port map( C1 => n22144, C2 => DATA1(13), A => n21405, B => 
                           n21382, ZN => n21282);
   U367 : NAND2_X1 port map( A1 => DATA1(12), A2 => n21978, ZN => n21389);
   U368 : OAI211_X1 port map( C1 => n21981, C2 => n22458, A => n21282, B => 
                           n21389, ZN => n21301);
   U369 : AOI222_X1 port map( A1 => n21283, A2 => n22516, B1 => n21302, B2 => 
                           n22518, C1 => n21301, C2 => n21982, ZN => n21551);
   U370 : CLKBUF_X1 port map( A => n21284, Z => n22866);
   U371 : NOR2_X1 port map( A1 => n22969, A2 => n21981, ZN => n21383);
   U372 : NAND2_X1 port map( A1 => n22144, A2 => n19444, ZN => n21406);
   U373 : NAND2_X1 port map( A1 => n19299, A2 => n22047, ZN => n21979);
   U374 : OAI211_X1 port map( C1 => n19428, C2 => n21472, A => n21406, B => 
                           n21979, ZN => n21285);
   U375 : AOI211_X1 port map( C1 => n21978, C2 => n19298, A => n21383, B => 
                           n21285, ZN => n21441);
   U376 : INV_X1 port map( A => n21441, ZN => n21287);
   U377 : AOI222_X1 port map( A1 => n21287, A2 => n22516, B1 => n21292, B2 => 
                           n22518, C1 => n21286, C2 => n21982, ZN => n21794);
   U378 : OAI22_X1 port map( A1 => n22874, A2 => n21551, B1 => n22866, B2 => 
                           n21794, ZN => n21288);
   U379 : AOI211_X1 port map( C1 => n22945, C2 => n21540, A => n21289, B => 
                           n21288, ZN => n1803);
   U380 : NOR2_X1 port map( A1 => n22970, A2 => n21802, ZN => n21430);
   U381 : NOR2_X1 port map( A1 => n19426, A2 => n22016, ZN => n21739);
   U382 : NOR2_X1 port map( A1 => n19428, A2 => n22017, ZN => n22149);
   U383 : OAI22_X1 port map( A1 => n21165, A2 => n21981, B1 => n19311, B2 => 
                           n21472, ZN => n21290);
   U384 : NOR4_X1 port map( A1 => n21430, A2 => n21739, A3 => n22149, A4 => 
                           n21290, ZN => n21444);
   U385 : INV_X1 port map( A => n22518, ZN => n22048);
   U386 : OAI22_X1 port map( A1 => n22061, A2 => n21444, B1 => n21441, B2 => 
                           n22048, ZN => n21291);
   U387 : AOI21_X1 port map( B1 => n21982, B2 => n21292, A => n21291, ZN => 
                           n21793);
   U388 : INV_X1 port map( A => n21793, ZN => n21437);
   U389 : OAI22_X1 port map( A1 => n22874, A2 => n21541, B1 => n21792, B2 => 
                           n22530, ZN => n21295);
   U390 : INV_X1 port map( A => n21293, ZN => n22864);
   U391 : OAI22_X1 port map( A1 => n21794, A2 => n22864, B1 => n21791, B2 => 
                           n22948, ZN => n21294);
   U392 : AOI211_X1 port map( C1 => n22939, C2 => n21437, A => n21295, B => 
                           n21294, ZN => n22273);
   U393 : OAI22_X1 port map( A1 => n17728, A2 => n22273, B1 => n22997, B2 => 
                           n1803, ZN => n21296);
   U394 : INV_X1 port map( A => n21296, ZN => n16713);
   U395 : INV_X1 port map( A => n22518, ZN => n21495);
   U396 : NOR2_X1 port map( A1 => n22458, A2 => n22016, ZN => n21322);
   U397 : NAND2_X1 port map( A1 => DATA1(12), A2 => n21440, ZN => n21380);
   U398 : NAND2_X1 port map( A1 => DATA1(13), A2 => n22047, ZN => n21388);
   U399 : OAI211_X1 port map( C1 => n21802, C2 => n22399, A => n21380, B => 
                           n21388, ZN => n21297);
   U400 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(16), A => n21322, B => 
                           n21297, ZN => n21372);
   U401 : NOR2_X1 port map( A1 => n22399, A2 => n22016, ZN => n21318);
   U402 : INV_X1 port map( A => DATA1(16), ZN => n22398);
   U403 : NAND2_X1 port map( A1 => DATA1(13), A2 => n21440, ZN => n21393);
   U404 : NAND2_X1 port map( A1 => DATA1(14), A2 => n22047, ZN => n21412);
   U405 : OAI211_X1 port map( C1 => n21802, C2 => n22398, A => n21393, B => 
                           n21412, ZN => n21298);
   U406 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(17), A => n21318, B => 
                           n21298, ZN => n21374);
   U407 : NOR2_X1 port map( A1 => n21324, A2 => n22016, ZN => n21409);
   U408 : NAND2_X1 port map( A1 => DATA1(11), A2 => n21440, ZN => n21402);
   U409 : NAND2_X1 port map( A1 => DATA1(12), A2 => n22047, ZN => n21394);
   U410 : OAI211_X1 port map( C1 => n21802, C2 => n22458, A => n21402, B => 
                           n21394, ZN => n21299);
   U411 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(15), A => n21409, B => 
                           n21299, ZN => n21304);
   U412 : OAI222_X1 port map( A1 => n21495, A2 => n21372, B1 => n22086, B2 => 
                           n21374, C1 => n21304, C2 => n22083, ZN => n21554);
   U413 : INV_X1 port map( A => n21541, ZN => n21300);
   U414 : AOI22_X1 port map( A1 => n22943, A2 => n21554, B1 => n22939, B2 => 
                           n21300, ZN => n21307);
   U415 : INV_X1 port map( A => n21301, ZN => n21305);
   U416 : OAI222_X1 port map( A1 => n21495, A2 => n21304, B1 => n22086, B2 => 
                           n21372, C1 => n21305, C2 => n22083, ZN => n21543);
   U417 : INV_X1 port map( A => n22948, ZN => n22524);
   U418 : INV_X1 port map( A => n21302, ZN => n21303);
   U419 : OAI222_X1 port map( A1 => n21495, A2 => n21305, B1 => n22086, B2 => 
                           n21304, C1 => n21303, C2 => n22083, ZN => n21544);
   U420 : AOI22_X1 port map( A1 => n22941, A2 => n21543, B1 => n22524, B2 => 
                           n21544, ZN => n21306);
   U421 : OAI211_X1 port map( C1 => n21551, C2 => n22864, A => n21307, B => 
                           n21306, ZN => n1805);
   U422 : NOR2_X1 port map( A1 => n22398, A2 => n21981, ZN => n21310);
   U423 : NAND2_X1 port map( A1 => DATA1(19), A2 => n22047, ZN => n21369);
   U424 : NAND2_X1 port map( A1 => DATA1(17), A2 => n22144, ZN => n21308);
   U425 : OAI211_X1 port map( C1 => n22511, C2 => n22127, A => n21369, B => 
                           n21308, ZN => n21309);
   U426 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(18), A => n21310, B => 
                           n21309, ZN => n21316);
   U427 : INV_X1 port map( A => DATA1(17), ZN => n22205);
   U428 : NOR2_X1 port map( A1 => n22205, A2 => n22016, ZN => n21358);
   U429 : NAND2_X1 port map( A1 => n21440, A2 => DATA1(19), ZN => n21454);
   U430 : NAND2_X1 port map( A1 => DATA1(18), A2 => n22047, ZN => n21365);
   U431 : OAI211_X1 port map( C1 => n21802, C2 => n22398, A => n21454, B => 
                           n21365, ZN => n21311);
   U432 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(15), A => n21358, B => 
                           n21311, ZN => n21321);
   U433 : INV_X1 port map( A => DATA1(21), ZN => n21471);
   U434 : NOR2_X1 port map( A1 => n21472, A2 => n21471, ZN => n21313);
   U435 : NOR2_X1 port map( A1 => n22127, A2 => n22017, ZN => n21457);
   U436 : AND2_X1 port map( A1 => DATA1(19), A2 => n21978, ZN => n21364);
   U437 : INV_X1 port map( A => DATA1(18), ZN => n22191);
   U438 : OAI22_X1 port map( A1 => n22191, A2 => n21802, B1 => n22205, B2 => 
                           n21981, ZN => n21312);
   U439 : NOR4_X1 port map( A1 => n21313, A2 => n21457, A3 => n21364, A4 => 
                           n21312, ZN => n21331);
   U440 : OAI222_X1 port map( A1 => n21495, A2 => n21316, B1 => n22086, B2 => 
                           n21321, C1 => n21331, C2 => n22083, ZN => n21558);
   U441 : INV_X1 port map( A => n21558, ZN => n21565);
   U442 : NOR2_X1 port map( A1 => n21472, A2 => n22191, ZN => n21367);
   U443 : NOR2_X1 port map( A1 => n22205, A2 => n22017, ZN => n21360);
   U444 : NOR2_X1 port map( A1 => n22398, A2 => n22016, ZN => n21355);
   U445 : OAI22_X1 port map( A1 => n22399, A2 => n21802, B1 => n22458, B2 => 
                           n21981, ZN => n21314);
   U446 : NOR4_X1 port map( A1 => n21367, A2 => n21360, A3 => n21355, A4 => 
                           n21314, ZN => n21325);
   U447 : OAI222_X1 port map( A1 => n21495, A2 => n21321, B1 => n22086, B2 => 
                           n21325, C1 => n21316, C2 => n22083, ZN => n21559);
   U448 : NOR2_X1 port map( A1 => n21471, A2 => n22017, ZN => n21468);
   U449 : NOR2_X1 port map( A1 => n22127, A2 => n22016, ZN => n21368);
   U450 : AOI211_X1 port map( C1 => DATA1(22), C2 => n21440, A => n21468, B => 
                           n21368, ZN => n21315);
   U451 : NAND2_X1 port map( A1 => DATA1(19), A2 => n22144, ZN => n21361);
   U452 : OAI211_X1 port map( C1 => n21981, C2 => n22191, A => n21315, B => 
                           n21361, ZN => n21421);
   U453 : INV_X1 port map( A => n21982, ZN => n22520);
   U454 : OAI22_X1 port map( A1 => n21316, A2 => n22520, B1 => n21331, B2 => 
                           n22048, ZN => n21317);
   U455 : AOI21_X1 port map( B1 => n22516, B2 => n21421, A => n21317, ZN => 
                           n21498);
   U456 : INV_X1 port map( A => n21498, ZN => n22942);
   U457 : AOI22_X1 port map( A1 => n22524, A2 => n21559, B1 => n22939, B2 => 
                           n22942, ZN => n21328);
   U458 : NOR2_X1 port map( A1 => n21472, A2 => n22205, ZN => n21363);
   U459 : AOI211_X1 port map( C1 => n22047, C2 => DATA1(16), A => n21363, B => 
                           n21318, ZN => n21320);
   U460 : NAND2_X1 port map( A1 => DATA1(13), A2 => n22002, ZN => n21319);
   U461 : OAI211_X1 port map( C1 => n21802, C2 => n22458, A => n21320, B => 
                           n21319, ZN => n21449);
   U462 : INV_X1 port map( A => n21449, ZN => n21326);
   U463 : OAI222_X1 port map( A1 => n21495, A2 => n21325, B1 => n22086, B2 => 
                           n21326, C1 => n21321, C2 => n22083, ZN => n21568);
   U464 : NOR2_X1 port map( A1 => n21472, A2 => n22398, ZN => n21359);
   U465 : AOI211_X1 port map( C1 => n22002, C2 => DATA1(12), A => n21359, B => 
                           n21322, ZN => n21323);
   U466 : NAND2_X1 port map( A1 => DATA1(15), A2 => n22047, ZN => n21353);
   U467 : OAI211_X1 port map( C1 => n21802, C2 => n21324, A => n21323, B => 
                           n21353, ZN => n21448);
   U468 : INV_X1 port map( A => n21448, ZN => n21416);
   U469 : OAI222_X1 port map( A1 => n21495, A2 => n21326, B1 => n22086, B2 => 
                           n21416, C1 => n21325, C2 => n22083, ZN => n21573);
   U470 : AOI22_X1 port map( A1 => n22941, A2 => n21568, B1 => n22943, B2 => 
                           n21573, ZN => n21327);
   U471 : OAI211_X1 port map( C1 => n21565, C2 => n22864, A => n21328, B => 
                           n21327, ZN => n1828);
   U472 : NAND2_X1 port map( A1 => DATA1(23), A2 => n21440, ZN => n21503);
   U473 : INV_X1 port map( A => n21503, ZN => n21329);
   U474 : INV_X1 port map( A => DATA1(22), ZN => n22475);
   U475 : NOR2_X1 port map( A1 => n22475, A2 => n22017, ZN => n21474);
   U476 : AOI211_X1 port map( C1 => n22144, C2 => DATA1(20), A => n21329, B => 
                           n21474, ZN => n21330);
   U477 : NAND2_X1 port map( A1 => DATA1(19), A2 => n22002, ZN => n21356);
   U478 : OAI211_X1 port map( C1 => n22016, C2 => n21471, A => n21330, B => 
                           n21356, ZN => n21422);
   U479 : INV_X1 port map( A => n21331, ZN => n21332);
   U480 : AOI222_X1 port map( A1 => n21422, A2 => n22516, B1 => n21421, B2 => 
                           n22518, C1 => n21332, C2 => n21982, ZN => n21563);
   U481 : INV_X1 port map( A => n21563, ZN => n22940);
   U482 : AOI22_X1 port map( A1 => n22524, A2 => n21558, B1 => n22939, B2 => 
                           n22940, ZN => n21334);
   U483 : AOI22_X1 port map( A1 => n22941, A2 => n21559, B1 => n22943, B2 => 
                           n21568, ZN => n21333);
   U484 : OAI211_X1 port map( C1 => n21498, C2 => n22864, A => n21334, B => 
                           n21333, ZN => n14003);
   U485 : NOR2_X1 port map( A1 => n22475, A2 => n21981, ZN => n21336);
   U486 : INV_X1 port map( A => DATA1(26), ZN => n22489);
   U487 : NAND2_X1 port map( A1 => DATA1(25), A2 => n22047, ZN => n21771);
   U488 : NAND2_X1 port map( A1 => DATA1(23), A2 => n22144, ZN => n21465);
   U489 : OAI211_X1 port map( C1 => n22511, C2 => n22489, A => n21771, B => 
                           n21465, ZN => n21335);
   U490 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(24), A => n21336, B => 
                           n21335, ZN => n21350);
   U491 : AOI22_X1 port map( A1 => DATA1(22), A2 => n22144, B1 => DATA1(21), B2
                           => n22002, ZN => n21338);
   U492 : NAND2_X1 port map( A1 => DATA1(24), A2 => n22047, ZN => n21337);
   U493 : NAND2_X1 port map( A1 => DATA1(23), A2 => n21978, ZN => n21469);
   U494 : NAND2_X1 port map( A1 => DATA1(25), A2 => n21440, ZN => n21780);
   U495 : NAND4_X1 port map( A1 => n21338, A2 => n21337, A3 => n21469, A4 => 
                           n21780, ZN => n21348);
   U496 : INV_X1 port map( A => n21348, ZN => n21340);
   U497 : NOR2_X1 port map( A1 => n1825, A2 => n21981, ZN => n21458);
   U498 : INV_X1 port map( A => DATA1(24), ZN => n22483);
   U499 : NAND2_X1 port map( A1 => DATA1(25), A2 => n21978, ZN => n21504);
   U500 : NAND2_X1 port map( A1 => DATA1(27), A2 => n21440, ZN => n21803);
   U501 : OAI211_X1 port map( C1 => n21802, C2 => n22483, A => n21504, B => 
                           n21803, ZN => n21339);
   U502 : AOI211_X1 port map( C1 => n22047, C2 => DATA1(26), A => n21458, B => 
                           n21339, ZN => n21343);
   U503 : OAI222_X1 port map( A1 => n21495, A2 => n21350, B1 => n22086, B2 => 
                           n21340, C1 => n21343, C2 => n22083, ZN => n22872);
   U504 : INV_X1 port map( A => DATA1(25), ZN => n22065);
   U505 : NOR2_X1 port map( A1 => n22065, A2 => n21802, ZN => n21476);
   U506 : INV_X1 port map( A => DATA1(28), ZN => n22495);
   U507 : NAND2_X1 port map( A1 => DATA1(27), A2 => n22047, ZN => n21799);
   U508 : NAND2_X1 port map( A1 => DATA1(24), A2 => n22002, ZN => n21466);
   U509 : OAI211_X1 port map( C1 => n22511, C2 => n22495, A => n21799, B => 
                           n21466, ZN => n21341);
   U510 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(26), A => n21476, B => 
                           n21341, ZN => n22085);
   U511 : NOR2_X1 port map( A1 => n22489, A2 => n21802, ZN => n21502);
   U512 : INV_X1 port map( A => DATA1(29), ZN => n22001);
   U513 : NAND2_X1 port map( A1 => DATA1(27), A2 => n21978, ZN => n21781);
   U514 : NAND2_X1 port map( A1 => DATA1(25), A2 => n22002, ZN => n21470);
   U515 : OAI211_X1 port map( C1 => n22511, C2 => n22001, A => n21781, B => 
                           n21470, ZN => n21342);
   U516 : AOI211_X1 port map( C1 => n22047, C2 => DATA1(28), A => n21502, B => 
                           n21342, ZN => n22087);
   U517 : OAI222_X1 port map( A1 => n22520, A2 => n21343, B1 => n22048, B2 => 
                           n22085, C1 => n22087, C2 => n22083, ZN => n22114);
   U518 : INV_X1 port map( A => n22114, ZN => n22865);
   U519 : INV_X1 port map( A => n21343, ZN => n21345);
   U520 : OAI22_X1 port map( A1 => n22061, A2 => n22085, B1 => n21350, B2 => 
                           n22520, ZN => n21344);
   U521 : AOI21_X1 port map( B1 => n22518, B2 => n21345, A => n21344, ZN => 
                           n22868);
   U522 : OAI22_X1 port map( A1 => n22865, A2 => n22866, B1 => n22868, B2 => 
                           n22864, ZN => n21352);
   U523 : NOR2_X1 port map( A1 => n1825, A2 => n22017, ZN => n21475);
   U524 : NOR2_X1 port map( A1 => n22127, A2 => n21981, ZN => n21346);
   U525 : AOI211_X1 port map( C1 => n22144, C2 => DATA1(21), A => n21475, B => 
                           n21346, ZN => n21347);
   U526 : NAND2_X1 port map( A1 => DATA1(24), A2 => n21440, ZN => n21772);
   U527 : OAI211_X1 port map( C1 => n22016, C2 => n22475, A => n21347, B => 
                           n21772, ZN => n21423);
   U528 : AOI222_X1 port map( A1 => n21348, A2 => n22516, B1 => n21423, B2 => 
                           n22518, C1 => n21422, C2 => n21982, ZN => n21564);
   U529 : AOI22_X1 port map( A1 => n21982, A2 => n21423, B1 => n22518, B2 => 
                           n21348, ZN => n21349);
   U530 : OAI21_X1 port map( B1 => n22061, B2 => n21350, A => n21349, ZN => 
                           n22938);
   U531 : INV_X1 port map( A => n22938, ZN => n22869);
   U532 : OAI22_X1 port map( A1 => n22874, A2 => n21564, B1 => n22869, B2 => 
                           n22530, ZN => n21351);
   U533 : AOI211_X1 port map( C1 => n22524, C2 => n22872, A => n21352, B => 
                           n21351, ZN => n1816);
   U534 : NAND2_X1 port map( A1 => DATA1(14), A2 => n21440, ZN => n21387);
   U535 : OAI211_X1 port map( C1 => n21802, C2 => n22205, A => n21387, B => 
                           n21353, ZN => n21354);
   U536 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(18), A => n21355, B => 
                           n21354, ZN => n21373);
   U537 : NAND2_X1 port map( A1 => DATA1(15), A2 => n21440, ZN => n21411);
   U538 : OAI211_X1 port map( C1 => n22017, C2 => n22398, A => n21356, B => 
                           n21411, ZN => n21357);
   U539 : AOI211_X1 port map( C1 => n22144, C2 => DATA1(18), A => n21358, B => 
                           n21357, ZN => n21375);
   U540 : OAI222_X1 port map( A1 => n21495, A2 => n21373, B1 => n22086, B2 => 
                           n21375, C1 => n21374, C2 => n22083, ZN => n21534);
   U541 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(18), A => n21360, B => 
                           n21359, ZN => n21362);
   U542 : OAI211_X1 port map( C1 => n21981, C2 => n22127, A => n21362, B => 
                           n21361, ZN => n21376);
   U543 : AOI211_X1 port map( C1 => n22002, C2 => DATA1(21), A => n21364, B => 
                           n21363, ZN => n21366);
   U544 : OAI211_X1 port map( C1 => n21802, C2 => n22127, A => n21366, B => 
                           n21365, ZN => n21452);
   U545 : AOI211_X1 port map( C1 => n22144, C2 => DATA1(21), A => n21368, B => 
                           n21367, ZN => n21370);
   U546 : OAI211_X1 port map( C1 => n21981, C2 => n22475, A => n21370, B => 
                           n21369, ZN => n21453);
   U547 : AOI222_X1 port map( A1 => n21376, A2 => n22516, B1 => n21452, B2 => 
                           n22518, C1 => n21453, C2 => n21982, ZN => n21770);
   U548 : OAI22_X1 port map( A1 => n22061, A2 => n21373, B1 => n21375, B2 => 
                           n22048, ZN => n21371);
   U549 : AOI21_X1 port map( B1 => n21982, B2 => n21376, A => n21371, ZN => 
                           n21488);
   U550 : OAI22_X1 port map( A1 => n22874, A2 => n21770, B1 => n21488, B2 => 
                           n22948, ZN => n21379);
   U551 : OAI222_X1 port map( A1 => n21495, A2 => n21374, B1 => n22086, B2 => 
                           n21373, C1 => n21372, C2 => n22083, ZN => n21535);
   U552 : INV_X1 port map( A => n21535, ZN => n21549);
   U553 : INV_X1 port map( A => n21375, ZN => n21377);
   U554 : AOI222_X1 port map( A1 => n21377, A2 => n22516, B1 => n21376, B2 => 
                           n22518, C1 => n21452, C2 => n21982, ZN => n21487);
   U555 : OAI22_X1 port map( A1 => n22866, A2 => n21549, B1 => n21487, B2 => 
                           n22530, ZN => n21378);
   U556 : AOI211_X1 port map( C1 => n22945, C2 => n21534, A => n21379, B => 
                           n21378, ZN => n14407);
   U557 : INV_X1 port map( A => n21380, ZN => n21381);
   U558 : NOR3_X1 port map( A1 => n21383, A2 => n21382, A3 => n21381, ZN => 
                           n21386);
   U559 : NAND3_X1 port map( A1 => n21386, A2 => n21385, A3 => n21384, ZN => 
                           n21408);
   U560 : NAND2_X1 port map( A1 => DATA1(10), A2 => n22002, ZN => n21390);
   U561 : NAND4_X1 port map( A1 => n21390, A2 => n21389, A3 => n21388, A4 => 
                           n21387, ZN => n21391);
   U562 : NOR2_X1 port map( A1 => n21392, A2 => n21391, ZN => n21417);
   U563 : AND4_X1 port map( A1 => n21396, A2 => n21395, A3 => n21394, A4 => 
                           n21393, ZN => n21397);
   U564 : NAND2_X1 port map( A1 => n21398, A2 => n21397, ZN => n21404);
   U565 : INV_X1 port map( A => n21404, ZN => n21415);
   U566 : OAI22_X1 port map( A1 => n22061, A2 => n21417, B1 => n21415, B2 => 
                           n22048, ZN => n21399);
   U567 : AOI21_X1 port map( B1 => n21982, B2 => n21408, A => n21399, ZN => 
                           n21716);
   U568 : NOR2_X1 port map( A1 => n22969, A2 => n21802, ZN => n21401);
   U569 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(9), A => n21401, B => 
                           n21400, ZN => n21403);
   U570 : OAI211_X1 port map( C1 => n21165, C2 => n21981, A => n21403, B => 
                           n21402, ZN => n21433);
   U571 : AOI222_X1 port map( A1 => n21404, A2 => n22516, B1 => n21408, B2 => 
                           n22518, C1 => n21433, C2 => n21982, ZN => n21744);
   U572 : INV_X1 port map( A => n21744, ZN => n21712);
   U573 : INV_X1 port map( A => DATA1(9), ZN => n21432);
   U574 : NOR2_X1 port map( A1 => n19427, A2 => n21981, ZN => n21439);
   U575 : AOI211_X1 port map( C1 => n21978, C2 => n19446, A => n21439, B => 
                           n21405, ZN => n21407);
   U576 : OAI211_X1 port map( C1 => n22017, C2 => n21432, A => n21407, B => 
                           n21406, ZN => n21709);
   U577 : AOI222_X1 port map( A1 => n21408, A2 => n22516, B1 => n21433, B2 => 
                           n22518, C1 => n21709, C2 => n21982, ZN => n21984);
   U578 : INV_X1 port map( A => n21984, ZN => n21713);
   U579 : AOI22_X1 port map( A1 => n22941, A2 => n21712, B1 => n22943, B2 => 
                           n21713, ZN => n21420);
   U580 : NOR2_X1 port map( A1 => n21410, A2 => n21409, ZN => n21414);
   U581 : NAND2_X1 port map( A1 => DATA1(11), A2 => n22002, ZN => n21413);
   U582 : NAND4_X1 port map( A1 => n21414, A2 => n21413, A3 => n21412, A4 => 
                           n21411, ZN => n21447);
   U583 : INV_X1 port map( A => n21447, ZN => n21418);
   U584 : OAI222_X1 port map( A1 => n21495, A2 => n21417, B1 => n22086, B2 => 
                           n21415, C1 => n21418, C2 => n22083, ZN => n21578);
   U585 : OAI222_X1 port map( A1 => n21495, A2 => n21418, B1 => n22086, B2 => 
                           n21417, C1 => n21416, C2 => n22083, ZN => n21571);
   U586 : AOI22_X1 port map( A1 => n22945, A2 => n21578, B1 => n22939, B2 => 
                           n21571, ZN => n21419);
   U587 : OAI211_X1 port map( C1 => n21716, C2 => n22948, A => n21420, B => 
                           n21419, ZN => n1808);
   U588 : AOI222_X1 port map( A1 => n21423, A2 => n22516, B1 => n21422, B2 => 
                           n22518, C1 => n21421, C2 => n21982, ZN => n22949);
   U589 : INV_X1 port map( A => n22868, ZN => n22122);
   U590 : AOI22_X1 port map( A1 => n22945, A2 => n22872, B1 => n22939, B2 => 
                           n22122, ZN => n21425);
   U591 : INV_X1 port map( A => n21564, ZN => n22944);
   U592 : AOI22_X1 port map( A1 => n22941, A2 => n22944, B1 => n22524, B2 => 
                           n22938, ZN => n21424);
   U593 : OAI211_X1 port map( C1 => n22874, C2 => n22949, A => n21425, B => 
                           n21424, ZN => n1817);
   U594 : AOI22_X1 port map( A1 => n22524, A2 => n22944, B1 => n22945, B2 => 
                           n22938, ZN => n21427);
   U595 : AOI22_X1 port map( A1 => n22943, A2 => n22940, B1 => n22939, B2 => 
                           n22872, ZN => n21426);
   U596 : OAI211_X1 port map( C1 => n22949, C2 => n22530, A => n21427, B => 
                           n21426, ZN => n1821);
   U597 : NOR3_X1 port map( A1 => n21430, A2 => n21429, A3 => n21428, ZN => 
                           n21431);
   U598 : NAND2_X1 port map( A1 => n19299, A2 => n22002, ZN => n21442);
   U599 : OAI211_X1 port map( C1 => n22511, C2 => n21432, A => n21431, B => 
                           n21442, ZN => n21743);
   U600 : AOI222_X1 port map( A1 => n21433, A2 => n22516, B1 => n21709, B2 => 
                           n22518, C1 => n21743, C2 => n21982, ZN => n22155);
   U601 : OAI22_X1 port map( A1 => n22874, A2 => n22155, B1 => n21744, B2 => 
                           n22948, ZN => n21435);
   U602 : OAI22_X1 port map( A1 => n21716, A2 => n22864, B1 => n21984, B2 => 
                           n22530, ZN => n21434);
   U603 : AOI211_X1 port map( C1 => n22939, C2 => n21578, A => n21435, B => 
                           n21434, ZN => n1807);
   U604 : NAND2_X1 port map( A1 => n21436, A2 => n1815, ZN => n1814);
   U605 : AOI22_X1 port map( A1 => n22524, A2 => n21437, B1 => n22943, B2 => 
                           n21540, ZN => n21446);
   U606 : NAND2_X1 port map( A1 => n19443, A2 => n22047, ZN => n22509);
   U607 : NAND2_X1 port map( A1 => n22144, A2 => n22986, ZN => n21706);
   U608 : OAI211_X1 port map( C1 => n19428, C2 => n22016, A => n22509, B => 
                           n21706, ZN => n21438);
   U609 : AOI211_X1 port map( C1 => n19442, C2 => n21440, A => n21439, B => 
                           n21438, ZN => n21494);
   U610 : OAI222_X1 port map( A1 => n22048, A2 => n21444, B1 => n22086, B2 => 
                           n21441, C1 => n21494, C2 => n22083, ZN => n21797);
   U611 : NOR2_X1 port map( A1 => n19428, A2 => n21802, ZN => n21740);
   U612 : NAND2_X1 port map( A1 => n19443, A2 => n21978, ZN => n22152);
   U613 : OAI211_X1 port map( C1 => n22511, C2 => n19430, A => n21442, B => 
                           n22152, ZN => n21443);
   U614 : AOI211_X1 port map( C1 => n22047, C2 => n19442, A => n21740, B => 
                           n21443, ZN => n21664);
   U615 : OAI222_X1 port map( A1 => n21495, A2 => n21494, B1 => n22520, B2 => 
                           n21444, C1 => n21664, C2 => n22083, ZN => n21652);
   U616 : AOI22_X1 port map( A1 => n22945, A2 => n21797, B1 => n21652, B2 => 
                           n22939, ZN => n21445);
   U617 : OAI211_X1 port map( C1 => n21794, C2 => n22530, A => n21446, B => 
                           n21445, ZN => n1804);
   U618 : AOI222_X1 port map( A1 => n21449, A2 => n22516, B1 => n21448, B2 => 
                           n22518, C1 => n21447, C2 => n21982, ZN => n21574);
   U619 : AOI22_X1 port map( A1 => n22943, A2 => n21571, B1 => n22939, B2 => 
                           n21559, ZN => n21451);
   U620 : AOI22_X1 port map( A1 => n22524, A2 => n21573, B1 => n22945, B2 => 
                           n21568, ZN => n21450);
   U621 : OAI211_X1 port map( C1 => n21574, C2 => n22530, A => n21451, B => 
                           n21450, ZN => n1830);
   U622 : INV_X1 port map( A => n21487, ZN => n21767);
   U623 : INV_X1 port map( A => n21452, ZN => n21459);
   U624 : INV_X1 port map( A => n21453, ZN => n21481);
   U625 : INV_X1 port map( A => n21454, ZN => n21456);
   U626 : OAI22_X1 port map( A1 => n22475, A2 => n21802, B1 => n21471, B2 => 
                           n22016, ZN => n21455);
   U627 : NOR4_X1 port map( A1 => n21458, A2 => n21457, A3 => n21456, A4 => 
                           n21455, ZN => n21480);
   U628 : OAI222_X1 port map( A1 => n21459, A2 => n22061, B1 => n21481, B2 => 
                           n22048, C1 => n21480, C2 => n22520, ZN => n21766);
   U629 : AOI22_X1 port map( A1 => n22524, A2 => n21767, B1 => n22943, B2 => 
                           n21766, ZN => n21461);
   U630 : INV_X1 port map( A => n21488, ZN => n21762);
   U631 : AOI22_X1 port map( A1 => n22945, A2 => n21762, B1 => n22939, B2 => 
                           n21534, ZN => n21460);
   U632 : OAI211_X1 port map( C1 => n21770, C2 => n22530, A => n21461, B => 
                           n21460, ZN => n1826);
   U633 : INV_X1 port map( A => n21578, ZN => n21462);
   U634 : OAI22_X1 port map( A1 => n21462, A2 => n22948, B1 => n21716, B2 => 
                           n22530, ZN => n21464);
   U635 : OAI22_X1 port map( A1 => n22874, A2 => n21744, B1 => n22866, B2 => 
                           n21574, ZN => n21463);
   U636 : AOI211_X1 port map( C1 => n22945, C2 => n21571, A => n21464, B => 
                           n21463, ZN => n1810);
   U637 : OAI211_X1 port map( C1 => n21472, C2 => n22127, A => n21466, B => 
                           n21465, ZN => n21467);
   U638 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(22), A => n21468, B => 
                           n21467, ZN => n21479);
   U639 : OAI211_X1 port map( C1 => n21472, C2 => n21471, A => n21470, B => 
                           n21469, ZN => n21473);
   U640 : AOI211_X1 port map( C1 => n22144, C2 => DATA1(24), A => n21474, B => 
                           n21473, ZN => n21506);
   U641 : OAI222_X1 port map( A1 => n21495, A2 => n21479, B1 => n22086, B2 => 
                           n21506, C1 => n21480, C2 => n22061, ZN => n21784);
   U642 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(24), A => n21476, B => 
                           n21475, ZN => n21477);
   U643 : NAND2_X1 port map( A1 => DATA1(26), A2 => n22002, ZN => n22043);
   U644 : OAI211_X1 port map( C1 => n22511, C2 => n22475, A => n21477, B => 
                           n22043, ZN => n21478);
   U645 : INV_X1 port map( A => n21478, ZN => n21774);
   U646 : OAI222_X1 port map( A1 => n21479, A2 => n22061, B1 => n21506, B2 => 
                           n22048, C1 => n21774, C2 => n22520, ZN => n21815);
   U647 : INV_X1 port map( A => n21815, ZN => n21787);
   U648 : OAI222_X1 port map( A1 => n21481, A2 => n22061, B1 => n21480, B2 => 
                           n22048, C1 => n21479, C2 => n22520, ZN => n21775);
   U649 : INV_X1 port map( A => n21775, ZN => n21507);
   U650 : OAI22_X1 port map( A1 => n22874, A2 => n21787, B1 => n21507, B2 => 
                           n22948, ZN => n21483);
   U651 : INV_X1 port map( A => n21766, ZN => n21765);
   U652 : OAI22_X1 port map( A1 => n22866, A2 => n21770, B1 => n21765, B2 => 
                           n22864, ZN => n21482);
   U653 : AOI211_X1 port map( C1 => n22941, C2 => n21784, A => n21483, B => 
                           n21482, ZN => n1823);
   U654 : OAI21_X2 port map( B1 => DATA2(1), B2 => n1834, A => n21526, ZN => 
                           n1836);
   U655 : INV_X1 port map( A => n21534, ZN => n21486);
   U656 : OAI22_X1 port map( A1 => n22874, A2 => n21488, B1 => n21486, B2 => 
                           n22530, ZN => n21485);
   U657 : INV_X1 port map( A => n21543, ZN => n21550);
   U658 : INV_X1 port map( A => n21554, ZN => n21489);
   U659 : OAI22_X1 port map( A1 => n22866, A2 => n21550, B1 => n21489, B2 => 
                           n22864, ZN => n21484);
   U660 : AOI211_X1 port map( C1 => n22524, C2 => n21535, A => n21485, B => 
                           n21484, ZN => n1831);
   U661 : INV_X1 port map( A => n1836, ZN => n13151);
   U662 : NOR3_X4 port map( A1 => n13151, A2 => n21527, A3 => n22933, ZN => 
                           n1894);
   U663 : INV_X1 port map( A => n1894, ZN => n1837);
   U664 : OAI22_X1 port map( A1 => n22874, A2 => n21487, B1 => n21486, B2 => 
                           n22948, ZN => n21491);
   U665 : OAI22_X1 port map( A1 => n22866, A2 => n21489, B1 => n21488, B2 => 
                           n22530, ZN => n21490);
   U666 : AOI211_X1 port map( C1 => n22945, C2 => n21535, A => n21491, B => 
                           n21490, ZN => n21838);
   U667 : OAI22_X1 port map( A1 => n1836, A2 => n1831, B1 => n1837, B2 => 
                           n21838, ZN => n21492);
   U668 : INV_X1 port map( A => n21492, ZN => n1829);
   U669 : INV_X1 port map( A => n21652, ZN => n21590);
   U670 : OAI22_X1 port map( A1 => n21590, A2 => n22864, B1 => n21793, B2 => 
                           n22530, ZN => n21497);
   U671 : NOR2_X1 port map( A1 => n19309, A2 => n22016, ZN => n22513);
   U672 : NAND2_X1 port map( A1 => n19300, A2 => n22002, ZN => n21705);
   U673 : NAND2_X1 port map( A1 => n19443, A2 => n22144, ZN => n21975);
   U674 : OAI211_X1 port map( C1 => n19429, C2 => n22511, A => n21705, B => 
                           n21975, ZN => n21493);
   U675 : AOI211_X1 port map( C1 => n22047, C2 => n19302, A => n22513, B => 
                           n21493, ZN => n21696);
   U676 : OAI222_X1 port map( A1 => n21495, A2 => n21664, B1 => n22520, B2 => 
                           n21494, C1 => n21696, C2 => n22083, ZN => n22887);
   U677 : INV_X1 port map( A => n22887, ZN => n21588);
   U678 : OAI22_X1 port map( A1 => n22874, A2 => n21794, B1 => n21588, B2 => 
                           n22866, ZN => n21496);
   U679 : AOI211_X1 port map( C1 => n22524, C2 => n21797, A => n21497, B => 
                           n21496, ZN => n12526);
   U680 : OR3_X1 port map( A1 => n22997, A2 => n1814, A3 => n12526, ZN => 
                           n14146);
   U681 : CLKBUF_X1 port map( A => n22941, Z => n22873);
   U682 : OAI22_X1 port map( A1 => n21498, A2 => n22948, B1 => n21563, B2 => 
                           n22864, ZN => n21501);
   U683 : INV_X1 port map( A => n21559, ZN => n21499);
   U684 : OAI22_X1 port map( A1 => n22874, A2 => n21499, B1 => n22866, B2 => 
                           n22949, ZN => n21500);
   U685 : AOI211_X1 port map( C1 => n22873, C2 => n21558, A => n21501, B => 
                           n21500, ZN => n1824);
   U686 : AOI21_X1 port map( B1 => n22047, B2 => DATA1(24), A => n21502, ZN => 
                           n21505);
   U687 : NAND2_X1 port map( A1 => DATA1(27), A2 => n22002, ZN => n22025);
   U688 : AND4_X1 port map( A1 => n21505, A2 => n22025, A3 => n21504, A4 => 
                           n21503, ZN => n21783);
   U689 : OAI222_X1 port map( A1 => n21506, A2 => n22061, B1 => n21774, B2 => 
                           n22048, C1 => n21783, C2 => n22520, ZN => n21808);
   U690 : INV_X1 port map( A => n21808, ZN => n21819);
   U691 : INV_X1 port map( A => n21784, ZN => n21778);
   U692 : OAI22_X1 port map( A1 => n22874, A2 => n21819, B1 => n21778, B2 => 
                           n22948, ZN => n21509);
   U693 : OAI22_X1 port map( A1 => n22866, A2 => n21765, B1 => n21507, B2 => 
                           n22864, ZN => n21508);
   U694 : AOI211_X1 port map( C1 => n22941, C2 => n21815, A => n21509, B => 
                           n21508, ZN => n1819);
   U695 : OAI211_X1 port map( C1 => n19356, C2 => n18953, A => n19003, B => 
                           n21168, ZN => n21510);
   U696 : INV_X1 port map( A => n21510, ZN => n21847);
   U697 : OAI211_X1 port map( C1 => n19363, C2 => n18956, A => n19005, B => 
                           n19004, ZN => n21511);
   U698 : INV_X1 port map( A => n21511, ZN => n21520);
   U699 : AOI211_X1 port map( C1 => n19014, C2 => n19206, A => n18952, B => 
                           n18951, ZN => n21512);
   U700 : OAI222_X1 port map( A1 => n19307, A2 => n21847, B1 => n19412, B2 => 
                           n21520, C1 => n19288, C2 => n21512, ZN => n21896);
   U701 : INV_X1 port map( A => n21896, ZN => n21914);
   U702 : AOI211_X1 port map( C1 => n19204, C2 => n19014, A => n18950, B => 
                           n19001, ZN => n21513);
   U703 : AOI211_X1 port map( C1 => n19014, C2 => n19422, A => n18949, B => 
                           n19000, ZN => n21517);
   U704 : OAI222_X1 port map( A1 => n19307, A2 => n21512, B1 => n19412, B2 => 
                           n21513, C1 => n19288, C2 => n21517, ZN => n22200);
   U705 : OAI222_X1 port map( A1 => n19307, A2 => n21520, B1 => n19412, B2 => 
                           n21512, C1 => n19288, C2 => n21513, ZN => n22182);
   U706 : AOI22_X1 port map( A1 => n19405, A2 => n22200, B1 => n18889, B2 => 
                           n22182, ZN => n21519);
   U707 : AOI211_X1 port map( C1 => n19009, C2 => n19204, A => n18948, B => 
                           n18999, ZN => n22246);
   U708 : OAI22_X1 port map( A1 => n19307, A2 => n21513, B1 => n19288, B2 => 
                           n22246, ZN => n21514);
   U709 : INV_X1 port map( A => n21514, ZN => n21515);
   U710 : OAI21_X1 port map( B1 => n19412, B2 => n21517, A => n21515, ZN => 
                           n22214);
   U711 : AOI22_X1 port map( A1 => n19422, A2 => n19009, B1 => n19204, B2 => 
                           n19414, ZN => n21516);
   U712 : OAI211_X1 port map( C1 => n19313, C2 => n19013, A => n18997, B => 
                           n21516, ZN => n22248);
   U713 : INV_X1 port map( A => n22248, ZN => n22266);
   U714 : OAI222_X1 port map( A1 => n19307, A2 => n21517, B1 => n19412, B2 => 
                           n22246, C1 => n19288, C2 => n22266, ZN => n22227);
   U715 : AOI22_X1 port map( A1 => n19211, A2 => n22214, B1 => n19368, B2 => 
                           n22227, ZN => n21518);
   U716 : OAI211_X1 port map( C1 => n19141, C2 => n21914, A => n21519, B => 
                           n21518, ZN => n22138);
   U717 : INV_X1 port map( A => n22200, ZN => n21523);
   U718 : AOI211_X1 port map( C1 => n19402, C2 => n19386, A => n18955, B => 
                           n18998, ZN => n21848);
   U719 : OAI222_X1 port map( A1 => n19288, A2 => n21520, B1 => n21848, B2 => 
                           n19307, C1 => n21847, C2 => n19412, ZN => n21900);
   U720 : AOI22_X1 port map( A1 => n21900, A2 => n19396, B1 => n22214, B2 => 
                           n19368, ZN => n21522);
   U721 : AOI22_X1 port map( A1 => n22982, A2 => n21896, B1 => n22182, B2 => 
                           n19405, ZN => n21521);
   U722 : OAI211_X1 port map( C1 => n22960, C2 => n21523, A => n21522, B => 
                           n21521, ZN => n21927);
   U723 : AOI22_X1 port map( A1 => n19226, A2 => n22138, B1 => n19320, B2 => 
                           n21927, ZN => n21524);
   U724 : OAI22_X1 port map( A1 => n19316, A2 => n21524, B1 => n19284, B2 => 
                           n18877, ZN => n21525);
   U725 : OR4_X1 port map( A1 => n19435, A2 => n19433, A3 => n21182, A4 => 
                           n21525, ZN => OUTALU(21));
   U726 : INV_X1 port map( A => n9084, ZN => n1795);
   U727 : INV_X1 port map( A => n9081, ZN => n1794);
   U728 : NAND3_X1 port map( A1 => n21527, A2 => n21526, A3 => n1836, ZN => 
                           n1896);
   U729 : INV_X1 port map( A => n1896, ZN => n1835);
   U730 : INV_X1 port map( A => n22081, ZN => n22050);
   U731 : AOI211_X1 port map( C1 => n21528, C2 => n21529, A => n21822, B => 
                           n22050, ZN => n21532);
   U732 : AOI211_X1 port map( C1 => n21530, C2 => n21529, A => n21820, B => 
                           n22063, ZN => n21531);
   U733 : NOR2_X1 port map( A1 => n21532, A2 => n21531, ZN => n13929);
   U734 : INV_X1 port map( A => n21533, ZN => n22953);
   U735 : INV_X1 port map( A => n21544, ZN => n21548);
   U736 : AOI22_X1 port map( A1 => n22941, A2 => n21535, B1 => n22943, B2 => 
                           n21534, ZN => n21537);
   U737 : AOI22_X1 port map( A1 => n22524, A2 => n21554, B1 => n22945, B2 => 
                           n21543, ZN => n21536);
   U738 : OAI211_X1 port map( C1 => n22866, C2 => n21548, A => n21537, B => 
                           n21536, ZN => n21779);
   U739 : AOI22_X1 port map( A1 => n1835, A2 => n1805, B1 => n22953, B2 => 
                           n21779, ZN => n16696);
   U740 : OAI22_X1 port map( A1 => n22530, A2 => n21551, B1 => n22864, B2 => 
                           n21792, ZN => n21539);
   U741 : OAI22_X1 port map( A1 => n22948, A2 => n21541, B1 => n22874, B2 => 
                           n21548, ZN => n21538);
   U742 : AOI211_X1 port map( C1 => n22939, C2 => n21540, A => n21539, B => 
                           n21538, ZN => n21790);
   U743 : INV_X1 port map( A => n21790, ZN => n21547);
   U744 : OAI22_X1 port map( A1 => n22864, A2 => n21541, B1 => n22866, B2 => 
                           n21792, ZN => n21542);
   U745 : INV_X1 port map( A => n21542, ZN => n21546);
   U746 : AOI22_X1 port map( A1 => n22941, A2 => n21544, B1 => n22943, B2 => 
                           n21543, ZN => n21545);
   U747 : OAI211_X1 port map( C1 => n21551, C2 => n22948, A => n21546, B => 
                           n21545, ZN => n21789);
   U748 : AOI22_X1 port map( A1 => n13151, A2 => n21547, B1 => n1894, B2 => 
                           n21789, ZN => n16695);
   U749 : AOI22_X1 port map( A1 => n1843, A2 => n21779, B1 => n13151, B2 => 
                           n21789, ZN => n16700);
   U750 : OAI22_X1 port map( A1 => n22874, A2 => n21549, B1 => n21548, B2 => 
                           n22864, ZN => n21553);
   U751 : OAI22_X1 port map( A1 => n22866, A2 => n21551, B1 => n21550, B2 => 
                           n22948, ZN => n21552);
   U752 : AOI211_X1 port map( C1 => n22873, C2 => n21554, A => n21553, B => 
                           n21552, ZN => n13963);
   U753 : OAI22_X1 port map( A1 => n1831, A2 => n22997, B1 => n13963, B2 => 
                           n1896, ZN => n16698);
   U754 : INV_X1 port map( A => n1805, ZN => n21788);
   U755 : OAI22_X1 port map( A1 => n22273, A2 => n1836, B1 => n21788, B2 => 
                           n22997, ZN => n16702);
   U756 : OAI22_X1 port map( A1 => n22273, A2 => n1837, B1 => n21790, B2 => 
                           n17728, ZN => n16705);
   U757 : OAI22_X1 port map( A1 => n22273, A2 => n1896, B1 => n21790, B2 => 
                           n22997, ZN => n16706);
   U758 : OAI22_X1 port map( A1 => n1831, A2 => n17728, B1 => n21838, B2 => 
                           n22997, ZN => n16709);
   U759 : NAND2_X1 port map( A1 => n7769, A2 => n8978, ZN => n22700);
   U760 : OAI21_X1 port map( B1 => n7769, B2 => n8978, A => n22700, ZN => n1798
                           );
   U761 : INV_X1 port map( A => n4302, ZN => n22926);
   U762 : NOR2_X1 port map( A1 => n22926, A2 => n1798, ZN => n14285);
   U763 : NOR2_X1 port map( A1 => n7769, A2 => n21555, ZN => n21184);
   U764 : NOR2_X1 port map( A1 => n21556, A2 => n21184, ZN => n14281);
   U765 : INV_X1 port map( A => n21557, ZN => n22222);
   U766 : NOR2_X1 port map( A1 => n22222, A2 => n22207, ZN => n14278);
   U767 : AOI22_X1 port map( A1 => n22945, A2 => n21559, B1 => n22939, B2 => 
                           n21558, ZN => n21561);
   U768 : AOI22_X1 port map( A1 => n22941, A2 => n21573, B1 => n22524, B2 => 
                           n21568, ZN => n21560);
   U769 : OAI211_X1 port map( C1 => n22874, C2 => n21574, A => n21561, B => 
                           n21560, ZN => n14004);
   U770 : INV_X1 port map( A => n1824, ZN => n21562);
   U771 : AOI22_X1 port map( A1 => n1894, A2 => n21562, B1 => n22953, B2 => 
                           n14004, ZN => n14000);
   U772 : AOI22_X1 port map( A1 => n1843, A2 => n1828, B1 => n1835, B2 => 
                           n14003, ZN => n13999);
   U773 : OAI22_X1 port map( A1 => n22949, A2 => n22864, B1 => n21563, B2 => 
                           n22948, ZN => n21567);
   U774 : OAI22_X1 port map( A1 => n22874, A2 => n21565, B1 => n22866, B2 => 
                           n21564, ZN => n21566);
   U775 : AOI211_X1 port map( C1 => n22941, C2 => n22942, A => n21567, B => 
                           n21566, ZN => n11449);
   U776 : OAI22_X1 port map( A1 => n1824, A2 => n1896, B1 => n11449, B2 => 
                           n1837, ZN => n13997);
   U777 : OAI22_X1 port map( A1 => n1824, A2 => n17728, B1 => n11449, B2 => 
                           n1896, ZN => n13992);
   U778 : AOI22_X1 port map( A1 => n22941, A2 => n21571, B1 => n22943, B2 => 
                           n21578, ZN => n21570);
   U779 : AOI22_X1 port map( A1 => n22945, A2 => n21573, B1 => n22939, B2 => 
                           n21568, ZN => n21569);
   U780 : OAI211_X1 port map( C1 => n21574, C2 => n22948, A => n21570, B => 
                           n21569, ZN => n21675);
   U781 : AOI22_X1 port map( A1 => n1894, A2 => n1828, B1 => n22953, B2 => 
                           n21675, ZN => n13990);
   U782 : AOI22_X1 port map( A1 => n13151, A2 => n14003, B1 => n1835, B2 => 
                           n14004, ZN => n13989);
   U783 : INV_X1 port map( A => n21571, ZN => n21572);
   U784 : OAI22_X1 port map( A1 => n22874, A2 => n21716, B1 => n21572, B2 => 
                           n22948, ZN => n21577);
   U785 : INV_X1 port map( A => n21573, ZN => n21575);
   U786 : OAI22_X1 port map( A1 => n22866, A2 => n21575, B1 => n21574, B2 => 
                           n22864, ZN => n21576);
   U787 : AOI211_X1 port map( C1 => n22941, C2 => n21578, A => n21577, B => 
                           n21576, ZN => n22893);
   U788 : OAI22_X1 port map( A1 => n22893, A2 => n17728, B1 => n1810, B2 => 
                           n22997, ZN => n13988);
   U789 : OAI22_X1 port map( A1 => n22893, A2 => n1896, B1 => n1810, B2 => 
                           n17728, ZN => n13987);
   U790 : NOR2_X1 port map( A1 => n22881, A2 => n22882, ZN => n22899);
   U791 : INV_X1 port map( A => DATA2(22), ZN => n22578);
   U792 : NOR3_X1 port map( A1 => n22899, A2 => n22578, A3 => n22475, ZN => 
                           n14184);
   U793 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_5_port,
                           ZN => n22928);
   U794 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n22928, ZN => n2808);
   U795 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n2808, ZN => n14182);
   U796 : NOR3_X1 port map( A1 => n19439, A2 => n19213, A3 => n1796, ZN => 
                           n3026);
   U797 : AOI221_X1 port map( B1 => n19213, B2 => n19439, C1 => n1796, C2 => 
                           n19439, A => n3026, ZN => n13884);
   U798 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, ZN => 
                           n21579);
   U799 : NOR3_X1 port map( A1 => n19384, A2 => n1796, A3 => n21579, ZN => 
                           n3030);
   U800 : AOI221_X1 port map( B1 => n19384, B2 => n21579, C1 => n1796, C2 => 
                           n21579, A => n3030, ZN => n13878);
   U801 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_4_8_port, ZN => 
                           n21580);
   U802 : NOR3_X1 port map( A1 => n19387, A2 => n1796, A3 => n21580, ZN => 
                           n3029);
   U803 : AOI21_X1 port map( B1 => n19214, B2 => data1_mul_0_port, A => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, ZN => n21581
                           );
   U804 : NOR2_X1 port map( A1 => n3029, A2 => n21581, ZN => n14176);
   U805 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_5_10_port, ZN => 
                           n21582);
   U806 : NOR3_X1 port map( A1 => n19199, A2 => n1796, A3 => n21582, ZN => 
                           n3028);
   U807 : AOI221_X1 port map( B1 => n19199, B2 => n21582, C1 => n1796, C2 => 
                           n21582, A => n3028, ZN => n13873);
   U808 : NAND2_X1 port map( A1 => n19292, A2 => n21161, ZN => n21583);
   U809 : OAI21_X1 port map( B1 => n19292, B2 => n21161, A => n21583, ZN => 
                           n22765);
   U810 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_6_12_port, ZN => 
                           n21584);
   U811 : NOR3_X1 port map( A1 => n1796, A2 => n22765, A3 => n21584, ZN => 
                           n3027);
   U812 : OR2_X1 port map( A1 => n1796, A2 => n22765, ZN => n21585);
   U813 : AOI21_X1 port map( B1 => n21585, B2 => n21584, A => n3027, ZN => 
                           n13868);
   U814 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n22854);
   U815 : INV_X1 port map( A => n22854, ZN => n22858);
   U816 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN 
                           => n22600);
   U817 : NAND2_X1 port map( A1 => n22600, A2 => data2_mul_1_port, ZN => n22852
                           );
   U818 : INV_X1 port map( A => n22852, ZN => n22857);
   U819 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => n22600, ZN => n22840)
                           ;
   U820 : AOI222_X1 port map( A1 => n22858, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           n22857, B2 => n21214, C1 => n22840, C2 => n9081, ZN 
                           => n21587);
   U821 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n22639);
   U822 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n22639, ZN => n22601);
   U823 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n22601, ZN => n21586
                           );
   U824 : NOR2_X1 port map( A1 => n21587, A2 => n21586, ZN => n3036);
   U825 : AOI21_X1 port map( B1 => n21587, B2 => n21586, A => n3036, ZN => 
                           n14170);
   U826 : OAI22_X1 port map( A1 => n21588, A2 => n22864, B1 => n22874, B2 => 
                           n21793, ZN => n21592);
   U827 : INV_X1 port map( A => n21797, ZN => n21589);
   U828 : OAI22_X1 port map( A1 => n21590, A2 => n22948, B1 => n21589, B2 => 
                           n22530, ZN => n21591);
   U829 : INV_X1 port map( A => n1814, ZN => n22274);
   U830 : OAI21_X1 port map( B1 => n21592, B2 => n21591, A => n22274, ZN => 
                           n14168);
   U831 : INV_X1 port map( A => n1816, ZN => n21593);
   U832 : AOI22_X1 port map( A1 => n1835, A2 => n21593, B1 => n22953, B2 => 
                           n1821, ZN => n16766);
   U833 : INV_X1 port map( A => n1821, ZN => n22950);
   U834 : OAI22_X1 port map( A1 => n22950, A2 => n1896, B1 => n1816, B2 => 
                           n1836, ZN => n16770);
   U835 : INV_X1 port map( A => n1817, ZN => n21594);
   U836 : OAI22_X1 port map( A1 => n22950, A2 => n1837, B1 => n21594, B2 => 
                           n1836, ZN => n16771);
   U837 : AOI22_X1 port map( A1 => n1894, A2 => n14003, B1 => n22953, B2 => 
                           n1830, ZN => n16783);
   U838 : AOI22_X1 port map( A1 => n1843, A2 => n14004, B1 => n1835, B2 => 
                           n1828, ZN => n16782);
   U839 : NOR2_X1 port map( A1 => n21596, A2 => n21595, ZN => n22315);
   U840 : NAND2_X1 port map( A1 => n22268, A2 => n22568, ZN => n22900);
   U841 : AOI211_X1 port map( C1 => n21596, C2 => n21595, A => n22315, B => 
                           n22900, ZN => n21602);
   U842 : INV_X1 port map( A => DATA2(9), ZN => n22590);
   U843 : NAND2_X1 port map( A1 => DATA1(9), A2 => n22590, ZN => n22385);
   U844 : INV_X1 port map( A => n22385, ZN => n22446);
   U845 : NOR2_X1 port map( A1 => DATA1(9), A2 => n22590, ZN => n22444);
   U846 : NOR2_X1 port map( A1 => n22446, A2 => n22444, ZN => n22341);
   U847 : AND2_X1 port map( A1 => n19446, A2 => DATA2_I_8_port, ZN => n21597);
   U848 : NOR2_X1 port map( A1 => n22999, A2 => n22268, ZN => n22283);
   U849 : OAI211_X1 port map( C1 => n21598, C2 => n21597, A => n22283, B => 
                           n22309, ZN => n21600);
   U850 : INV_X1 port map( A => n22899, ZN => n22272);
   U851 : NAND3_X1 port map( A1 => DATA2(9), A2 => DATA1(9), A3 => n22272, ZN 
                           => n21599);
   U852 : OAI211_X1 port map( C1 => n22341, C2 => n22958, A => n21600, B => 
                           n21599, ZN => n21601);
   U853 : AOI211_X1 port map( C1 => n19100, C2 => n22998, A => n21602, B => 
                           n21601, ZN => n16797);
   U854 : OAI22_X1 port map( A1 => n18992, A2 => n19203, B1 => n19205, B2 => 
                           n19008, ZN => n21603);
   U855 : AOI211_X1 port map( C1 => n19216, C2 => n19012, A => n18983, B => 
                           n21603, ZN => n21617);
   U856 : AOI211_X1 port map( C1 => n19204, C2 => n22977, A => n18990, B => 
                           n19419, ZN => n21619);
   U857 : OAI22_X1 port map( A1 => n18992, A2 => n19425, B1 => n19203, B2 => 
                           n19008, ZN => n21604);
   U858 : AOI211_X1 port map( C1 => n19399, C2 => n19204, A => n18984, B => 
                           n21604, ZN => n21623);
   U859 : OAI22_X1 port map( A1 => n19210, A2 => n21619, B1 => n19289, B2 => 
                           n21623, ZN => n21605);
   U860 : INV_X1 port map( A => n21605, ZN => n21606);
   U861 : OAI21_X1 port map( B1 => n19412, B2 => n21617, A => n21606, ZN => 
                           n22277);
   U862 : OAI211_X1 port map( C1 => n19313, C2 => n18992, A => n18995, B => 
                           n18993, ZN => n21626);
   U863 : INV_X1 port map( A => n21626, ZN => n21610);
   U864 : OAI22_X1 port map( A1 => n19408, A2 => n19011, B1 => n19423, B2 => 
                           n21169, ZN => n21607);
   U865 : AOI211_X1 port map( C1 => n19420, C2 => n18994, A => n18991, B => 
                           n21607, ZN => n21618);
   U866 : OAI22_X1 port map( A1 => n19412, A2 => n21618, B1 => n19289, B2 => 
                           n21619, ZN => n21608);
   U867 : INV_X1 port map( A => n21608, ZN => n21609);
   U868 : OAI21_X1 port map( B1 => n19210, B2 => n21610, A => n21609, ZN => 
                           n21661);
   U869 : INV_X1 port map( A => n21661, ZN => n21639);
   U870 : OAI211_X1 port map( C1 => n19398, C2 => n19423, A => n18982, B => 
                           n18981, ZN => n21627);
   U871 : INV_X1 port map( A => n21627, ZN => n21638);
   U872 : OAI222_X1 port map( A1 => n19315, A2 => n21610, B1 => n21638, B2 => 
                           n19210, C1 => n21618, C2 => n19289, ZN => n21611);
   U873 : INV_X1 port map( A => n21611, ZN => n21683);
   U874 : OAI22_X1 port map( A1 => n19409, A2 => n21639, B1 => n19141, B2 => 
                           n21683, ZN => n21621);
   U875 : AOI22_X1 port map( A1 => n19420, A2 => n19400, B1 => n19386, B2 => 
                           n21167, ZN => n21613);
   U876 : AOI22_X1 port map( A1 => n19216, A2 => n22977, B1 => n19422, B2 => 
                           n19399, ZN => n21612);
   U877 : OAI211_X1 port map( C1 => n19421, C2 => n19401, A => n21613, B => 
                           n21612, ZN => n21614);
   U878 : INV_X1 port map( A => n21614, ZN => n22224);
   U879 : OAI22_X1 port map( A1 => n19315, A2 => n21623, B1 => n21617, B2 => 
                           n19334, ZN => n21615);
   U880 : INV_X1 port map( A => n21615, ZN => n21616);
   U881 : OAI21_X1 port map( B1 => n19288, B2 => n22224, A => n21616, ZN => 
                           n22278);
   U882 : INV_X1 port map( A => n22278, ZN => n22286);
   U883 : OAI222_X1 port map( A1 => n19412, A2 => n21619, B1 => n19210, B2 => 
                           n21618, C1 => n19289, C2 => n21617, ZN => n21642);
   U884 : INV_X1 port map( A => n21642, ZN => n22288);
   U885 : OAI22_X1 port map( A1 => n19230, A2 => n22286, B1 => n19146, B2 => 
                           n22288, ZN => n21620);
   U886 : AOI211_X1 port map( C1 => n19211, C2 => n22277, A => n21621, B => 
                           n21620, ZN => n21691);
   U887 : INV_X1 port map( A => n21691, ZN => n22324);
   U888 : AOI22_X1 port map( A1 => n19420, A2 => n19399, B1 => n19206, B2 => 
                           n18921, ZN => n21622);
   U889 : OAI211_X1 port map( C1 => n19356, C2 => n22980, A => n18985, B => 
                           n21622, ZN => n22217);
   U890 : INV_X1 port map( A => n22217, ZN => n22225);
   U891 : OAI222_X1 port map( A1 => n19288, A2 => n22225, B1 => n19315, B2 => 
                           n22224, C1 => n19334, C2 => n21623, ZN => n22279);
   U892 : AOI22_X1 port map( A1 => n19333, A2 => n21661, B1 => n22971, B2 => 
                           n22279, ZN => n21625);
   U893 : AOI22_X1 port map( A1 => n19405, A2 => n22277, B1 => n18889, B2 => 
                           n21642, ZN => n21624);
   U894 : OAI211_X1 port map( C1 => n22286, C2 => n22960, A => n21625, B => 
                           n21624, ZN => n22325);
   U895 : OAI211_X1 port map( C1 => n19363, C2 => n18888, A => n18989, B => 
                           n18988, ZN => n21637);
   U896 : AOI222_X1 port map( A1 => n21627, A2 => n19222, B1 => n21626, B2 => 
                           n19306, C1 => n21637, C2 => n19385, ZN => n21685);
   U897 : OAI22_X1 port map( A1 => n19141, A2 => n21685, B1 => n21683, B2 => 
                           n22968, ZN => n21629);
   U898 : INV_X1 port map( A => n22277, ZN => n22289);
   U899 : OAI22_X1 port map( A1 => n19146, A2 => n21639, B1 => n19229, B2 => 
                           n22289, ZN => n21628);
   U900 : AOI211_X1 port map( C1 => n19211, C2 => n21642, A => n21629, B => 
                           n21628, ZN => n21692);
   U901 : INV_X1 port map( A => n21692, ZN => n21630);
   U902 : AOI222_X1 port map( A1 => n22324, A2 => n19226, B1 => n22325, B2 => 
                           n19319, C1 => n21630, C2 => n19320, ZN => n21631);
   U903 : OAI211_X1 port map( C1 => n19326, C2 => n21631, A => n19186, B => 
                           n19185, ZN => OUTALU(9));
   U904 : NAND2_X1 port map( A1 => n19446, A2 => n22591, ZN => n22382);
   U905 : OAI21_X1 port map( B1 => n19446, B2 => n22591, A => n22382, ZN => 
                           n22354);
   U906 : AOI22_X1 port map( A1 => n19272, A2 => n22998, B1 => n22908, B2 => 
                           n22354, ZN => n13980);
   U907 : NOR3_X1 port map( A1 => n22899, A2 => n22591, A3 => n22969, ZN => 
                           n21634);
   U908 : AOI222_X1 port map( A1 => n21797, A2 => n22092, B1 => n22887, B2 => 
                           n22524, C1 => n21652, C2 => n22873, ZN => n21632);
   U909 : OAI22_X1 port map( A1 => n21635, A2 => n22900, B1 => n21632, B2 => 
                           n1814, ZN => n21633);
   U910 : AOI211_X1 port map( C1 => n22283, C2 => n21635, A => n21634, B => 
                           n21633, ZN => n13978);
   U911 : INV_X1 port map( A => n21675, ZN => n21677);
   U912 : OAI22_X1 port map( A1 => n21677, A2 => n17728, B1 => n22893, B2 => 
                           n22997, ZN => n16808);
   U913 : INV_X1 port map( A => n1828, ZN => n21636);
   U914 : INV_X1 port map( A => n1830, ZN => n21676);
   U915 : OAI22_X1 port map( A1 => n21636, A2 => n1836, B1 => n21676, B2 => 
                           n1896, ZN => n16807);
   U916 : AOI211_X1 port map( C1 => n18996, C2 => n19204, A => n18978, B => 
                           n18977, ZN => n21678);
   U917 : INV_X1 port map( A => n21637, ZN => n21658);
   U918 : OAI222_X1 port map( A1 => n19210, A2 => n21678, B1 => n19289, B2 => 
                           n21638, C1 => n19315, C2 => n21658, ZN => n21719);
   U919 : INV_X1 port map( A => n21719, ZN => n21684);
   U920 : OAI22_X1 port map( A1 => n19141, A2 => n21684, B1 => n21683, B2 => 
                           n22974, ZN => n21641);
   U921 : OAI22_X1 port map( A1 => n19409, A2 => n21685, B1 => n19364, B2 => 
                           n21639, ZN => n21640);
   U922 : AOI211_X1 port map( C1 => n22971, C2 => n21642, A => n21641, B => 
                           n21640, ZN => n21690);
   U923 : INV_X1 port map( A => n21690, ZN => n21723);
   U924 : AOI22_X1 port map( A1 => n19224, A2 => n22325, B1 => n19319, B2 => 
                           n22324, ZN => n21643);
   U925 : OAI21_X1 port map( B1 => n19392, B2 => n21692, A => n21643, ZN => 
                           n21644);
   U926 : AOI21_X1 port map( B1 => n19320, B2 => n21723, A => n21644, ZN => 
                           n21645);
   U927 : OAI211_X1 port map( C1 => n19326, C2 => n21645, A => n18980, B => 
                           n18979, ZN => OUTALU(8));
   U928 : OAI221_X1 port map( B1 => n21165, B2 => n22328, C1 => n19444, C2 => 
                           n22958, A => n22221, ZN => n21649);
   U929 : AOI21_X1 port map( B1 => n22880, B2 => n22877, A => n21646, ZN => 
                           n21651);
   U930 : AOI21_X1 port map( B1 => n22880, B2 => n22875, A => n21646, ZN => 
                           n21650);
   U931 : AOI22_X1 port map( A1 => n22331, A2 => n21651, B1 => n17537, B2 => 
                           n21650, ZN => n21647);
   U932 : NOR2_X1 port map( A1 => n21657, A2 => n21647, ZN => n21648);
   U933 : AOI21_X1 port map( B1 => DATA2(7), B2 => n21649, A => n21648, ZN => 
                           n13977);
   U934 : INV_X1 port map( A => n22331, ZN => n22878);
   U935 : INV_X1 port map( A => n17537, ZN => n22876);
   U936 : OAI22_X1 port map( A1 => n21651, A2 => n22878, B1 => n21650, B2 => 
                           n22876, ZN => n21656);
   U937 : AOI22_X1 port map( A1 => n22941, A2 => n22887, B1 => n22943, B2 => 
                           n21652, ZN => n21654);
   U938 : NOR2_X1 port map( A1 => n21165, A2 => DATA2(7), ZN => n22439);
   U939 : AOI22_X1 port map( A1 => n22439, A2 => n22908, B1 => n22998, B2 => 
                           n19108, ZN => n21653);
   U940 : OAI21_X1 port map( B1 => n21654, B2 => n1814, A => n21653, ZN => 
                           n21655);
   U941 : AOI21_X1 port map( B1 => n21657, B2 => n21656, A => n21655, ZN => 
                           n13976);
   U942 : OAI22_X1 port map( A1 => n21677, A2 => n1896, B1 => n21676, B2 => 
                           n1837, ZN => n16831);
   U943 : AOI211_X1 port map( C1 => n18996, C2 => n19386, A => n18987, B => 
                           n18975, ZN => n21679);
   U944 : OAI222_X1 port map( A1 => n19210, A2 => n21679, B1 => n21678, B2 => 
                           n19315, C1 => n19289, C2 => n21658, ZN => n21751);
   U945 : INV_X1 port map( A => n21751, ZN => n21682);
   U946 : OAI22_X1 port map( A1 => n21683, A2 => n22960, B1 => n21682, B2 => 
                           n22981, ZN => n21660);
   U947 : OAI22_X1 port map( A1 => n19146, A2 => n21685, B1 => n21684, B2 => 
                           n22968, ZN => n21659);
   U948 : AOI211_X1 port map( C1 => n19367, C2 => n21661, A => n21660, B => 
                           n21659, ZN => n21727);
   U949 : OAI22_X1 port map( A1 => n19142, A2 => n21727, B1 => n19392, B2 => 
                           n21690, ZN => n21663);
   U950 : OAI22_X1 port map( A1 => n18890, A2 => n21692, B1 => n19391, B2 => 
                           n21691, ZN => n21662);
   U951 : AOI211_X1 port map( C1 => n19287, C2 => n22325, A => n21663, B => 
                           n21662, ZN => n22889);
   U952 : OAI211_X1 port map( C1 => n22889, C2 => n19271, A => n18976, B => 
                           n19184, ZN => OUTALU(7));
   U953 : OAI21_X1 port map( B1 => n19426, B2 => n22328, A => n22221, ZN => 
                           n21666);
   U954 : OAI22_X1 port map( A1 => n21696, A2 => n22048, B1 => n21664, B2 => 
                           n22520, ZN => n21665);
   U955 : AOI22_X1 port map( A1 => DATA2(5), A2 => n21666, B1 => n22274, B2 => 
                           n21665, ZN => n13974);
   U956 : AOI22_X1 port map( A1 => DATA2(5), A2 => n19299, B1 => n19426, B2 => 
                           n22596, ZN => n22349);
   U957 : AOI22_X1 port map( A1 => n22998, A2 => n19115, B1 => n22908, B2 => 
                           n22349, ZN => n13973);
   U958 : OAI22_X1 port map( A1 => n21668, A2 => n22878, B1 => n21667, B2 => 
                           n22876, ZN => n21673);
   U959 : OAI22_X1 port map( A1 => n22878, A2 => n21670, B1 => n22876, B2 => 
                           n21669, ZN => n21672);
   U960 : INV_X1 port map( A => n21674, ZN => n21671);
   U961 : AOI22_X1 port map( A1 => n21674, A2 => n21673, B1 => n21672, B2 => 
                           n21671, ZN => n13972);
   U962 : INV_X1 port map( A => n1807, ZN => n22896);
   U963 : AOI22_X1 port map( A1 => n13151, A2 => n21675, B1 => n22953, B2 => 
                           n22896, ZN => n13971);
   U964 : OAI22_X1 port map( A1 => n21677, A2 => n1837, B1 => n21676, B2 => 
                           n1836, ZN => n16857);
   U965 : AOI211_X1 port map( C1 => n19406, C2 => n19216, A => n18986, B => 
                           n18970, ZN => n21718);
   U966 : OAI222_X1 port map( A1 => n19210, A2 => n21718, B1 => n21678, B2 => 
                           n19289, C1 => n19315, C2 => n21679, ZN => n21990);
   U967 : AOI22_X1 port map( A1 => n18889, A2 => n21990, B1 => n19211, B2 => 
                           n21719, ZN => n21681);
   U968 : OAI211_X1 port map( C1 => n19363, C2 => n18880, A => n18881, B => 
                           n18971, ZN => n21748);
   U969 : INV_X1 port map( A => n21748, ZN => n21717);
   U970 : OAI222_X1 port map( A1 => n22979, A2 => n21717, B1 => n19289, B2 => 
                           n21679, C1 => n21718, C2 => n19315, ZN => n22160);
   U971 : AOI22_X1 port map( A1 => n19317, A2 => n21751, B1 => n19333, B2 => 
                           n22160, ZN => n21680);
   U972 : OAI211_X1 port map( C1 => n21685, C2 => n19229, A => n21681, B => 
                           n21680, ZN => n22164);
   U973 : OAI22_X1 port map( A1 => n19304, A2 => n21692, B1 => n21727, B2 => 
                           n22978, ZN => n21689);
   U974 : OAI22_X1 port map( A1 => n21683, A2 => n19229, B1 => n21682, B2 => 
                           n22968, ZN => n21687);
   U975 : OAI22_X1 port map( A1 => n19364, A2 => n21685, B1 => n19146, B2 => 
                           n21684, ZN => n21686);
   U976 : AOI211_X1 port map( C1 => n22959, C2 => n21990, A => n21687, B => 
                           n21686, ZN => n21995);
   U977 : OAI22_X1 port map( A1 => n19391, A2 => n21690, B1 => n19392, B2 => 
                           n21995, ZN => n21688);
   U978 : AOI211_X1 port map( C1 => n22976, C2 => n22164, A => n21689, B => 
                           n21688, ZN => n21757);
   U979 : INV_X1 port map( A => n21727, ZN => n21754);
   U980 : OAI22_X1 port map( A1 => n19142, A2 => n21995, B1 => n18890, B2 => 
                           n21690, ZN => n21694);
   U981 : OAI22_X1 port map( A1 => n19332, A2 => n21692, B1 => n21691, B2 => 
                           n22962, ZN => n21693);
   U982 : AOI211_X1 port map( C1 => n22972, C2 => n21754, A => n21694, B => 
                           n21693, ZN => n22890);
   U983 : OAI222_X1 port map( A1 => n19394, A2 => n21757, B1 => n19144, B2 => 
                           n22889, C1 => n19212, C2 => n22890, ZN => n22171);
   U984 : NAND3_X1 port map( A1 => n19321, A2 => n19282, A3 => n22171, ZN => 
                           n21695);
   U985 : NAND4_X1 port map( A1 => n18974, A2 => n18973, A3 => n18972, A4 => 
                           n21695, ZN => OUTALU(5));
   U986 : AOI22_X1 port map( A1 => n21702, A2 => n22331, B1 => n17537, B2 => 
                           n21701, ZN => n13970);
   U987 : NOR3_X1 port map( A1 => n21696, A2 => n1814, A3 => n22520, ZN => 
                           n21700);
   U988 : NAND2_X1 port map( A1 => n22913, A2 => n19300, ZN => n22433);
   U989 : NAND2_X1 port map( A1 => DATA2(4), A2 => n19428, ZN => n22437);
   U990 : AND2_X1 port map( A1 => n22433, A2 => n22437, ZN => n21698);
   U991 : AOI21_X1 port map( B1 => n22881, B2 => n19300, A => n22882, ZN => 
                           n21697);
   U992 : OAI22_X1 port map( A1 => n21698, A2 => n22958, B1 => n21697, B2 => 
                           n22913, ZN => n21699);
   U993 : AOI211_X1 port map( C1 => n22998, C2 => n18872, A => n21700, B => 
                           n21699, ZN => n13969);
   U994 : OAI22_X1 port map( A1 => n21702, A2 => n22878, B1 => n21701, B2 => 
                           n22876, ZN => n13968);
   U995 : INV_X1 port map( A => n1810, ZN => n22894);
   U996 : INV_X1 port map( A => n22155, ZN => n21711);
   U997 : INV_X1 port map( A => n21703, ZN => n21704);
   U998 : NAND3_X1 port map( A1 => n21706, A2 => n21705, A3 => n21704, ZN => 
                           n21707);
   U999 : AOI211_X1 port map( C1 => n21978, C2 => n19298, A => n21708, B => 
                           n21707, ZN => n21737);
   U1000 : AOI22_X1 port map( A1 => n22518, A2 => n21743, B1 => n22516, B2 => 
                           n21709, ZN => n21710);
   U1001 : OAI21_X1 port map( B1 => n21737, B2 => n22520, A => n21710, ZN => 
                           n22526);
   U1002 : AOI22_X1 port map( A1 => n22941, A2 => n21711, B1 => n22943, B2 => 
                           n22526, ZN => n21715);
   U1003 : AOI22_X1 port map( A1 => n22524, A2 => n21713, B1 => n22945, B2 => 
                           n21712, ZN => n21714);
   U1004 : OAI211_X1 port map( C1 => n22866, C2 => n21716, A => n21715, B => 
                           n21714, ZN => n21747);
   U1005 : AOI22_X1 port map( A1 => n1894, A2 => n22894, B1 => n22953, B2 => 
                           n21747, ZN => n13967);
   U1006 : INV_X1 port map( A => n22171, ZN => n21988);
   U1007 : INV_X1 port map( A => n22160, ZN => n21722);
   U1008 : OAI211_X1 port map( C1 => n19308, C2 => n18880, A => n18966, B => 
                           n18879, ZN => n21749);
   U1009 : INV_X1 port map( A => n21749, ZN => n21989);
   U1010 : OAI222_X1 port map( A1 => n21718, A2 => n19289, B1 => n21989, B2 => 
                           n22979, C1 => n21717, C2 => n22963, ZN => n22542);
   U1011 : AOI22_X1 port map( A1 => n19405, A2 => n21990, B1 => n19329, B2 => 
                           n22542, ZN => n21721);
   U1012 : AOI22_X1 port map( A1 => n19211, A2 => n21751, B1 => n22971, B2 => 
                           n21719, ZN => n21720);
   U1013 : OAI211_X1 port map( C1 => n21722, C2 => n22968, A => n21721, B => 
                           n21720, ZN => n22550);
   U1014 : AOI22_X1 port map( A1 => n19287, A2 => n21723, B1 => n19397, B2 => 
                           n22550, ZN => n21726);
   U1015 : INV_X1 port map( A => n21995, ZN => n21724);
   U1016 : AOI22_X1 port map( A1 => n19227, A2 => n22164, B1 => n19319, B2 => 
                           n21724, ZN => n21725);
   U1017 : OAI211_X1 port map( C1 => n19391, C2 => n21727, A => n21726, B => 
                           n21725, ZN => n21996);
   U1018 : OAI22_X1 port map( A1 => n19144, A2 => n22890, B1 => n19212, B2 => 
                           n21757, ZN => n21728);
   U1019 : AOI21_X1 port map( B1 => n22985, B2 => n21996, A => n21728, ZN => 
                           n22560);
   U1020 : OAI22_X1 port map( A1 => n19228, A2 => n21988, B1 => n19143, B2 => 
                           n22560, ZN => n21729);
   U1021 : AOI22_X1 port map( A1 => n19282, A2 => n21729, B1 => n18967, B2 => 
                           n19209, ZN => n21730);
   U1022 : OAI211_X1 port map( C1 => n19209, C2 => n18969, A => n18968, B => 
                           n21730, ZN => OUTALU(4));
   U1023 : NAND2_X1 port map( A1 => n19443, A2 => n22933, ZN => n22432);
   U1024 : NAND2_X1 port map( A1 => DATA2(3), A2 => n19311, ZN => n22431);
   U1025 : NAND2_X1 port map( A1 => n22432, A2 => n22431, ZN => n22355);
   U1026 : NOR2_X1 port map( A1 => n19309, A2 => n21802, ZN => n22148);
   U1027 : AOI21_X1 port map( B1 => n21978, B2 => n19335, A => n22148, ZN => 
                           n21731);
   U1028 : NAND2_X1 port map( A1 => n19443, A2 => n22514, ZN => n21741);
   U1029 : OAI211_X1 port map( C1 => n22017, C2 => n22987, A => n21731, B => 
                           n21741, ZN => n21732);
   U1030 : AOI22_X1 port map( A1 => n22908, A2 => n22355, B1 => n22274, B2 => 
                           n21732, ZN => n13966);
   U1031 : OAI21_X1 port map( B1 => n19311, B2 => n22328, A => n22221, ZN => 
                           n21733);
   U1032 : AOI22_X1 port map( A1 => DATA2(3), A2 => n21733, B1 => n22998, B2 =>
                           n19135, ZN => n13965);
   U1033 : AOI21_X1 port map( B1 => n22862, B2 => n21735, A => n21734, ZN => 
                           n21736);
   U1034 : NAND2_X1 port map( A1 => n22331, A2 => n21736, ZN => n14271);
   U1035 : INV_X1 port map( A => n21737, ZN => n21983);
   U1036 : NOR3_X1 port map( A1 => n21740, A2 => n21739, A3 => n21738, ZN => 
                           n21742);
   U1037 : OAI211_X1 port map( C1 => n22017, C2 => n22970, A => n21742, B => 
                           n21741, ZN => n22154);
   U1038 : AOI222_X1 port map( A1 => n21743, A2 => n22516, B1 => n21983, B2 => 
                           n22518, C1 => n22154, C2 => n21982, ZN => n22525);
   U1039 : OAI22_X1 port map( A1 => n22874, A2 => n22525, B1 => n22155, B2 => 
                           n22948, ZN => n21746);
   U1040 : OAI22_X1 port map( A1 => n22866, A2 => n21744, B1 => n21984, B2 => 
                           n22864, ZN => n21745);
   U1041 : AOI211_X1 port map( C1 => n22941, C2 => n22526, A => n21746, B => 
                           n21745, ZN => n22533);
   U1042 : OAI22_X1 port map( A1 => n1807, A2 => n1896, B1 => n22533, B2 => 
                           n22997, ZN => n13964);
   U1043 : INV_X1 port map( A => n21747, ZN => n22534);
   U1044 : INV_X1 port map( A => n1808, ZN => n21987);
   U1045 : OAI22_X1 port map( A1 => n22534, A2 => n17728, B1 => n21987, B2 => 
                           n1837, ZN => n16909);
   U1046 : INV_X1 port map( A => n22542, ZN => n22163);
   U1047 : AOI211_X1 port map( C1 => n19015, C2 => n19386, A => n18963, B => 
                           n18962, ZN => n22158);
   U1048 : AOI22_X1 port map( A1 => n19222, A2 => n21749, B1 => n19306, B2 => 
                           n21748, ZN => n21750);
   U1049 : OAI21_X1 port map( B1 => n19210, B2 => n22158, A => n21750, ZN => 
                           n22159);
   U1050 : AOI22_X1 port map( A1 => n19396, A2 => n22159, B1 => n22961, B2 => 
                           n22160, ZN => n21753);
   U1051 : AOI22_X1 port map( A1 => n19211, A2 => n21990, B1 => n19368, B2 => 
                           n21751, ZN => n21752);
   U1052 : OAI211_X1 port map( C1 => n22163, C2 => n22968, A => n21753, B => 
                           n21752, ZN => n22536);
   U1053 : AOI22_X1 port map( A1 => n19397, A2 => n22536, B1 => n22972, B2 => 
                           n22550, ZN => n21756);
   U1054 : AOI22_X1 port map( A1 => n19287, A2 => n21754, B1 => n19404, B2 => 
                           n22164, ZN => n21755);
   U1055 : OAI211_X1 port map( C1 => n21995, C2 => n22984, A => n21756, B => 
                           n21755, ZN => n22168);
   U1056 : INV_X1 port map( A => n21757, ZN => n21758);
   U1057 : AOI222_X1 port map( A1 => n22168, A2 => n19285, B1 => n21758, B2 => 
                           n19361, C1 => n21996, C2 => n19389, ZN => n22559);
   U1058 : OAI222_X1 port map( A1 => n19228, A2 => n22560, B1 => n19359, B2 => 
                           n21988, C1 => n19143, C2 => n22559, ZN => n21759);
   U1059 : AOI22_X1 port map( A1 => n19282, A2 => n21759, B1 => n19353, B2 => 
                           n19147, ZN => n21760);
   U1060 : NAND4_X1 port map( A1 => n18964, A2 => n19269, A3 => n18965, A4 => 
                           n21760, ZN => OUTALU(3));
   U1061 : INV_X1 port map( A => n21770, ZN => n21761);
   U1062 : AOI22_X1 port map( A1 => n22524, A2 => n21761, B1 => n22943, B2 => 
                           n21775, ZN => n21764);
   U1063 : AOI22_X1 port map( A1 => n22945, A2 => n21767, B1 => n22939, B2 => 
                           n21762, ZN => n21763);
   U1064 : OAI211_X1 port map( C1 => n21765, C2 => n22530, A => n21764, B => 
                           n21763, ZN => n11966);
   U1065 : AOI22_X1 port map( A1 => n22524, A2 => n21766, B1 => n22943, B2 => 
                           n21784, ZN => n21769);
   U1066 : AOI22_X1 port map( A1 => n22941, A2 => n21775, B1 => n22939, B2 => 
                           n21767, ZN => n21768);
   U1067 : OAI211_X1 port map( C1 => n21770, C2 => n22864, A => n21769, B => 
                           n21768, ZN => n21841);
   U1068 : AOI22_X1 port map( A1 => n1835, A2 => n21841, B1 => n1894, B2 => 
                           n11966, ZN => n13956);
   U1069 : AOI22_X1 port map( A1 => n1843, A2 => n21841, B1 => n1835, B2 => 
                           n11966, ZN => n13955);
   U1070 : INV_X1 port map( A => n1823, ZN => n21840);
   U1071 : AOI22_X1 port map( A1 => n1835, A2 => n21840, B1 => n1894, B2 => 
                           n21841, ZN => n13954);
   U1072 : NOR2_X1 port map( A1 => n22032, A2 => n21802, ZN => n22046);
   U1073 : OAI211_X1 port map( C1 => n21981, C2 => n22495, A => n21772, B => 
                           n21771, ZN => n21773);
   U1074 : AOI211_X1 port map( C1 => n21978, C2 => DATA1(26), A => n22046, B =>
                           n21773, ZN => n21801);
   U1075 : OAI222_X1 port map( A1 => n21495, A2 => n21783, B1 => n22086, B2 => 
                           n21801, C1 => n21774, C2 => n22083, ZN => n21814);
   U1076 : AOI22_X1 port map( A1 => n22524, A2 => n21815, B1 => n22092, B2 => 
                           n21814, ZN => n21777);
   U1077 : AOI22_X1 port map( A1 => n22941, A2 => n21808, B1 => n22939, B2 => 
                           n21775, ZN => n21776);
   U1078 : OAI211_X1 port map( C1 => n21778, C2 => n22864, A => n21777, B => 
                           n21776, ZN => n21843);
   U1079 : AOI22_X1 port map( A1 => n13151, A2 => n11966, B1 => n22953, B2 => 
                           n21843, ZN => n13953);
   U1080 : INV_X1 port map( A => n21779, ZN => n21839);
   U1081 : OAI22_X1 port map( A1 => n21839, A2 => n1896, B1 => n13963, B2 => 
                           n1837, ZN => n13950);
   U1082 : NOR2_X1 port map( A1 => n22495, A2 => n21802, ZN => n22029);
   U1083 : OAI211_X1 port map( C1 => n22017, C2 => n22489, A => n21781, B => 
                           n21780, ZN => n21782);
   U1084 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(29), A => n22029, B =>
                           n21782, ZN => n21805);
   U1085 : OAI222_X1 port map( A1 => n21495, A2 => n21801, B1 => n22086, B2 => 
                           n21805, C1 => n21783, C2 => n22083, ZN => n21816);
   U1086 : AOI22_X1 port map( A1 => n22524, A2 => n21808, B1 => n22943, B2 => 
                           n21816, ZN => n21786);
   U1087 : AOI22_X1 port map( A1 => n22941, A2 => n21814, B1 => n22939, B2 => 
                           n21784, ZN => n21785);
   U1088 : OAI211_X1 port map( C1 => n21787, C2 => n22864, A => n21786, B => 
                           n21785, ZN => n21844);
   U1089 : AOI22_X1 port map( A1 => n1843, A2 => n21843, B1 => n22953, B2 => 
                           n21844, ZN => n13949);
   U1090 : OAI22_X1 port map( A1 => n21788, A2 => n17728, B1 => n21790, B2 => 
                           n1837, ZN => n13947);
   U1091 : INV_X1 port map( A => n21789, ZN => n21798);
   U1092 : OAI22_X1 port map( A1 => n21798, A2 => n1896, B1 => n13963, B2 => 
                           n22997, ZN => n13946);
   U1093 : OAI22_X1 port map( A1 => n21790, A2 => n1896, B1 => n21798, B2 => 
                           n17728, ZN => n13945);
   U1094 : OAI22_X1 port map( A1 => n22874, A2 => n21792, B1 => n21791, B2 => 
                           n22530, ZN => n21796);
   U1095 : OAI22_X1 port map( A1 => n21794, A2 => n22948, B1 => n21793, B2 => 
                           n22864, ZN => n21795);
   U1096 : AOI211_X1 port map( C1 => n21797, C2 => n22939, A => n21796, B => 
                           n21795, ZN => n1802);
   U1097 : OAI22_X1 port map( A1 => n1802, A2 => n1836, B1 => n21798, B2 => 
                           n22997, ZN => n13944);
   U1098 : INV_X1 port map( A => n1804, ZN => n22301);
   U1099 : OAI22_X1 port map( A1 => n22301, A2 => n1836, B1 => n1803, B2 => 
                           n17728, ZN => n13943);
   U1100 : NOR2_X1 port map( A1 => n22001, A2 => n21802, ZN => n22019);
   U1101 : NAND2_X1 port map( A1 => DATA1(28), A2 => n21978, ZN => n22044);
   U1102 : OAI211_X1 port map( C1 => n22511, C2 => n22489, A => n21799, B => 
                           n22044, ZN => n21800);
   U1103 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(30), A => n22019, B =>
                           n21800, ZN => n21807);
   U1104 : OAI222_X1 port map( A1 => n22048, A2 => n21805, B1 => n22086, B2 => 
                           n21807, C1 => n21801, C2 => n22083, ZN => n21813);
   U1105 : AOI22_X1 port map( A1 => n22941, A2 => n21813, B1 => n22945, B2 => 
                           n21814, ZN => n21811);
   U1106 : NOR2_X1 port map( A1 => n22502, A2 => n21802, ZN => n22003);
   U1107 : NAND2_X1 port map( A1 => DATA1(29), A2 => n21978, ZN => n22026);
   U1108 : OAI211_X1 port map( C1 => n22017, C2 => n22495, A => n22026, B => 
                           n21803, ZN => n21804);
   U1109 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(31), A => n22003, B =>
                           n21804, ZN => n21806);
   U1110 : OAI222_X1 port map( A1 => n21495, A2 => n21807, B1 => n22086, B2 => 
                           n21806, C1 => n21805, C2 => n22083, ZN => n21809);
   U1111 : AOI22_X1 port map( A1 => n22943, A2 => n21809, B1 => n22939, B2 => 
                           n21808, ZN => n21810);
   U1112 : NAND2_X1 port map( A1 => n21811, A2 => n21810, ZN => n21812);
   U1113 : AOI21_X1 port map( B1 => n22524, B2 => n21816, A => n21812, ZN => 
                           n13942);
   U1114 : INV_X1 port map( A => n1819, ZN => n22952);
   U1115 : AOI22_X1 port map( A1 => n13151, A2 => n22952, B1 => n1894, B2 => 
                           n21843, ZN => n13941);
   U1116 : AOI22_X1 port map( A1 => n22524, A2 => n21814, B1 => n22943, B2 => 
                           n21813, ZN => n21818);
   U1117 : AOI22_X1 port map( A1 => n22941, A2 => n21816, B1 => n22939, B2 => 
                           n21815, ZN => n21817);
   U1118 : OAI211_X1 port map( C1 => n21819, C2 => n22864, A => n21818, B => 
                           n21817, ZN => n21842);
   U1119 : AOI22_X1 port map( A1 => n1843, A2 => n21842, B1 => n1835, B2 => 
                           n21844, ZN => n13940);
   U1120 : INV_X1 port map( A => n22009, ZN => n21823);
   U1121 : INV_X1 port map( A => n8847, ZN => n21821);
   U1122 : OAI21_X1 port map( B1 => n21823, B2 => n21820, A => n21821, ZN => 
                           n21825);
   U1123 : OAI21_X1 port map( B1 => n21823, B2 => n21822, A => n21821, ZN => 
                           n21824);
   U1124 : OAI22_X1 port map( A1 => n22063, A2 => n21825, B1 => n22050, B2 => 
                           n21824, ZN => n1778);
   U1125 : INV_X1 port map( A => DATA1(31), ZN => n22027);
   U1126 : XNOR2_X1 port map( A => n4293, B => n22027, ZN => n21835);
   U1127 : AOI22_X1 port map( A1 => n22079, A2 => n21825, B1 => n22081, B2 => 
                           n21824, ZN => n22008);
   U1128 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n21826);
   U1129 : OAI21_X1 port map( B1 => n21957, B2 => n21827, A => n21826, ZN => 
                           n21830);
   U1130 : AOI211_X1 port map( C1 => n1801, C2 => n22008, A => n22999, B => 
                           n21830, ZN => n21834);
   U1131 : INV_X1 port map( A => DATA2(31), ZN => n22569);
   U1132 : NAND2_X1 port map( A1 => DATA1(31), A2 => n22569, ZN => n22507);
   U1133 : INV_X1 port map( A => n22507, ZN => n22501);
   U1134 : NAND2_X1 port map( A1 => DATA2(31), A2 => n22027, ZN => n22422);
   U1135 : INV_X1 port map( A => n22422, ZN => n22504);
   U1136 : NOR2_X1 port map( A1 => n22501, A2 => n22504, ZN => n22347);
   U1137 : AOI22_X1 port map( A1 => DATA2(31), A2 => n22882, B1 => n22998, B2 
                           => n19018, ZN => n21829);
   U1138 : NOR2_X1 port map( A1 => n21981, A2 => n1813, ZN => n21952);
   U1139 : OAI221_X1 port map( B1 => n21952, B2 => DATA2(31), C1 => n21952, C2 
                           => n22881, A => DATA1(31), ZN => n21828);
   U1140 : OAI211_X1 port map( C1 => n22347, C2 => n22958, A => n21829, B => 
                           n21828, ZN => n21833);
   U1141 : AOI22_X1 port map( A1 => n22568, A2 => n21830, B1 => n1801, B2 => 
                           n1778, ZN => n21831);
   U1142 : NOR2_X1 port map( A1 => n21831, A2 => n21835, ZN => n21832);
   U1143 : AOI211_X1 port map( C1 => n21835, C2 => n21834, A => n21833, B => 
                           n21832, ZN => n14165);
   U1144 : OAI22_X1 port map( A1 => n21838, A2 => n17728, B1 => n14407, B2 => 
                           n22997, ZN => n17012);
   U1145 : OAI22_X1 port map( A1 => n21839, A2 => n1837, B1 => n13963, B2 => 
                           n1836, ZN => n17011);
   U1146 : AOI22_X1 port map( A1 => n1843, A2 => n1826, B1 => n22953, B2 => 
                           n11966, ZN => n17016);
   U1147 : INV_X1 port map( A => n21841, ZN => n21836);
   U1148 : OAI22_X1 port map( A1 => n21836, A2 => n22997, B1 => n14407, B2 => 
                           n1837, ZN => n17018);
   U1149 : INV_X1 port map( A => n1826, ZN => n21837);
   U1150 : OAI22_X1 port map( A1 => n21838, A2 => n1836, B1 => n21837, B2 => 
                           n1896, ZN => n17017);
   U1151 : OAI22_X1 port map( A1 => n21839, A2 => n1836, B1 => n21838, B2 => 
                           n1896, ZN => n17020);
   U1152 : OAI22_X1 port map( A1 => n1831, A2 => n1837, B1 => n14407, B2 => 
                           n17728, ZN => n17019);
   U1153 : AOI22_X1 port map( A1 => n13151, A2 => n21841, B1 => n1894, B2 => 
                           n21840, ZN => n17068);
   U1154 : AOI22_X1 port map( A1 => n22953, A2 => n21842, B1 => n1894, B2 => 
                           n22952, ZN => n21846);
   U1155 : AOI22_X1 port map( A1 => n1843, A2 => n21844, B1 => n1835, B2 => 
                           n21843, ZN => n21845);
   U1156 : OAI211_X1 port map( C1 => n1823, C2 => n1836, A => n21846, B => 
                           n21845, ZN => n17089);
   U1157 : INV_X1 port map( A => n21900, ZN => n21913);
   U1158 : AOI211_X1 port map( C1 => n18887, C2 => n19422, A => n18944, B => 
                           n18943, ZN => n21849);
   U1159 : OAI222_X1 port map( A1 => n19307, A2 => n21849, B1 => n19288, B2 => 
                           n21847, C1 => n21848, C2 => n19330, ZN => n21911);
   U1160 : AOI211_X1 port map( C1 => n18961, C2 => n19420, A => n18941, B => 
                           n18940, ZN => n21854);
   U1161 : OAI211_X1 port map( C1 => n19308, C2 => n18886, A => n18942, B => 
                           n19418, ZN => n21855);
   U1162 : INV_X1 port map( A => n21855, ZN => n21851);
   U1163 : AOI211_X1 port map( C1 => n19318, C2 => n19216, A => n18939, B => 
                           n18938, ZN => n21850);
   U1164 : OAI222_X1 port map( A1 => n21854, A2 => n19307, B1 => n21851, B2 => 
                           n19412, C1 => n19288, C2 => n21850, ZN => n21857);
   U1165 : AOI22_X1 port map( A1 => n19211, A2 => n21911, B1 => n19325, B2 => 
                           n21857, ZN => n21853);
   U1166 : OAI222_X1 port map( A1 => n19307, A2 => n21850, B1 => n19412, B2 => 
                           n21849, C1 => n19288, C2 => n21848, ZN => n21902);
   U1167 : OAI222_X1 port map( A1 => n21851, A2 => n19307, B1 => n19412, B2 => 
                           n21850, C1 => n19288, C2 => n21849, ZN => n21901);
   U1168 : AOI22_X1 port map( A1 => n19317, A2 => n21902, B1 => n18889, B2 => 
                           n21901, ZN => n21852);
   U1169 : OAI211_X1 port map( C1 => n19230, C2 => n21913, A => n21853, B => 
                           n21852, ZN => n21930);
   U1170 : INV_X1 port map( A => n21901, ZN => n21867);
   U1171 : INV_X1 port map( A => n21854, ZN => n21856);
   U1172 : OAI211_X1 port map( C1 => n19388, C2 => n19408, A => n18959, B => 
                           n19417, ZN => n21860);
   U1173 : AOI222_X1 port map( A1 => n21856, A2 => n19222, B1 => n21855, B2 => 
                           n19305, C1 => n21860, C2 => n19437, ZN => n21875);
   U1174 : OAI22_X1 port map( A1 => n21867, A2 => n22960, B1 => n19409, B2 => 
                           n21875, ZN => n21859);
   U1175 : OAI211_X1 port map( C1 => n19363, C2 => n19388, A => n18960, B => 
                           n19416, ZN => n21864);
   U1176 : AOI222_X1 port map( A1 => n21860, A2 => n19222, B1 => n21864, B2 => 
                           n19437, C1 => n21856, C2 => n19305, ZN => n21863);
   U1177 : INV_X1 port map( A => n21857, ZN => n21868);
   U1178 : OAI22_X1 port map( A1 => n21863, A2 => n19141, B1 => n21868, B2 => 
                           n19146, ZN => n21858);
   U1179 : AOI211_X1 port map( C1 => n22971, C2 => n21902, A => n21859, B => 
                           n21858, ZN => n21907);
   U1180 : OAI211_X1 port map( C1 => n19363, C2 => n19403, A => n18958, B => 
                           n18957, ZN => n21874);
   U1181 : AOI222_X1 port map( A1 => n21864, A2 => n19222, B1 => n21860, B2 => 
                           n19305, C1 => n21874, C2 => n19437, ZN => n21884);
   U1182 : OAI22_X1 port map( A1 => n21868, A2 => n22960, B1 => n21884, B2 => 
                           n19141, ZN => n21862);
   U1183 : OAI22_X1 port map( A1 => n19409, A2 => n21863, B1 => n21875, B2 => 
                           n19146, ZN => n21861);
   U1184 : AOI211_X1 port map( C1 => n22971, C2 => n21901, A => n21862, B => 
                           n21861, ZN => n21908);
   U1185 : OAI22_X1 port map( A1 => n21907, A2 => n18891, B1 => n21908, B2 => 
                           n19331, ZN => n21873);
   U1186 : INV_X1 port map( A => n21863, ZN => n21888);
   U1187 : OAI211_X1 port map( C1 => n19403, C2 => n19308, A => n18954, B => 
                           n18937, ZN => n21880);
   U1188 : AOI222_X1 port map( A1 => n21874, A2 => n19222, B1 => n21864, B2 => 
                           n19305, C1 => n21880, C2 => n19437, ZN => n21882);
   U1189 : OAI22_X1 port map( A1 => n19230, A2 => n21868, B1 => n19141, B2 => 
                           n21882, ZN => n21866);
   U1190 : OAI22_X1 port map( A1 => n19409, A2 => n21884, B1 => n19364, B2 => 
                           n21875, ZN => n21865);
   U1191 : AOI211_X1 port map( C1 => n19317, C2 => n21888, A => n21866, B => 
                           n21865, ZN => n21891);
   U1192 : OAI22_X1 port map( A1 => n19409, A2 => n21868, B1 => n21867, B2 => 
                           n22974, ZN => n21871);
   U1193 : INV_X1 port map( A => n21911, ZN => n21869);
   U1194 : OAI22_X1 port map( A1 => n21875, A2 => n19141, B1 => n19230, B2 => 
                           n21869, ZN => n21870);
   U1195 : AOI211_X1 port map( C1 => n22973, C2 => n21902, A => n21871, B => 
                           n21870, ZN => n21917);
   U1196 : OAI22_X1 port map( A1 => n19142, A2 => n21891, B1 => n21917, B2 => 
                           n22984, ZN => n21872);
   U1197 : AOI211_X1 port map( C1 => n19287, C2 => n21930, A => n21873, B => 
                           n21872, ZN => n21922);
   U1198 : INV_X1 port map( A => n21917, ZN => n21899);
   U1199 : AOI222_X1 port map( A1 => n21880, A2 => n19222, B1 => n19437, B2 => 
                           n18936, C1 => n21874, C2 => n19305, ZN => n21885);
   U1200 : OAI22_X1 port map( A1 => n21884, A2 => n19146, B1 => n19141, B2 => 
                           n21885, ZN => n21877);
   U1201 : OAI22_X1 port map( A1 => n19409, A2 => n21882, B1 => n21875, B2 => 
                           n19230, ZN => n21876);
   U1202 : AOI211_X1 port map( C1 => n19211, C2 => n21888, A => n21877, B => 
                           n21876, ZN => n21890);
   U1203 : OAI22_X1 port map( A1 => n19142, A2 => n21890, B1 => n21907, B2 => 
                           n19391, ZN => n21879);
   U1204 : OAI22_X1 port map( A1 => n21891, A2 => n19393, B1 => n21908, B2 => 
                           n18890, ZN => n21878);
   U1205 : AOI211_X1 port map( C1 => n19287, C2 => n21899, A => n21879, B => 
                           n21878, ZN => n21921);
   U1206 : INV_X1 port map( A => n21907, ZN => n21894);
   U1207 : OAI211_X1 port map( C1 => n19408, C2 => n19183, A => n18947, B => 
                           n18946, ZN => n21881);
   U1208 : AOI222_X1 port map( A1 => n21881, A2 => n19385, B1 => n19222, B2 => 
                           n18936, C1 => n21880, C2 => n19306, ZN => n21883);
   U1209 : OAI22_X1 port map( A1 => n19141, A2 => n21883, B1 => n21882, B2 => 
                           n19146, ZN => n21887);
   U1210 : OAI22_X1 port map( A1 => n19409, A2 => n21885, B1 => n21884, B2 => 
                           n19324, ZN => n21886);
   U1211 : AOI211_X1 port map( C1 => n19368, C2 => n21888, A => n21887, B => 
                           n21886, ZN => n21889);
   U1212 : OAI22_X1 port map( A1 => n19142, A2 => n21889, B1 => n21908, B2 => 
                           n19391, ZN => n21893);
   U1213 : OAI22_X1 port map( A1 => n21891, A2 => n18891, B1 => n19392, B2 => 
                           n21890, ZN => n21892);
   U1214 : AOI211_X1 port map( C1 => n19287, C2 => n21894, A => n21893, B => 
                           n21892, ZN => n21895);
   U1215 : OAI222_X1 port map( A1 => n22994, A2 => n21922, B1 => n19212, B2 => 
                           n21921, C1 => n19328, C2 => n21895, ZN => n21938);
   U1216 : AOI22_X1 port map( A1 => n19368, A2 => n22182, B1 => n19333, B2 => 
                           n21902, ZN => n21898);
   U1217 : AOI22_X1 port map( A1 => n19211, A2 => n21896, B1 => n18889, B2 => 
                           n21911, ZN => n21897);
   U1218 : OAI211_X1 port map( C1 => n21913, C2 => n19146, A => n21898, B => 
                           n21897, ZN => n21931);
   U1219 : AOI22_X1 port map( A1 => n19287, A2 => n21931, B1 => n19226, B2 => 
                           n21899, ZN => n21906);
   U1220 : AOI22_X1 port map( A1 => n19405, A2 => n21911, B1 => n22973, B2 => 
                           n21900, ZN => n21904);
   U1221 : AOI22_X1 port map( A1 => n22982, A2 => n21902, B1 => n22959, B2 => 
                           n21901, ZN => n21903);
   U1222 : OAI211_X1 port map( C1 => n19230, C2 => n21914, A => n21904, B => 
                           n21903, ZN => n21928);
   U1223 : AOI22_X1 port map( A1 => n19225, A2 => n21928, B1 => n19407, B2 => 
                           n21930, ZN => n21905);
   U1224 : OAI211_X1 port map( C1 => n19142, C2 => n21907, A => n21906, B => 
                           n21905, ZN => n21935);
   U1225 : INV_X1 port map( A => n21928, ZN => n21939);
   U1226 : OAI22_X1 port map( A1 => n21917, A2 => n18890, B1 => n21939, B2 => 
                           n19304, ZN => n21910);
   U1227 : OAI22_X1 port map( A1 => n19142, A2 => n21908, B1 => n21907, B2 => 
                           n19393, ZN => n21909);
   U1228 : AOI211_X1 port map( C1 => n19224, C2 => n21930, A => n21910, B => 
                           n21909, ZN => n21923);
   U1229 : AOI22_X1 port map( A1 => n21911, A2 => n19396, B1 => n22182, B2 => 
                           n19211, ZN => n21912);
   U1230 : INV_X1 port map( A => n21912, ZN => n21916);
   U1231 : OAI22_X1 port map( A1 => n19146, A2 => n21914, B1 => n21913, B2 => 
                           n22968, ZN => n21915);
   U1232 : AOI211_X1 port map( C1 => n19368, C2 => n22200, A => n21916, B => 
                           n21915, ZN => n22119);
   U1233 : OAI22_X1 port map( A1 => n21939, A2 => n22978, B1 => n22119, B2 => 
                           n22962, ZN => n21919);
   U1234 : INV_X1 port map( A => n21931, ZN => n22105);
   U1235 : OAI22_X1 port map( A1 => n22105, A2 => n19391, B1 => n21917, B2 => 
                           n22989, ZN => n21918);
   U1236 : AOI211_X1 port map( C1 => n19227, C2 => n21930, A => n21919, B => 
                           n21918, ZN => n21943);
   U1237 : OAI22_X1 port map( A1 => n21923, A2 => n19327, B1 => n21943, B2 => 
                           n22990, ZN => n21920);
   U1238 : AOI21_X1 port map( B1 => n19389, B2 => n21935, A => n21920, ZN => 
                           n21946);
   U1239 : INV_X1 port map( A => n21921, ZN => n21924);
   U1240 : INV_X1 port map( A => n21922, ZN => n21926);
   U1241 : INV_X1 port map( A => n21923, ZN => n21925);
   U1242 : AOI222_X1 port map( A1 => n21924, A2 => n19285, B1 => n21926, B2 => 
                           n19389, C1 => n21925, C2 => n19361, ZN => n21944);
   U1243 : OAI22_X1 port map( A1 => n21946, A2 => n22964, B1 => n19228, B2 => 
                           n21944, ZN => n21937);
   U1244 : AOI222_X1 port map( A1 => n21926, A2 => n19285, B1 => n21935, B2 => 
                           n19361, C1 => n21925, C2 => n19389, ZN => n22010);
   U1245 : INV_X1 port map( A => n21927, ZN => n22117);
   U1246 : INV_X1 port map( A => n22119, ZN => n21929);
   U1247 : AOI22_X1 port map( A1 => n19225, A2 => n21929, B1 => n21928, B2 => 
                           n22972, ZN => n21933);
   U1248 : AOI22_X1 port map( A1 => n19407, A2 => n21931, B1 => n19397, B2 => 
                           n21930, ZN => n21932);
   U1249 : OAI211_X1 port map( C1 => n22117, C2 => n22962, A => n21933, B => 
                           n21932, ZN => n22075);
   U1250 : INV_X1 port map( A => n21943, ZN => n21934);
   U1251 : AOI222_X1 port map( A1 => n21935, A2 => n19285, B1 => n22075, B2 => 
                           n19361, C1 => n21934, C2 => n19389, ZN => n21947);
   U1252 : OAI22_X1 port map( A1 => n22010, A2 => n19359, B1 => n21947, B2 => 
                           n19221, ZN => n21936);
   U1253 : AOI211_X1 port map( C1 => n22988, C2 => n21938, A => n21937, B => 
                           n21936, ZN => n21951);
   U1254 : INV_X1 port map( A => n22075, ZN => n21942);
   U1255 : OAI22_X1 port map( A1 => n19142, A2 => n21939, B1 => n18890, B2 => 
                           n22119, ZN => n21941);
   U1256 : OAI22_X1 port map( A1 => n22105, A2 => n19392, B1 => n22117, B2 => 
                           n19332, ZN => n21940);
   U1257 : AOI211_X1 port map( C1 => n19287, C2 => n22138, A => n21941, B => 
                           n21940, ZN => n22089);
   U1258 : OAI222_X1 port map( A1 => n21943, A2 => n19394, B1 => n21942, B2 => 
                           n19212, C1 => n19144, C2 => n22089, ZN => n22059);
   U1259 : INV_X1 port map( A => n21944, ZN => n21945);
   U1260 : AOI22_X1 port map( A1 => n19366, A2 => n22059, B1 => n19321, B2 => 
                           n21945, ZN => n21949);
   U1261 : INV_X1 port map( A => n21946, ZN => n22023);
   U1262 : INV_X1 port map( A => n21947, ZN => n22041);
   U1263 : AOI22_X1 port map( A1 => n19223, A2 => n22023, B1 => n19220, B2 => 
                           n22041, ZN => n21948);
   U1264 : OAI211_X1 port map( C1 => n19228, C2 => n22010, A => n21949, B => 
                           n21948, ZN => n21958);
   U1265 : NAND3_X1 port map( A1 => n19436, A2 => n19260, A3 => n21958, ZN => 
                           n21950);
   U1266 : OAI211_X1 port map( C1 => n19354, C2 => n21951, A => n18945, B => 
                           n21950, ZN => OUTALU(31));
   U1267 : AOI21_X1 port map( B1 => DATA2(30), B2 => n22272, A => n21952, ZN =>
                           n21955);
   U1268 : INV_X1 port map( A => DATA2(30), ZN => n22570);
   U1269 : AOI22_X1 port map( A1 => DATA1(30), A2 => n22570, B1 => DATA2(30), 
                           B2 => n22502, ZN => n22420);
   U1270 : INV_X1 port map( A => n22420, ZN => n22496);
   U1271 : AOI22_X1 port map( A1 => n19021, A2 => n22313, B1 => n22908, B2 => 
                           n22496, ZN => n21954);
   U1272 : NAND3_X1 port map( A1 => DATA1(31), A2 => n22126, A3 => n22144, ZN 
                           => n21953);
   U1273 : OAI211_X1 port map( C1 => n21955, C2 => n22502, A => n21954, B => 
                           n21953, ZN => n13938);
   U1274 : NOR3_X1 port map( A1 => n1801, A2 => n21957, A3 => n22999, ZN => 
                           n14269);
   U1275 : INV_X1 port map( A => n22008, ZN => n21956);
   U1276 : NAND3_X1 port map( A1 => n1801, A2 => n21957, A3 => n21956, ZN => 
                           n17140);
   U1277 : AOI21_X1 port map( B1 => n21958, B2 => n19281, A => n19182, ZN => 
                           n21959);
   U1278 : NAND2_X1 port map( A1 => n19268, A2 => n21959, ZN => n21960);
   U1279 : NOR2_X1 port map( A1 => n21960, A2 => n18935, ZN => n21961);
   U1280 : OAI21_X1 port map( B1 => n19310, B2 => n19016, A => n21961, ZN => 
                           OUTALU(30));
   U1281 : NOR2_X1 port map( A1 => n19309, A2 => n21981, ZN => n21963);
   U1282 : NAND2_X1 port map( A1 => n19335, A2 => n22144, ZN => n22510);
   U1283 : INV_X1 port map( A => n22510, ZN => n21962);
   U1284 : AOI211_X1 port map( C1 => n21978, C2 => n19303, A => n21963, B => 
                           n21962, ZN => n13936);
   U1285 : AOI211_X1 port map( C1 => n21966, C2 => n21965, A => n21964, B => 
                           n22878, ZN => n21974);
   U1286 : NAND2_X1 port map( A1 => DATA2(2), A2 => n19442, ZN => n21972);
   U1287 : OAI211_X1 port map( C1 => n21969, C2 => n21968, A => n17537, B => 
                           n21967, ZN => n21971);
   U1288 : AOI22_X1 port map( A1 => DATA2(2), A2 => n19442, B1 => n19309, B2 =>
                           n22934, ZN => n22428);
   U1289 : NAND2_X1 port map( A1 => n22428, A2 => n22908, ZN => n21970);
   U1290 : OAI211_X1 port map( C1 => n22899, C2 => n21972, A => n21971, B => 
                           n21970, ZN => n21973);
   U1291 : AOI211_X1 port map( C1 => n19187, C2 => n22998, A => n21974, B => 
                           n21973, ZN => n13935);
   U1292 : OAI22_X1 port map( A1 => n22534, A2 => n1896, B1 => n22533, B2 => 
                           n17728, ZN => n13933);
   U1293 : INV_X1 port map( A => n21975, ZN => n21977);
   U1294 : AOI211_X1 port map( C1 => n21978, C2 => n19300, A => n21977, B => 
                           n21976, ZN => n21980);
   U1295 : OAI211_X1 port map( C1 => n19309, C2 => n21981, A => n21980, B => 
                           n21979, ZN => n22515);
   U1296 : AOI222_X1 port map( A1 => n21983, A2 => n22516, B1 => n22154, B2 => 
                           n22518, C1 => n22515, C2 => n21982, ZN => n22508);
   U1297 : OAI22_X1 port map( A1 => n22874, A2 => n22508, B1 => n22155, B2 => 
                           n22864, ZN => n21986);
   U1298 : OAI22_X1 port map( A1 => n22866, A2 => n21984, B1 => n22525, B2 => 
                           n22530, ZN => n21985);
   U1299 : AOI211_X1 port map( C1 => n22524, C2 => n22526, A => n21986, B => 
                           n21985, ZN => n1806);
   U1300 : OAI22_X1 port map( A1 => n21987, A2 => n1836, B1 => n1806, B2 => 
                           n22997, ZN => n17160);
   U1301 : OAI22_X1 port map( A1 => n19359, A2 => n22560, B1 => n21988, B2 => 
                           n19362, ZN => n21998);
   U1302 : INV_X1 port map( A => n22159, ZN => n22546);
   U1303 : AOI211_X1 port map( C1 => n19006, C2 => n19204, A => n18932, B => 
                           n18931, ZN => n22537);
   U1304 : OAI222_X1 port map( A1 => n19412, A2 => n22158, B1 => n19210, B2 => 
                           n22537, C1 => n19289, C2 => n21989, ZN => n22540);
   U1305 : AOI22_X1 port map( A1 => n19405, A2 => n22542, B1 => n19396, B2 => 
                           n22540, ZN => n21992);
   U1306 : AOI22_X1 port map( A1 => n19368, A2 => n21990, B1 => n22973, B2 => 
                           n22160, ZN => n21991);
   U1307 : OAI211_X1 port map( C1 => n22546, C2 => n22968, A => n21992, B => 
                           n21991, ZN => n22547);
   U1308 : AOI22_X1 port map( A1 => n19397, A2 => n22547, B1 => n19404, B2 => 
                           n22550, ZN => n21994);
   U1309 : AOI22_X1 port map( A1 => n19225, A2 => n22164, B1 => n19227, B2 => 
                           n22536, ZN => n21993);
   U1310 : OAI211_X1 port map( C1 => n19304, C2 => n21995, A => n21994, B => 
                           n21993, ZN => n22554);
   U1311 : AOI222_X1 port map( A1 => n22554, A2 => n19285, B1 => n21996, B2 => 
                           n19361, C1 => n22168, C2 => n19389, ZN => n22558);
   U1312 : OAI22_X1 port map( A1 => n19228, A2 => n22559, B1 => n19143, B2 => 
                           n22558, ZN => n21997);
   U1313 : OAI21_X1 port map( B1 => n21998, B2 => n21997, A => n19282, ZN => 
                           n21999);
   U1314 : OAI211_X1 port map( C1 => n19354, C2 => n18934, A => n18933, B => 
                           n21999, ZN => OUTALU(2));
   U1315 : NOR2_X1 port map( A1 => DATA2(29), A2 => n22001, ZN => n22497);
   U1316 : NAND2_X1 port map( A1 => DATA2(29), A2 => n22001, ZN => n22498);
   U1317 : INV_X1 port map( A => n22498, ZN => n22343);
   U1318 : OR2_X1 port map( A1 => n22497, A2 => n22343, ZN => n22000);
   U1319 : AOI22_X1 port map( A1 => n22998, A2 => n19024, B1 => n22908, B2 => 
                           n22000, ZN => n13932);
   U1320 : OAI21_X1 port map( B1 => n22328, B2 => n22001, A => n22221, ZN => 
                           n22007);
   U1321 : NAND2_X1 port map( A1 => DATA1(29), A2 => n22002, ZN => n22005);
   U1322 : INV_X1 port map( A => n22003, ZN => n22004);
   U1323 : OAI211_X1 port map( C1 => n22016, C2 => n22027, A => n22005, B => 
                           n22004, ZN => n22006);
   U1324 : AOI22_X1 port map( A1 => DATA2(29), A2 => n22007, B1 => n22126, B2 
                           => n22006, ZN => n13931);
   U1325 : AOI21_X1 port map( B1 => n8847, B2 => n22009, A => n22008, ZN => 
                           n14164);
   U1326 : AOI22_X1 port map( A1 => n19223, A2 => n22041, B1 => n19390, B2 => 
                           n22023, ZN => n22013);
   U1327 : INV_X1 port map( A => n22010, ZN => n22011);
   U1328 : AOI22_X1 port map( A1 => n19220, A2 => n22059, B1 => n19395, B2 => 
                           n22011, ZN => n22012);
   U1329 : AOI21_X1 port map( B1 => n22013, B2 => n22012, A => n19354, ZN => 
                           n22014);
   U1330 : AOI211_X1 port map( C1 => n19208, C2 => n18928, A => n19181, B => 
                           n22014, ZN => n22015);
   U1331 : NAND3_X1 port map( A1 => n18930, A2 => n18929, A3 => n22015, ZN => 
                           OUTALU(29));
   U1332 : INV_X1 port map( A => DATA2(28), ZN => n22572);
   U1333 : NOR3_X1 port map( A1 => n22899, A2 => n22572, A3 => n22495, ZN => 
                           n22022);
   U1334 : AOI22_X1 port map( A1 => DATA1(28), A2 => n22572, B1 => DATA2(28), 
                           B2 => n22495, ZN => n22417);
   U1335 : OAI22_X1 port map( A1 => n22027, A2 => n22017, B1 => n22502, B2 => 
                           n22016, ZN => n22018);
   U1336 : AOI211_X1 port map( C1 => n22514, C2 => DATA1(28), A => n22019, B =>
                           n22018, ZN => n22020);
   U1337 : OAI22_X1 port map( A1 => n22417, A2 => n22958, B1 => n22020, B2 => 
                           n1813, ZN => n22021);
   U1338 : AOI211_X1 port map( C1 => n22998, C2 => n19027, A => n22022, B => 
                           n22021, ZN => n14163);
   U1339 : AOI222_X1 port map( A1 => n22059, A2 => n19223, B1 => n22023, B2 => 
                           n19395, C1 => n22041, C2 => n19390, ZN => n22024);
   U1340 : OAI211_X1 port map( C1 => n19354, C2 => n22024, A => n18927, B => 
                           n19283, ZN => OUTALU(28));
   U1341 : OAI22_X1 port map( A1 => n22063, A2 => n22031, B1 => n22050, B2 => 
                           n22030, ZN => n22039);
   U1342 : OAI211_X1 port map( C1 => n22511, C2 => n22027, A => n22026, B => 
                           n22025, ZN => n22028);
   U1343 : AOI211_X1 port map( C1 => DATA1(30), C2 => n22047, A => n22029, B =>
                           n22028, ZN => n22062);
   U1344 : NOR3_X1 port map( A1 => n22062, A2 => n22086, A3 => n1813, ZN => 
                           n22038);
   U1345 : AOI22_X1 port map( A1 => n22079, A2 => n22031, B1 => n22081, B2 => 
                           n22030, ZN => n22036);
   U1346 : NOR2_X1 port map( A1 => DATA2(27), A2 => n22032, ZN => n22491);
   U1347 : INV_X1 port map( A => n22491, ZN => n22033);
   U1348 : NAND2_X1 port map( A1 => DATA2(27), A2 => n22032, ZN => n22492);
   U1349 : NAND2_X1 port map( A1 => n22033, A2 => n22492, ZN => n22350);
   U1350 : AOI22_X1 port map( A1 => n22313, A2 => n19030, B1 => n22908, B2 => 
                           n22350, ZN => n22035);
   U1351 : OAI211_X1 port map( C1 => n22882, C2 => n22881, A => DATA2(27), B =>
                           DATA1(27), ZN => n22034);
   U1352 : OAI211_X1 port map( C1 => n22040, C2 => n22036, A => n22035, B => 
                           n22034, ZN => n22037);
   U1353 : AOI211_X1 port map( C1 => n22040, C2 => n22039, A => n22038, B => 
                           n22037, ZN => n13928);
   U1354 : AOI22_X1 port map( A1 => n19390, A2 => n22059, B1 => n19395, B2 => 
                           n22041, ZN => n22042);
   U1355 : OAI21_X1 port map( B1 => n19354, B2 => n22042, A => n18926, ZN => 
                           OUTALU(27));
   U1356 : OAI211_X1 port map( C1 => n22511, C2 => n22502, A => n22044, B => 
                           n22043, ZN => n22045);
   U1357 : AOI211_X1 port map( C1 => n22047, C2 => DATA1(29), A => n22046, B =>
                           n22045, ZN => n22084);
   U1358 : OAI22_X1 port map( A1 => n22062, A2 => n22048, B1 => n22084, B2 => 
                           n22520, ZN => n22049);
   U1359 : NAND2_X1 port map( A1 => n22126, A2 => n22049, ZN => n14268);
   U1360 : INV_X1 port map( A => DATA2(26), ZN => n22574);
   U1361 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2(26), B1 => n22574, 
                           B2 => n22489, ZN => n22484);
   U1362 : NOR3_X1 port map( A1 => n22899, A2 => n22574, A3 => n22489, ZN => 
                           n22058);
   U1363 : AOI22_X1 port map( A1 => n22079, A2 => n22052, B1 => n22081, B2 => 
                           n22051, ZN => n22056);
   U1364 : OAI22_X1 port map( A1 => n22052, A2 => n22063, B1 => n22051, B2 => 
                           n22050, ZN => n22053);
   U1365 : AOI22_X1 port map( A1 => n19033, A2 => n22313, B1 => n22055, B2 => 
                           n22053, ZN => n22054);
   U1366 : OAI21_X1 port map( B1 => n22056, B2 => n22055, A => n22054, ZN => 
                           n22057);
   U1367 : AOI211_X1 port map( C1 => n22908, C2 => n22484, A => n22058, B => 
                           n22057, ZN => n13927);
   U1368 : NAND3_X1 port map( A1 => n19281, A2 => n19395, A3 => n22059, ZN => 
                           n22060);
   U1369 : NAND3_X1 port map( A1 => n19267, A2 => n18925, A3 => n22060, ZN => 
                           OUTALU(26));
   U1370 : OAI222_X1 port map( A1 => n21495, A2 => n22084, B1 => n22086, B2 => 
                           n22087, C1 => n22062, C2 => n22061, ZN => n22123);
   U1371 : NAND3_X1 port map( A1 => n22126, A2 => n22943, A3 => n22123, ZN => 
                           n14161);
   U1372 : AOI211_X1 port map( C1 => n22078, C2 => n22068, A => n22064, B => 
                           n22063, ZN => n22073);
   U1373 : NOR2_X1 port map( A1 => DATA2(25), A2 => n22065, ZN => n22485);
   U1374 : NAND2_X1 port map( A1 => DATA2(25), A2 => n22065, ZN => n22486);
   U1375 : INV_X1 port map( A => n22486, ZN => n22066);
   U1376 : NOR2_X1 port map( A1 => n22485, A2 => n22066, ZN => n22359);
   U1377 : AOI21_X1 port map( B1 => n22068, B2 => n22080, A => n22067, ZN => 
                           n22069);
   U1378 : NAND2_X1 port map( A1 => n22081, A2 => n22069, ZN => n22071);
   U1379 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n22272, 
                           ZN => n22070);
   U1380 : OAI211_X1 port map( C1 => n22359, C2 => n22958, A => n22071, B => 
                           n22070, ZN => n22072);
   U1381 : AOI211_X1 port map( C1 => n22998, C2 => n19038, A => n22073, B => 
                           n22072, ZN => n17254);
   U1382 : INV_X1 port map( A => n22089, ZN => n22074);
   U1383 : AOI22_X1 port map( A1 => n22075, A2 => n22985, B1 => n22074, B2 => 
                           n22965, ZN => n22076);
   U1384 : OAI211_X1 port map( C1 => n19316, C2 => n22076, A => n19180, B => 
                           n19179, ZN => OUTALU(25));
   U1385 : INV_X1 port map( A => n22080, ZN => n22077);
   U1386 : NAND3_X1 port map( A1 => n22079, A2 => n22078, A3 => n22077, ZN => 
                           n14160);
   U1387 : NAND2_X1 port map( A1 => n22081, A2 => n22080, ZN => n14266);
   U1388 : AOI22_X1 port map( A1 => DATA2(24), A2 => n22881, B1 => 
                           DATA2_I_24_port, B2 => n22081, ZN => n22082);
   U1389 : AOI21_X1 port map( B1 => n22082, B2 => n22221, A => n22483, ZN => 
                           n17270);
   U1390 : INV_X1 port map( A => DATA2(24), ZN => n22576);
   U1391 : AOI22_X1 port map( A1 => DATA1(24), A2 => DATA2(24), B1 => n22576, 
                           B2 => n22483, ZN => n22478);
   U1392 : INV_X1 port map( A => n22478, ZN => n22352);
   U1393 : OAI222_X1 port map( A1 => n22048, A2 => n22087, B1 => n22086, B2 => 
                           n22085, C1 => n22084, C2 => n22083, ZN => n22863);
   U1394 : AOI22_X1 port map( A1 => n22941, A2 => n22123, B1 => n22943, B2 => 
                           n22863, ZN => n22088);
   U1395 : OAI22_X1 port map( A1 => n22352, A2 => n22958, B1 => n22088, B2 => 
                           n1813, ZN => n17269);
   U1396 : AOI211_X1 port map( C1 => n19431, C2 => n19042, A => n19177, B => 
                           n18924, ZN => n22091);
   U1397 : OR3_X1 port map( A1 => n19394, A2 => n22089, A3 => n19354, ZN => 
                           n22090);
   U1398 : NAND4_X1 port map( A1 => n19178, A2 => n19266, A3 => n22091, A4 => 
                           n22090, ZN => OUTALU(24));
   U1399 : AOI21_X1 port map( B1 => DATA2(23), B2 => n22881, A => n22882, ZN =>
                           n14159);
   U1400 : NAND2_X1 port map( A1 => n22998, A2 => n19047, ZN => n14265);
   U1401 : AOI222_X1 port map( A1 => n22114, A2 => n22092, B1 => n22863, B2 => 
                           n22873, C1 => n22123, C2 => n22524, ZN => n22104);
   U1402 : NOR2_X1 port map( A1 => DATA2(23), A2 => n1825, ZN => n22479);
   U1403 : INV_X1 port map( A => n22479, ZN => n22093);
   U1404 : NAND2_X1 port map( A1 => DATA2(23), A2 => n1825, ZN => n22480);
   U1405 : NAND2_X1 port map( A1 => n22093, A2 => n22480, ZN => n22361);
   U1406 : NOR2_X1 port map( A1 => n22100, A2 => n22112, ZN => n22094);
   U1407 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, B1 => 
                           n1809, B2 => n22911, ZN => n22096);
   U1408 : OAI22_X1 port map( A1 => n22098, A2 => n22210, B1 => n22096, B2 => 
                           n22207, ZN => n22110);
   U1409 : AOI22_X1 port map( A1 => n22908, A2 => n22361, B1 => n22094, B2 => 
                           n22110, ZN => n22103);
   U1410 : INV_X1 port map( A => n22095, ZN => n22101);
   U1411 : INV_X1 port map( A => n22207, ZN => n22912);
   U1412 : AND2_X1 port map( A1 => n22912, A2 => n22096, ZN => n22097);
   U1413 : AOI211_X1 port map( C1 => n22098, C2 => n22910, A => n22097, B => 
                           n22112, ZN => n22111);
   U1414 : OAI21_X1 port map( B1 => n22101, B2 => n22111, A => n22100, ZN => 
                           n22099);
   U1415 : OAI211_X1 port map( C1 => n22101, C2 => n22100, A => n22568, B => 
                           n22099, ZN => n22102);
   U1416 : OAI211_X1 port map( C1 => n22104, C2 => n1813, A => n22103, B => 
                           n22102, ZN => n14264);
   U1417 : INV_X1 port map( A => n22138, ZN => n22118);
   U1418 : OAI22_X1 port map( A1 => n18890, A2 => n22117, B1 => n19391, B2 => 
                           n22118, ZN => n22107);
   U1419 : OAI22_X1 port map( A1 => n19142, A2 => n22105, B1 => n22119, B2 => 
                           n19392, ZN => n22106);
   U1420 : AOI221_X1 port map( B1 => n22107, B2 => n19281, C1 => n22106, C2 => 
                           n19281, A => n18923, ZN => n22108);
   U1421 : OAI211_X1 port map( C1 => n19176, C2 => n19432, A => n19265, B => 
                           n22108, ZN => OUTALU(23));
   U1422 : AOI22_X1 port map( A1 => DATA1(22), A2 => n22578, B1 => DATA2(22), 
                           B2 => n22475, ZN => n22477);
   U1423 : INV_X1 port map( A => n22477, ZN => n22109);
   U1424 : AOI22_X1 port map( A1 => n19051, A2 => n22998, B1 => n22908, B2 => 
                           n22109, ZN => n13924);
   U1425 : INV_X1 port map( A => n22110, ZN => n22113);
   U1426 : AOI21_X1 port map( B1 => n22113, B2 => n22112, A => n22111, ZN => 
                           n14158);
   U1427 : AOI22_X1 port map( A1 => n22945, A2 => n22123, B1 => n22873, B2 => 
                           n22114, ZN => n22115);
   U1428 : OAI21_X1 port map( B1 => n22874, B2 => n22868, A => n22115, ZN => 
                           n22116);
   U1429 : AOI21_X1 port map( B1 => n22524, B2 => n22863, A => n22116, ZN => 
                           n14157);
   U1430 : OAI222_X1 port map( A1 => n19142, A2 => n22119, B1 => n18890, B2 => 
                           n22118, C1 => n22117, C2 => n19392, ZN => n22120);
   U1431 : AOI211_X1 port map( C1 => n19281, C2 => n22120, A => n19175, B => 
                           n19202, ZN => n22121);
   U1432 : OAI211_X1 port map( C1 => n19355, C2 => n19174, A => n18922, B => 
                           n22121, ZN => OUTALU(22));
   U1433 : AOI22_X1 port map( A1 => n22941, A2 => n22122, B1 => n22945, B2 => 
                           n22863, ZN => n22125);
   U1434 : AOI22_X1 port map( A1 => n22943, A2 => n22872, B1 => n22123, B2 => 
                           n22939, ZN => n22124);
   U1435 : OAI211_X1 port map( C1 => n22865, C2 => n22948, A => n22125, B => 
                           n22124, ZN => n13985);
   U1436 : NAND3_X1 port map( A1 => n22953, A2 => n22126, A3 => n13985, ZN => 
                           n12313);
   U1437 : INV_X1 port map( A => DATA2(20), ZN => n22580);
   U1438 : NAND2_X1 port map( A1 => DATA1(20), A2 => n22580, ZN => n22471);
   U1439 : NAND2_X1 port map( A1 => DATA2(20), A2 => n22127, ZN => n22474);
   U1440 : NAND2_X1 port map( A1 => n22471, A2 => n22474, ZN => n22338);
   U1441 : NOR3_X1 port map( A1 => n22899, A2 => n22580, A3 => n22127, ZN => 
                           n22137);
   U1442 : NAND2_X1 port map( A1 => n19059, A2 => n22313, ZN => n22135);
   U1443 : OAI211_X1 port map( C1 => n22132, C2 => n22129, A => n22912, B => 
                           n22128, ZN => n22134);
   U1444 : OAI211_X1 port map( C1 => n22132, C2 => n22131, A => n22910, B => 
                           n22130, ZN => n22133);
   U1445 : NAND3_X1 port map( A1 => n22135, A2 => n22134, A3 => n22133, ZN => 
                           n22136);
   U1446 : AOI211_X1 port map( C1 => n22908, C2 => n22338, A => n22137, B => 
                           n22136, ZN => n14263);
   U1447 : AOI22_X1 port map( A1 => n19420, A2 => n18921, B1 => n19216, B2 => 
                           n21167, ZN => n22140);
   U1448 : NAND3_X1 port map( A1 => n19281, A2 => n19320, A3 => n22138, ZN => 
                           n22139);
   U1449 : OAI211_X1 port map( C1 => n19355, C2 => n22140, A => n19172, B => 
                           n22139, ZN => OUTALU(20));
   U1450 : AOI211_X1 port map( C1 => n22329, C2 => n22145, A => n22141, B => 
                           n22878, ZN => n22143);
   U1451 : NOR2_X1 port map( A1 => n19302, A2 => n22919, ZN => n22426);
   U1452 : NAND2_X1 port map( A1 => n19335, A2 => n22919, ZN => n22374);
   U1453 : INV_X1 port map( A => n22374, ZN => n22427);
   U1454 : NOR2_X1 port map( A1 => n22426, A2 => n22427, ZN => n22356);
   U1455 : NOR2_X1 port map( A1 => n22356, A2 => n22958, ZN => n22142);
   U1456 : AOI211_X1 port map( C1 => n18839, C2 => n22998, A => n22143, B => 
                           n22142, ZN => n13922);
   U1457 : AOI21_X1 port map( B1 => n22514, B2 => n22274, A => n22882, ZN => 
                           n22327);
   U1458 : OAI21_X1 port map( B1 => n22919, B2 => n22328, A => n22327, ZN => 
                           n14155);
   U1459 : NAND3_X1 port map( A1 => n19303, A2 => n22144, A3 => n22274, ZN => 
                           n14154);
   U1460 : INV_X1 port map( A => n22146, ZN => n22330);
   U1461 : INV_X1 port map( A => n22145, ZN => n22147);
   U1462 : OAI221_X1 port map( B1 => n22330, B2 => n22147, C1 => n22146, C2 => 
                           n22145, A => n17537, ZN => n13867);
   U1463 : AOI211_X1 port map( C1 => n22514, C2 => n19335, A => n22149, B => 
                           n22148, ZN => n22153);
   U1464 : INV_X1 port map( A => n22150, ZN => n22151);
   U1465 : NAND3_X1 port map( A1 => n22153, A2 => n22152, A3 => n22151, ZN => 
                           n22517);
   U1466 : AOI222_X1 port map( A1 => n22154, A2 => n22516, B1 => n22515, B2 => 
                           n22518, C1 => n22517, C2 => n21982, ZN => n22531);
   U1467 : OAI22_X1 port map( A1 => n22874, A2 => n22531, B1 => n22525, B2 => 
                           n22948, ZN => n22157);
   U1468 : OAI22_X1 port map( A1 => n22866, A2 => n22155, B1 => n22508, B2 => 
                           n22530, ZN => n22156);
   U1469 : AOI211_X1 port map( C1 => n22945, C2 => n22526, A => n22157, B => 
                           n22156, ZN => n22532);
   U1470 : OAI22_X1 port map( A1 => n22533, A2 => n1896, B1 => n22532, B2 => 
                           n22997, ZN => n17360);
   U1471 : OAI22_X1 port map( A1 => n1807, A2 => n1836, B1 => n22534, B2 => 
                           n1837, ZN => n17359);
   U1472 : INV_X1 port map( A => n22550, ZN => n22167);
   U1473 : AOI211_X1 port map( C1 => n19007, C2 => n19420, A => n18919, B => 
                           n18918, ZN => n22539);
   U1474 : OAI222_X1 port map( A1 => n19412, A2 => n22537, B1 => n19210, B2 => 
                           n22539, C1 => n19289, C2 => n22158, ZN => n22543);
   U1475 : AOI22_X1 port map( A1 => n19405, A2 => n22159, B1 => n22959, B2 => 
                           n22543, ZN => n22162);
   U1476 : AOI22_X1 port map( A1 => n18889, A2 => n22540, B1 => n19367, B2 => 
                           n22160, ZN => n22161);
   U1477 : OAI211_X1 port map( C1 => n22163, C2 => n22960, A => n22162, B => 
                           n22161, ZN => n22549);
   U1478 : AOI22_X1 port map( A1 => n19397, A2 => n22549, B1 => n19404, B2 => 
                           n22536, ZN => n22166);
   U1479 : AOI22_X1 port map( A1 => n19226, A2 => n22547, B1 => n22991, B2 => 
                           n22164, ZN => n22165);
   U1480 : OAI211_X1 port map( C1 => n22167, C2 => n19322, A => n22166, B => 
                           n22165, ZN => n22556);
   U1481 : AOI222_X1 port map( A1 => n22556, A2 => n22995, B1 => n22168, B2 => 
                           n19360, C1 => n22554, C2 => n19389, ZN => n22535);
   U1482 : OAI22_X1 port map( A1 => n22559, A2 => n22967, B1 => n22535, B2 => 
                           n22992, ZN => n22170);
   U1483 : OAI22_X1 port map( A1 => n19228, A2 => n22558, B1 => n22560, B2 => 
                           n22964, ZN => n22169);
   U1484 : AOI211_X1 port map( C1 => n19366, C2 => n22171, A => n22170, B => 
                           n22169, ZN => n22567);
   U1485 : INV_X1 port map( A => n22567, ZN => n22172);
   U1486 : AOI22_X1 port map( A1 => n19171, A2 => n19301, B1 => n19282, B2 => 
                           n22172, ZN => n22173);
   U1487 : NAND4_X1 port map( A1 => n19170, A2 => n18860, A3 => n18920, A4 => 
                           n22173, ZN => OUTALU(1));
   U1488 : AOI22_X1 port map( A1 => n22175, A2 => n22910, B1 => n22912, B2 => 
                           n22174, ZN => n22178);
   U1489 : OAI22_X1 port map( A1 => n22175, A2 => n22210, B1 => n22174, B2 => 
                           n22207, ZN => n22176);
   U1490 : NAND2_X1 port map( A1 => n22179, A2 => n22176, ZN => n22177);
   U1491 : OAI21_X1 port map( B1 => n22179, B2 => n22178, A => n22177, ZN => 
                           n13919);
   U1492 : INV_X1 port map( A => DATA2(19), ZN => n22581);
   U1493 : NAND2_X1 port map( A1 => n22581, A2 => DATA1(19), ZN => n22470);
   U1494 : INV_X1 port map( A => n22470, ZN => n22409);
   U1495 : NOR2_X1 port map( A1 => n22581, A2 => DATA1(19), ZN => n22407);
   U1496 : NOR2_X1 port map( A1 => n22409, A2 => n22407, ZN => n22339);
   U1497 : OAI21_X1 port map( B1 => n22328, B2 => n22581, A => n22221, ZN => 
                           n22180);
   U1498 : AOI22_X1 port map( A1 => DATA1(19), A2 => n22180, B1 => n22998, B2 
                           => n19063, ZN => n22181);
   U1499 : OAI21_X1 port map( B1 => n22339, B2 => n22958, A => n22181, ZN => 
                           n17388);
   U1500 : AOI222_X1 port map( A1 => n19420, A2 => n21167, B1 => n19216, B2 => 
                           n18884, C1 => n19422, C2 => n18921, ZN => n22187);
   U1501 : AOI22_X1 port map( A1 => n18889, A2 => n22200, B1 => n19211, B2 => 
                           n22227, ZN => n22184);
   U1502 : AOI22_X1 port map( A1 => n19405, A2 => n22214, B1 => n19396, B2 => 
                           n22182, ZN => n22183);
   U1503 : AOI21_X1 port map( B1 => n22184, B2 => n22183, A => n19354, ZN => 
                           n22185);
   U1504 : NOR3_X1 port map( A1 => n22185, A2 => n18917, A3 => n19264, ZN => 
                           n22186);
   U1505 : OAI21_X1 port map( B1 => n19355, B2 => n22187, A => n22186, ZN => 
                           OUTALU(19));
   U1506 : AOI211_X1 port map( C1 => n22189, C2 => n22194, A => n22188, B => 
                           n22210, ZN => n22199);
   U1507 : INV_X1 port map( A => DATA2(18), ZN => n22582);
   U1508 : NAND2_X1 port map( A1 => DATA1(18), A2 => n22582, ZN => n22464);
   U1509 : INV_X1 port map( A => n22464, ZN => n22190);
   U1510 : AOI21_X1 port map( B1 => DATA2(18), B2 => n22191, A => n22190, ZN =>
                           n22353);
   U1511 : NAND3_X1 port map( A1 => DATA2(18), A2 => DATA1(18), A3 => n22272, 
                           ZN => n22197);
   U1512 : AOI21_X1 port map( B1 => n22194, B2 => n22193, A => n22192, ZN => 
                           n22195);
   U1513 : NAND2_X1 port map( A1 => n22912, A2 => n22195, ZN => n22196);
   U1514 : OAI211_X1 port map( C1 => n22353, C2 => n22958, A => n22197, B => 
                           n22196, ZN => n22198);
   U1515 : AOI211_X1 port map( C1 => n22998, C2 => n19067, A => n22199, B => 
                           n22198, ZN => n14262);
   U1516 : AOI222_X1 port map( A1 => n22227, A2 => n19405, B1 => n22214, B2 => 
                           n18889, C1 => n22200, C2 => n19396, ZN => n22204);
   U1517 : AOI22_X1 port map( A1 => n19422, A2 => n21167, B1 => n18921, B2 => 
                           n19314, ZN => n22201);
   U1518 : OAI21_X1 port map( B1 => n19408, B2 => n18885, A => n22201, ZN => 
                           n22202);
   U1519 : OAI221_X1 port map( B1 => n22202, B2 => n19420, C1 => n22202, C2 => 
                           n18884, A => n19282, ZN => n22203);
   U1520 : OAI211_X1 port map( C1 => n19354, C2 => n22204, A => n18916, B => 
                           n22203, ZN => OUTALU(18));
   U1521 : NOR2_X1 port map( A1 => DATA2(17), A2 => n22205, ZN => n22402);
   U1522 : INV_X1 port map( A => n22402, ZN => n22463);
   U1523 : NAND2_X1 port map( A1 => DATA2(17), A2 => n22205, ZN => n22404);
   U1524 : NAND2_X1 port map( A1 => n22463, A2 => n22404, ZN => n22206);
   U1525 : AOI22_X1 port map( A1 => n22998, A2 => n19071, B1 => n22908, B2 => 
                           n22206, ZN => n13918);
   U1526 : AOI211_X1 port map( C1 => n22209, C2 => n22212, A => n22208, B => 
                           n22207, ZN => n13917);
   U1527 : AOI211_X1 port map( C1 => n22213, C2 => n22212, A => n22211, B => 
                           n22210, ZN => n13916);
   U1528 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n22272, 
                           ZN => n14152);
   U1529 : AOI22_X1 port map( A1 => n22214, A2 => n19396, B1 => n22227, B2 => 
                           n18889, ZN => n22215);
   U1530 : INV_X1 port map( A => n22215, ZN => n22216);
   U1531 : AOI211_X1 port map( C1 => n19281, C2 => n22216, A => n18914, B => 
                           n18913, ZN => n22219);
   U1532 : NAND3_X1 port map( A1 => n19437, A2 => n19282, A3 => n22217, ZN => 
                           n22218);
   U1533 : NAND4_X1 port map( A1 => n18915, A2 => n19169, A3 => n22219, A4 => 
                           n22218, ZN => OUTALU(17));
   U1534 : NOR2_X1 port map( A1 => DATA2(16), A2 => n22398, ZN => n22459);
   U1535 : AOI21_X1 port map( B1 => DATA2(16), B2 => n22398, A => n22459, ZN =>
                           n22340);
   U1536 : INV_X1 port map( A => n22340, ZN => n22220);
   U1537 : AOI22_X1 port map( A1 => n22998, A2 => n19075, B1 => n22908, B2 => 
                           n22220, ZN => n13915);
   U1538 : INV_X1 port map( A => DATA2(16), ZN => n22584);
   U1539 : OAI21_X1 port map( B1 => n22328, B2 => n22584, A => n22221, ZN => 
                           n22223);
   U1540 : AOI22_X1 port map( A1 => DATA1(16), A2 => n22223, B1 => n22222, B2 
                           => n22910, ZN => n14151);
   U1541 : OAI22_X1 port map( A1 => n19315, A2 => n22225, B1 => n22224, B2 => 
                           n19334, ZN => n22226);
   U1542 : AOI21_X1 port map( B1 => n19282, B2 => n22226, A => n19277, ZN => 
                           n22229);
   U1543 : NAND3_X1 port map( A1 => n19396, A2 => n19281, A3 => n22227, ZN => 
                           n22228);
   U1544 : NAND4_X1 port map( A1 => n18911, A2 => n18912, A3 => n22229, A4 => 
                           n22228, ZN => OUTALU(16));
   U1545 : INV_X1 port map( A => n22303, ZN => n22300);
   U1546 : INV_X1 port map( A => n22312, ZN => n22231);
   U1547 : INV_X1 port map( A => n22314, ZN => n22230);
   U1548 : OAI21_X1 port map( B1 => n22231, B2 => n22315, A => n22230, ZN => 
                           n22310);
   U1549 : NAND2_X1 port map( A1 => n22232, A2 => n22310, ZN => n22302);
   U1550 : NAND2_X1 port map( A1 => n22300, A2 => n22302, ZN => n17503);
   U1551 : INV_X1 port map( A => n22235, ZN => n22234);
   U1552 : INV_X1 port map( A => n22240, ZN => n22233);
   U1553 : INV_X1 port map( A => n22283, ZN => n22307);
   U1554 : AOI221_X1 port map( B1 => n22235, B2 => n22240, C1 => n22234, C2 => 
                           n22233, A => n22307, ZN => n22245);
   U1555 : AOI22_X1 port map( A1 => DATA1(15), A2 => n22585, B1 => DATA2(15), 
                           B2 => n22399, ZN => n22358);
   U1556 : NAND3_X1 port map( A1 => DATA2(15), A2 => DATA1(15), A3 => n22272, 
                           ZN => n22243);
   U1557 : NAND2_X1 port map( A1 => n22236, A2 => n17503, ZN => n22903);
   U1558 : AOI21_X1 port map( B1 => n22238, B2 => n22903, A => n22237, ZN => 
                           n22252);
   U1559 : NAND2_X1 port map( A1 => n22252, A2 => n22251, ZN => n22259);
   U1560 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n22263, B2 => n22259, ZN => n22241);
   U1561 : AOI21_X1 port map( B1 => n22241, B2 => n22240, A => n22900, ZN => 
                           n22239);
   U1562 : OAI21_X1 port map( B1 => n22241, B2 => n22240, A => n22239, ZN => 
                           n22242);
   U1563 : OAI211_X1 port map( C1 => n22358, C2 => n22958, A => n22243, B => 
                           n22242, ZN => n22244);
   U1564 : AOI211_X1 port map( C1 => n22998, C2 => n19079, A => n22245, B => 
                           n22244, ZN => n13914);
   U1565 : INV_X1 port map( A => n22246, ZN => n22247);
   U1566 : AOI22_X1 port map( A1 => n19222, A2 => n22248, B1 => n19437, B2 => 
                           n22247, ZN => n22250);
   U1567 : NAND3_X1 port map( A1 => n19325, A2 => n19282, A3 => n22279, ZN => 
                           n22249);
   U1568 : OAI211_X1 port map( C1 => n19354, C2 => n22250, A => n18910, B => 
                           n22249, ZN => OUTALU(15));
   U1569 : INV_X1 port map( A => n22251, ZN => n22255);
   U1570 : INV_X1 port map( A => n22900, ZN => n22316);
   U1571 : AOI22_X1 port map( A1 => n22253, A2 => n22283, B1 => n22316, B2 => 
                           n22252, ZN => n22269);
   U1572 : NOR3_X1 port map( A1 => n22255, A2 => n22269, A3 => n22254, ZN => 
                           n14150);
   U1573 : NAND2_X1 port map( A1 => n21159, A2 => n19294, ZN => n22256);
   U1574 : OAI21_X1 port map( B1 => n21159, B2 => n19294, A => n22256, ZN => 
                           n22802);
   U1575 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_7_14_port, ZN =>
                           n22257);
   U1576 : NOR3_X1 port map( A1 => n19440, A2 => n22802, A3 => n22257, ZN => 
                           n3020);
   U1577 : AOI221_X1 port map( B1 => n19440, B2 => n22257, C1 => n22802, C2 => 
                           n22257, A => n3020, ZN => n13864);
   U1578 : AOI22_X1 port map( A1 => n22316, A2 => n22259, B1 => n22283, B2 => 
                           n22258, ZN => n22262);
   U1579 : OAI22_X1 port map( A1 => n22458, A2 => DATA2(14), B1 => n22586, B2 
                           => DATA1(14), ZN => n22396);
   U1580 : AOI22_X1 port map( A1 => n18856, A2 => n22313, B1 => n22908, B2 => 
                           n22396, ZN => n22261);
   U1581 : NAND3_X1 port map( A1 => DATA2(14), A2 => DATA1(14), A3 => n22272, 
                           ZN => n22260);
   U1582 : OAI211_X1 port map( C1 => n22263, C2 => n22262, A => n22261, B => 
                           n22260, ZN => n13913);
   U1583 : NAND2_X1 port map( A1 => n22274, A2 => n1841, ZN => n17471);
   U1584 : INV_X1 port map( A => n22279, ZN => n22287);
   U1585 : OAI22_X1 port map( A1 => n19409, A2 => n22287, B1 => n19141, B2 => 
                           n22286, ZN => n22264);
   U1586 : AOI211_X1 port map( C1 => n19282, C2 => n22264, A => n19168, B => 
                           n18909, ZN => n22265);
   U1587 : OAI21_X1 port map( B1 => n22266, B2 => n19262, A => n22265, ZN => 
                           OUTALU(14));
   U1588 : INV_X1 port map( A => n22903, ZN => n22901);
   U1589 : NOR3_X1 port map( A1 => n22901, A2 => n22902, A3 => n22999, ZN => 
                           n22267);
   U1590 : OAI211_X1 port map( C1 => n22268, C2 => n22285, A => n22267, B => 
                           n22271, ZN => n13912);
   U1591 : AOI21_X1 port map( B1 => n22271, B2 => n22270, A => n22269, ZN => 
                           n14149);
   U1592 : OAI211_X1 port map( C1 => DATA2(13), C2 => n22882, A => DATA1(13), B
                           => n22272, ZN => n14261);
   U1593 : OAI22_X1 port map( A1 => n22273, A2 => n22997, B1 => n22301, B2 => 
                           n1896, ZN => n22276);
   U1594 : OAI22_X1 port map( A1 => n12526, A2 => n1837, B1 => n1802, B2 => 
                           n17728, ZN => n22275);
   U1595 : OAI21_X1 port map( B1 => n22276, B2 => n22275, A => n22274, ZN => 
                           n17479);
   U1596 : AOI222_X1 port map( A1 => n22961, A2 => n22279, B1 => n22278, B2 => 
                           n22982, C1 => n22277, C2 => n22959, ZN => n22282);
   U1597 : NAND2_X1 port map( A1 => n18908, A2 => n18907, ZN => n22280);
   U1598 : NOR3_X1 port map( A1 => n19167, A2 => n19434, A3 => n22280, ZN => 
                           n22281);
   U1599 : OAI211_X1 port map( C1 => n22282, C2 => n22983, A => n19166, B => 
                           n22281, ZN => OUTALU(13));
   U1600 : INV_X1 port map( A => n22902, ZN => n22904);
   U1601 : INV_X1 port map( A => n22285, ZN => n22284);
   U1602 : OAI221_X1 port map( B1 => n22904, B2 => n22285, C1 => n22902, C2 => 
                           n22284, A => n22283, ZN => n13863);
   U1603 : OAI222_X1 port map( A1 => n1896, A2 => n12526, B1 => n22997, B2 => 
                           n1802, C1 => n17728, C2 => n22301, ZN => n13858);
   U1604 : AOI22_X1 port map( A1 => n19281, A2 => n18849, B1 => n18861, B2 => 
                           n19017, ZN => n22293);
   U1605 : OAI22_X1 port map( A1 => n19364, A2 => n22287, B1 => n19146, B2 => 
                           n22286, ZN => n22291);
   U1606 : OAI22_X1 port map( A1 => n19409, A2 => n22289, B1 => n19141, B2 => 
                           n22288, ZN => n22290);
   U1607 : OAI21_X1 port map( B1 => n22291, B2 => n22290, A => n19282, ZN => 
                           n22292);
   U1608 : NAND4_X1 port map( A1 => n18855, A2 => n18878, A3 => n22293, A4 => 
                           n22292, ZN => OUTALU(12));
   U1609 : INV_X1 port map( A => DATA2(11), ZN => n22588);
   U1610 : NOR3_X1 port map( A1 => n22899, A2 => n22588, A3 => n22294, ZN => 
                           n22297);
   U1611 : NOR2_X1 port map( A1 => DATA1(11), A2 => n22588, ZN => n22450);
   U1612 : INV_X1 port map( A => n22450, ZN => n22363);
   U1613 : NOR2_X1 port map( A1 => DATA2(11), A2 => n22294, ZN => n22387);
   U1614 : INV_X1 port map( A => n22387, ZN => n22295);
   U1615 : AOI21_X1 port map( B1 => n22363, B2 => n22295, A => n22958, ZN => 
                           n22296);
   U1616 : AOI211_X1 port map( C1 => n19092, C2 => n22998, A => n22297, B => 
                           n22296, ZN => n13910);
   U1617 : INV_X1 port map( A => n22298, ZN => n22299);
   U1618 : AOI221_X1 port map( B1 => n22300, B2 => n22299, C1 => n22303, C2 => 
                           n22298, A => n22307, ZN => n13862);
   U1619 : OAI22_X1 port map( A1 => n12526, A2 => n17728, B1 => n22301, B2 => 
                           n22997, ZN => n17505);
   U1620 : INV_X1 port map( A => n22302, ZN => n22304);
   U1621 : AOI21_X1 port map( B1 => n22304, B2 => n22303, A => n22900, ZN => 
                           n17504);
   U1622 : AOI211_X1 port map( C1 => n19261, C2 => n22325, A => n18854, B => 
                           n22996, ZN => n22306);
   U1623 : AOI22_X1 port map( A1 => n19281, A2 => n18905, B1 => n19263, B2 => 
                           n19165, ZN => n22305);
   U1624 : NAND2_X1 port map( A1 => n22306, A2 => n22305, ZN => OUTALU(11));
   U1625 : NOR2_X1 port map( A1 => n22308, A2 => n22307, ZN => n22323);
   U1626 : INV_X1 port map( A => n22309, ZN => n22322);
   U1627 : AOI21_X1 port map( B1 => n22316, B2 => n22310, A => n22323, ZN => 
                           n22311);
   U1628 : AOI21_X1 port map( B1 => n22314, B2 => n22312, A => n22311, ZN => 
                           n22321);
   U1629 : AOI21_X1 port map( B1 => n22881, B2 => DATA2(10), A => n22882, ZN =>
                           n22319);
   U1630 : AOI22_X1 port map( A1 => DATA1(10), A2 => n22589, B1 => DATA2(10), 
                           B2 => n22451, ZN => n22390);
   U1631 : INV_X1 port map( A => n22390, ZN => n22445);
   U1632 : AOI22_X1 port map( A1 => n19194, A2 => n22313, B1 => n22908, B2 => 
                           n22445, ZN => n22318);
   U1633 : NAND3_X1 port map( A1 => n22316, A2 => n22315, A3 => n22314, ZN => 
                           n22317);
   U1634 : OAI211_X1 port map( C1 => n22319, C2 => n22451, A => n22318, B => 
                           n22317, ZN => n22320);
   U1635 : AOI211_X1 port map( C1 => n22323, C2 => n22322, A => n22321, B => 
                           n22320, ZN => n17527);
   U1636 : AOI22_X1 port map( A1 => n19227, A2 => n22325, B1 => n19320, B2 => 
                           n22324, ZN => n22326);
   U1637 : OAI211_X1 port map( C1 => n19326, C2 => n22326, A => n19207, B => 
                           n19164, ZN => OUTALU(10));
   U1638 : OAI21_X1 port map( B1 => n22597, B2 => n22328, A => n22327, ZN => 
                           n22333);
   U1639 : NAND2_X1 port map( A1 => n19303, A2 => n22597, ZN => n22373);
   U1640 : NAND2_X1 port map( A1 => DATA2(0), A2 => n19429, ZN => n22429);
   U1641 : NAND2_X1 port map( A1 => n22373, A2 => n22429, ZN => n22345);
   U1642 : NOR2_X1 port map( A1 => n22330, A2 => n22329, ZN => n22334);
   U1643 : INV_X1 port map( A => n22334, ZN => n22332);
   U1644 : AOI222_X1 port map( A1 => n22333, A2 => n19303, B1 => n22345, B2 => 
                           n22908, C1 => n22332, C2 => n22331, ZN => n13856);
   U1645 : AOI22_X1 port map( A1 => n22998, A2 => n19253, B1 => n17537, B2 => 
                           n22334, ZN => n13908);
   U1646 : INV_X1 port map( A => n22335, ZN => n22337);
   U1647 : NOR2_X1 port map( A1 => n22337, A2 => n22336, ZN => n8626);
   U1648 : NAND2_X1 port map( A1 => FUNC(3), A2 => n8626, ZN => n14259);
   U1649 : INV_X1 port map( A => n22338, ZN => n22342);
   U1650 : NAND4_X1 port map( A1 => n22342, A2 => n22341, A3 => n22340, A4 => 
                           n22339, ZN => n22344);
   U1651 : NOR4_X1 port map( A1 => n22497, A2 => n22345, A3 => n22344, A4 => 
                           n22343, ZN => n22346);
   U1652 : NAND4_X1 port map( A1 => n22347, A2 => n22346, A3 => n22433, A4 => 
                           n22437, ZN => n22370);
   U1653 : INV_X1 port map( A => DATA2(6), ZN => n22595);
   U1654 : AOI22_X1 port map( A1 => DATA2(6), A2 => n19312, B1 => n22970, B2 =>
                           n22595, ZN => n22425);
   U1655 : INV_X1 port map( A => DATA2(12), ZN => n22898);
   U1656 : NOR2_X1 port map( A1 => DATA1(12), A2 => n22898, ZN => n22391);
   U1657 : INV_X1 port map( A => n22391, ZN => n22452);
   U1658 : OAI21_X1 port map( B1 => n22897, B2 => DATA2(12), A => n22452, ZN =>
                           n22907);
   U1659 : OR2_X1 port map( A1 => n22907, A2 => n22387, ZN => n22454);
   U1660 : NAND2_X1 port map( A1 => DATA1(21), A2 => n22579, ZN => n22424);
   U1661 : NOR2_X1 port map( A1 => DATA1(21), A2 => n22579, ZN => n22954);
   U1662 : INV_X1 port map( A => n22954, ZN => n22472);
   U1663 : NAND4_X1 port map( A1 => n22424, A2 => n22472, A3 => n22453, A4 => 
                           n22457, ZN => n22348);
   U1664 : NOR4_X1 port map( A1 => n22425, A2 => n22484, A3 => n22454, A4 => 
                           n22348, ZN => n22368);
   U1665 : INV_X1 port map( A => n22417, ZN => n22490);
   U1666 : NOR4_X1 port map( A1 => n22490, A2 => n22496, A3 => n22350, A4 => 
                           n22349, ZN => n22351);
   U1667 : NAND3_X1 port map( A1 => n22353, A2 => n22352, A3 => n22351, ZN => 
                           n22366);
   U1668 : AOI21_X1 port map( B1 => n21165, B2 => DATA2(7), A => n22354, ZN => 
                           n22384);
   U1669 : INV_X1 port map( A => n22404, ZN => n22466);
   U1670 : INV_X1 port map( A => n22355, ZN => n22357);
   U1671 : NAND4_X1 port map( A1 => n22359, A2 => n22358, A3 => n22357, A4 => 
                           n22356, ZN => n22360);
   U1672 : NOR4_X1 port map( A1 => n22402, A2 => n22466, A3 => n22361, A4 => 
                           n22360, ZN => n22364);
   U1673 : INV_X1 port map( A => n22439, ZN => n22362);
   U1674 : NAND4_X1 port map( A1 => n22384, A2 => n22364, A3 => n22363, A4 => 
                           n22362, ZN => n22365);
   U1675 : NOR4_X1 port map( A1 => n22428, A2 => n22396, A3 => n22366, A4 => 
                           n22365, ZN => n22367);
   U1676 : NAND4_X1 port map( A1 => n22477, A2 => n22390, A3 => n22368, A4 => 
                           n22367, ZN => n22369);
   U1677 : OAI21_X1 port map( B1 => n22370, B2 => n22369, A => n1815, ZN => 
                           n22372);
   U1678 : AOI211_X1 port map( C1 => FUNC(2), C2 => n22372, A => FUNC(1), B => 
                           n22371, ZN => n13907);
   U1679 : NOR2_X1 port map( A1 => DATA2(24), A2 => n22483, ZN => n22415);
   U1680 : OAI22_X1 port map( A1 => n22399, A2 => DATA2(15), B1 => n22458, B2 
                           => DATA2(14), ZN => n22460);
   U1681 : NAND2_X1 port map( A1 => DATA1(12), A2 => n22898, ZN => n22393);
   U1682 : AOI211_X1 port map( C1 => n22374, C2 => n22373, A => n22428, B => 
                           n22426, ZN => n22375);
   U1683 : AOI21_X1 port map( B1 => n19442, B2 => n22934, A => n22375, ZN => 
                           n22376);
   U1684 : AOI22_X1 port map( A1 => DATA2(4), A2 => n19428, B1 => n22376, B2 =>
                           n22432, ZN => n22378);
   U1685 : INV_X1 port map( A => n22433, ZN => n22377);
   U1686 : AOI21_X1 port map( B1 => n22378, B2 => n22431, A => n22377, ZN => 
                           n22379);
   U1687 : OAI21_X1 port map( B1 => DATA2(5), B2 => n19426, A => n22379, ZN => 
                           n22380);
   U1688 : OAI21_X1 port map( B1 => n19299, B2 => n22596, A => n22380, ZN => 
                           n22381);
   U1689 : OAI22_X1 port map( A1 => DATA2(6), A2 => n19427, B1 => n22425, B2 =>
                           n22381, ZN => n22383);
   U1690 : INV_X1 port map( A => n22382, ZN => n22440);
   U1691 : AOI221_X1 port map( B1 => n22439, B2 => n22384, C1 => n22383, C2 => 
                           n22384, A => n22440, ZN => n22386);
   U1692 : OAI21_X1 port map( B1 => n22444, B2 => n22386, A => n22385, ZN => 
                           n22389);
   U1693 : NOR2_X1 port map( A1 => DATA2(10), A2 => n22451, ZN => n22388);
   U1694 : AOI211_X1 port map( C1 => n22390, C2 => n22389, A => n22388, B => 
                           n22387, ZN => n22392);
   U1695 : AOI221_X1 port map( B1 => n22450, B2 => n22393, C1 => n22392, C2 => 
                           n22393, A => n22391, ZN => n22394);
   U1696 : INV_X1 port map( A => n22394, ZN => n22397);
   U1697 : AOI211_X1 port map( C1 => n22457, C2 => n22397, A => n22396, B => 
                           n22395, ZN => n22400);
   U1698 : AOI22_X1 port map( A1 => n22399, A2 => DATA2(15), B1 => n22398, B2 
                           => DATA2(16), ZN => n22461);
   U1699 : OAI21_X1 port map( B1 => n22460, B2 => n22400, A => n22461, ZN => 
                           n22401);
   U1700 : INV_X1 port map( A => n22401, ZN => n22403);
   U1701 : AOI221_X1 port map( B1 => n22459, B2 => n22404, C1 => n22403, C2 => 
                           n22404, A => n22402, ZN => n22406);
   U1702 : NOR2_X1 port map( A1 => DATA1(18), A2 => n22582, ZN => n22405);
   U1703 : OAI21_X1 port map( B1 => n22406, B2 => n22405, A => n22464, ZN => 
                           n22408);
   U1704 : INV_X1 port map( A => n22407, ZN => n22467);
   U1705 : OAI211_X1 port map( C1 => n22409, C2 => n22408, A => n22467, B => 
                           n22474, ZN => n22410);
   U1706 : OAI221_X1 port map( B1 => n22954, B2 => n22471, C1 => n22954, C2 => 
                           n22410, A => n22424, ZN => n22412);
   U1707 : NOR2_X1 port map( A1 => DATA2(22), A2 => n22475, ZN => n22411);
   U1708 : AOI211_X1 port map( C1 => n22477, C2 => n22412, A => n22411, B => 
                           n22479, ZN => n22413);
   U1709 : AOI211_X1 port map( C1 => DATA2(23), C2 => n1825, A => n22413, B => 
                           n22478, ZN => n22414);
   U1710 : AOI221_X1 port map( B1 => n22415, B2 => n22486, C1 => n22414, C2 => 
                           n22486, A => n22485, ZN => n22416);
   U1711 : OAI22_X1 port map( A1 => DATA2(26), A2 => n22489, B1 => n22416, B2 
                           => n22484, ZN => n22418);
   U1712 : OAI211_X1 port map( C1 => n22491, C2 => n22418, A => n22417, B => 
                           n22492, ZN => n22419);
   U1713 : OAI21_X1 port map( B1 => DATA2(28), B2 => n22495, A => n22419, ZN =>
                           n22421);
   U1714 : OAI211_X1 port map( C1 => n22497, C2 => n22421, A => n22420, B => 
                           n22498, ZN => n22423);
   U1715 : OAI211_X1 port map( C1 => DATA2(30), C2 => n22502, A => n22423, B =>
                           n22422, ZN => n22506);
   U1716 : INV_X1 port map( A => n22424, ZN => n22955);
   U1717 : AOI22_X1 port map( A1 => DATA2(6), A2 => n19427, B1 => n21165, B2 =>
                           DATA2(7), ZN => n22442);
   U1718 : INV_X1 port map( A => n22425, ZN => n22885);
   U1719 : INV_X1 port map( A => n22426, ZN => n22430);
   U1720 : AOI211_X1 port map( C1 => n22430, C2 => n22429, A => n22428, B => 
                           n22427, ZN => n22435);
   U1721 : OAI21_X1 port map( B1 => n19442, B2 => n22934, A => n22431, ZN => 
                           n22434);
   U1722 : OAI211_X1 port map( C1 => n22435, C2 => n22434, A => n22433, B => 
                           n22432, ZN => n22436);
   U1723 : OAI211_X1 port map( C1 => n19299, C2 => n22596, A => n22437, B => 
                           n22436, ZN => n22438);
   U1724 : OAI211_X1 port map( C1 => DATA2(5), C2 => n19426, A => n22885, B => 
                           n22438, ZN => n22441);
   U1725 : AOI211_X1 port map( C1 => n22442, C2 => n22441, A => n22440, B => 
                           n22439, ZN => n22443);
   U1726 : AOI21_X1 port map( B1 => DATA2(8), B2 => n22969, A => n22443, ZN => 
                           n22448);
   U1727 : INV_X1 port map( A => n22444, ZN => n22447);
   U1728 : AOI211_X1 port map( C1 => n22448, C2 => n22447, A => n22446, B => 
                           n22445, ZN => n22449);
   U1729 : AOI211_X1 port map( C1 => DATA2(10), C2 => n22451, A => n22450, B =>
                           n22449, ZN => n22455);
   U1730 : OAI211_X1 port map( C1 => n22455, C2 => n22454, A => n22453, B => 
                           n22452, ZN => n22456);
   U1731 : AOI22_X1 port map( A1 => DATA2(14), A2 => n22458, B1 => n22457, B2 
                           => n22456, ZN => n22462);
   U1732 : AOI221_X1 port map( B1 => n22462, B2 => n22461, C1 => n22460, C2 => 
                           n22461, A => n22459, ZN => n22465);
   U1733 : OAI211_X1 port map( C1 => n22466, C2 => n22465, A => n22464, B => 
                           n22463, ZN => n22468);
   U1734 : OAI211_X1 port map( C1 => DATA1(18), C2 => n22582, A => n22468, B =>
                           n22467, ZN => n22469);
   U1735 : NAND3_X1 port map( A1 => n22471, A2 => n22470, A3 => n22469, ZN => 
                           n22473);
   U1736 : OAI221_X1 port map( B1 => n22955, B2 => n22474, C1 => n22955, C2 => 
                           n22473, A => n22472, ZN => n22476);
   U1737 : AOI22_X1 port map( A1 => n22477, A2 => n22476, B1 => DATA2(22), B2 
                           => n22475, ZN => n22481);
   U1738 : AOI211_X1 port map( C1 => n22481, C2 => n22480, A => n22479, B => 
                           n22478, ZN => n22482);
   U1739 : AOI21_X1 port map( B1 => DATA2(24), B2 => n22483, A => n22482, ZN =>
                           n22487);
   U1740 : AOI211_X1 port map( C1 => n22487, C2 => n22486, A => n22485, B => 
                           n22484, ZN => n22488);
   U1741 : AOI21_X1 port map( B1 => DATA2(26), B2 => n22489, A => n22488, ZN =>
                           n22493);
   U1742 : AOI211_X1 port map( C1 => n22493, C2 => n22492, A => n22491, B => 
                           n22490, ZN => n22494);
   U1743 : AOI21_X1 port map( B1 => DATA2(28), B2 => n22495, A => n22494, ZN =>
                           n22499);
   U1744 : AOI211_X1 port map( C1 => n22499, C2 => n22498, A => n22497, B => 
                           n22496, ZN => n22500);
   U1745 : AOI211_X1 port map( C1 => DATA2(30), C2 => n22502, A => n22501, B =>
                           n22500, ZN => n22503);
   U1746 : AOI221_X1 port map( B1 => n22504, B2 => n1815, C1 => n22503, C2 => 
                           n1815, A => FUNC(2), ZN => n22505);
   U1747 : OAI221_X1 port map( B1 => n1815, B2 => n22507, C1 => n1815, C2 => 
                           n22506, A => n22505, ZN => n13906);
   U1748 : INV_X1 port map( A => n22508, ZN => n22523);
   U1749 : OAI211_X1 port map( C1 => n19428, C2 => n22511, A => n22510, B => 
                           n22509, ZN => n22512);
   U1750 : AOI211_X1 port map( C1 => n22514, C2 => n19303, A => n22513, B => 
                           n22512, ZN => n22521);
   U1751 : AOI22_X1 port map( A1 => n22518, A2 => n22517, B1 => n22516, B2 => 
                           n22515, ZN => n22519);
   U1752 : OAI21_X1 port map( B1 => n22521, B2 => n22520, A => n22519, ZN => 
                           n22522);
   U1753 : AOI22_X1 port map( A1 => n22524, A2 => n22523, B1 => n22943, B2 => 
                           n22522, ZN => n22529);
   U1754 : INV_X1 port map( A => n22525, ZN => n22527);
   U1755 : AOI22_X1 port map( A1 => n22945, A2 => n22527, B1 => n22939, B2 => 
                           n22526, ZN => n22528);
   U1756 : OAI211_X1 port map( C1 => n22531, C2 => n22530, A => n22529, B => 
                           n22528, ZN => n17735);
   U1757 : OAI22_X1 port map( A1 => n1806, A2 => n1896, B1 => n22532, B2 => 
                           n17728, ZN => n17734);
   U1758 : OAI22_X1 port map( A1 => n22534, A2 => n1836, B1 => n22533, B2 => 
                           n1837, ZN => n17733);
   U1759 : INV_X1 port map( A => n22535, ZN => n22563);
   U1760 : INV_X1 port map( A => n22536, ZN => n22553);
   U1761 : AOI211_X1 port map( C1 => n18902, C2 => n19216, A => n18901, B => 
                           n18900, ZN => n22538);
   U1762 : OAI222_X1 port map( A1 => n19412, A2 => n22539, B1 => n19210, B2 => 
                           n22538, C1 => n19289, C2 => n22537, ZN => n22541);
   U1763 : AOI22_X1 port map( A1 => n19396, A2 => n22541, B1 => n22961, B2 => 
                           n22540, ZN => n22545);
   U1764 : AOI22_X1 port map( A1 => n18889, A2 => n22543, B1 => n19367, B2 => 
                           n22542, ZN => n22544);
   U1765 : OAI211_X1 port map( C1 => n22546, C2 => n22960, A => n22545, B => 
                           n22544, ZN => n22548);
   U1766 : AOI22_X1 port map( A1 => n19397, A2 => n22548, B1 => n19404, B2 => 
                           n22547, ZN => n22552);
   U1767 : AOI22_X1 port map( A1 => n19287, A2 => n22550, B1 => n19226, B2 => 
                           n22549, ZN => n22551);
   U1768 : OAI211_X1 port map( C1 => n22553, C2 => n19322, A => n22552, B => 
                           n22551, ZN => n22555);
   U1769 : AOI222_X1 port map( A1 => n22556, A2 => n22965, B1 => n22555, B2 => 
                           n19286, C1 => n22554, C2 => n19360, ZN => n22557);
   U1770 : OAI22_X1 port map( A1 => n19359, A2 => n22558, B1 => n19143, B2 => 
                           n22557, ZN => n22562);
   U1771 : OAI22_X1 port map( A1 => n22560, A2 => n22993, B1 => n22559, B2 => 
                           n22964, ZN => n22561);
   U1772 : AOI211_X1 port map( C1 => n19323, C2 => n22563, A => n22562, B => 
                           n22561, ZN => n22564);
   U1773 : OAI211_X1 port map( C1 => n19355, C2 => n22564, A => n18848, B => 
                           n18904, ZN => n22565);
   U1774 : AOI21_X1 port map( B1 => n18903, B2 => n18853, A => n22565, ZN => 
                           n22566);
   U1775 : OAI21_X1 port map( B1 => n19259, B2 => n22567, A => n22566, ZN => 
                           OUTALU(0));
   U1776 : NAND2_X1 port map( A1 => n22568, A2 => n1815, ZN => n22599);
   U1777 : CLKBUF_X1 port map( A => n22599, Z => n22593);
   U1778 : NAND2_X1 port map( A1 => FUNC(3), A2 => n22568, ZN => n22598);
   U1779 : AOI22_X1 port map( A1 => DATA2(31), A2 => n22593, B1 => n22592, B2 
                           => n22569, ZN => N2548);
   U1780 : AOI22_X1 port map( A1 => DATA2(30), A2 => n22599, B1 => n22598, B2 
                           => n22570, ZN => N2547);
   U1781 : INV_X1 port map( A => DATA2(29), ZN => n22571);
   U1782 : AOI22_X1 port map( A1 => DATA2(29), A2 => n22593, B1 => n22592, B2 
                           => n22571, ZN => N2546);
   U1783 : AOI22_X1 port map( A1 => DATA2(28), A2 => n22599, B1 => n22598, B2 
                           => n22572, ZN => N2545);
   U1784 : INV_X1 port map( A => DATA2(27), ZN => n22573);
   U1785 : AOI22_X1 port map( A1 => DATA2(27), A2 => n22593, B1 => n22592, B2 
                           => n22573, ZN => N2544);
   U1786 : AOI22_X1 port map( A1 => DATA2(26), A2 => n22599, B1 => n22598, B2 
                           => n22574, ZN => N2543);
   U1787 : INV_X1 port map( A => DATA2(25), ZN => n22575);
   U1788 : AOI22_X1 port map( A1 => DATA2(25), A2 => n22593, B1 => n22592, B2 
                           => n22575, ZN => N2542);
   U1789 : AOI22_X1 port map( A1 => DATA2(24), A2 => n22599, B1 => n22598, B2 
                           => n22576, ZN => N2541);
   U1790 : INV_X1 port map( A => DATA2(23), ZN => n22577);
   U1791 : AOI22_X1 port map( A1 => DATA2(23), A2 => n22593, B1 => n22592, B2 
                           => n22577, ZN => N2540);
   U1792 : AOI22_X1 port map( A1 => DATA2(22), A2 => n22599, B1 => n22598, B2 
                           => n22578, ZN => N2539);
   U1793 : AOI22_X1 port map( A1 => DATA2(21), A2 => n22599, B1 => n22598, B2 
                           => n22579, ZN => N2538);
   U1794 : AOI22_X1 port map( A1 => DATA2(20), A2 => n22599, B1 => n22598, B2 
                           => n22580, ZN => N2537);
   U1795 : AOI22_X1 port map( A1 => DATA2(19), A2 => n22593, B1 => n22592, B2 
                           => n22581, ZN => N2536);
   U1796 : AOI22_X1 port map( A1 => DATA2(18), A2 => n22593, B1 => n22592, B2 
                           => n22582, ZN => N2535);
   U1797 : INV_X1 port map( A => DATA2(17), ZN => n22583);
   U1798 : AOI22_X1 port map( A1 => DATA2(17), A2 => n22593, B1 => n22592, B2 
                           => n22583, ZN => N2534);
   U1799 : AOI22_X1 port map( A1 => DATA2(16), A2 => n22593, B1 => n22592, B2 
                           => n22584, ZN => N2533);
   U1800 : AOI22_X1 port map( A1 => DATA2(15), A2 => n22593, B1 => n22592, B2 
                           => n22585, ZN => N2532);
   U1801 : AOI22_X1 port map( A1 => DATA2(14), A2 => n22593, B1 => n22592, B2 
                           => n22586, ZN => N2531);
   U1802 : AOI22_X1 port map( A1 => DATA2(13), A2 => n22593, B1 => n22592, B2 
                           => n22587, ZN => N2530);
   U1803 : AOI22_X1 port map( A1 => DATA2(12), A2 => n22593, B1 => n22592, B2 
                           => n22898, ZN => N2529);
   U1804 : AOI22_X1 port map( A1 => DATA2(11), A2 => n22593, B1 => n22592, B2 
                           => n22588, ZN => N2528);
   U1805 : AOI22_X1 port map( A1 => DATA2(10), A2 => n22593, B1 => n22592, B2 
                           => n22589, ZN => N2527);
   U1806 : AOI22_X1 port map( A1 => DATA2(9), A2 => n22593, B1 => n22592, B2 =>
                           n22590, ZN => N2526);
   U1807 : AOI22_X1 port map( A1 => DATA2(8), A2 => n22593, B1 => n22592, B2 =>
                           n22591, ZN => N2525);
   U1808 : INV_X1 port map( A => DATA2(7), ZN => n22594);
   U1809 : AOI22_X1 port map( A1 => DATA2(7), A2 => n22599, B1 => n22598, B2 =>
                           n22594, ZN => N2524);
   U1810 : AOI22_X1 port map( A1 => DATA2(6), A2 => n22599, B1 => n22598, B2 =>
                           n22595, ZN => N2523);
   U1811 : AOI22_X1 port map( A1 => DATA2(5), A2 => n22599, B1 => n22598, B2 =>
                           n22596, ZN => N2522);
   U1812 : AOI22_X1 port map( A1 => DATA2(4), A2 => n22599, B1 => n22598, B2 =>
                           n22913, ZN => N2521);
   U1813 : AOI22_X1 port map( A1 => DATA2(3), A2 => n22599, B1 => n22598, B2 =>
                           n22933, ZN => N2520);
   U1814 : AOI22_X1 port map( A1 => DATA2(2), A2 => n22599, B1 => n22598, B2 =>
                           n22934, ZN => N2519);
   U1815 : AOI22_X1 port map( A1 => DATA2(1), A2 => n22599, B1 => n22598, B2 =>
                           n22919, ZN => N2518);
   U1816 : AOI22_X1 port map( A1 => DATA2(0), A2 => n22599, B1 => n22598, B2 =>
                           n22597, ZN => N2517);
   U1817 : NOR2_X1 port map( A1 => n22600, A2 => n1796, ZN => n14253);
   U1818 : NAND2_X1 port map( A1 => n22639, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n22604);
   U1819 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , ZN => n22635);
   U1820 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n22635, ZN => n22634);
   U1821 : INV_X1 port map( A => n22601, ZN => n22602);
   U1822 : AOI22_X1 port map( A1 => n21214, A2 => n22637, B1 => n9084, B2 => 
                           n22631, ZN => n22603);
   U1823 : OAI221_X1 port map( B1 => n1796, B2 => n22604, C1 => n1796, C2 => 
                           n22634, A => n22603, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1824 : INV_X1 port map( A => n22604, ZN => n22636);
   U1825 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n22637, B1 => n21214, B2 => n22636, ZN => 
                           n22606);
   U1826 : NAND2_X1 port map( A1 => n9081, A2 => n22631, ZN => n22605);
   U1827 : OAI211_X1 port map( C1 => n1795, C2 => n22634, A => n22606, B => 
                           n22605, ZN => boothmul_pipelined_i_mux_out_1_4_port)
                           ;
   U1828 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n22636, B1 => n22637, B2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n22608);
   U1829 : NAND2_X1 port map( A1 => n22631, A2 => n9078, ZN => n22607);
   U1830 : OAI211_X1 port map( C1 => n22634, C2 => n1794, A => n22608, B => 
                           n22607, ZN => boothmul_pipelined_i_mux_out_1_5_port)
                           ;
   U1831 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n22610);
   U1832 : NAND2_X1 port map( A1 => n22631, A2 => n9075, ZN => n22609);
   U1833 : OAI211_X1 port map( C1 => n1793, C2 => n22634, A => n22610, B => 
                           n22609, ZN => boothmul_pipelined_i_mux_out_1_6_port)
                           ;
   U1834 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n22612);
   U1835 : NAND2_X1 port map( A1 => n22631, A2 => n9072, ZN => n22611);
   U1836 : OAI211_X1 port map( C1 => n1792, C2 => n22634, A => n22612, B => 
                           n22611, ZN => boothmul_pipelined_i_mux_out_1_7_port)
                           ;
   U1837 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n22614);
   U1838 : NAND2_X1 port map( A1 => n22631, A2 => n9069, ZN => n22613);
   U1839 : OAI211_X1 port map( C1 => n1790, C2 => n22634, A => n22614, B => 
                           n22613, ZN => boothmul_pipelined_i_mux_out_1_8_port)
                           ;
   U1840 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n22616);
   U1841 : NAND2_X1 port map( A1 => n22631, A2 => n9066, ZN => n22615);
   U1842 : OAI211_X1 port map( C1 => n1789, C2 => n22634, A => n22616, B => 
                           n22615, ZN => boothmul_pipelined_i_mux_out_1_9_port)
                           ;
   U1843 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n22618);
   U1844 : NAND2_X1 port map( A1 => n22631, A2 => n9063, ZN => n22617);
   U1845 : OAI211_X1 port map( C1 => n1788, C2 => n22634, A => n22618, B => 
                           n22617, ZN => boothmul_pipelined_i_mux_out_1_10_port
                           );
   U1846 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n22620);
   U1847 : NAND2_X1 port map( A1 => n22631, A2 => n9060, ZN => n22619);
   U1848 : OAI211_X1 port map( C1 => n1787, C2 => n22634, A => n22620, B => 
                           n22619, ZN => boothmul_pipelined_i_mux_out_1_11_port
                           );
   U1849 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n22622);
   U1850 : NAND2_X1 port map( A1 => n22631, A2 => n9057, ZN => n22621);
   U1851 : OAI211_X1 port map( C1 => n1786, C2 => n22634, A => n22622, B => 
                           n22621, ZN => boothmul_pipelined_i_mux_out_1_12_port
                           );
   U1852 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n22624);
   U1853 : NAND2_X1 port map( A1 => n22631, A2 => n9054, ZN => n22623);
   U1854 : OAI211_X1 port map( C1 => n1785, C2 => n22634, A => n22624, B => 
                           n22623, ZN => boothmul_pipelined_i_mux_out_1_13_port
                           );
   U1855 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n22626);
   U1856 : NAND2_X1 port map( A1 => n22631, A2 => n9051, ZN => n22625);
   U1857 : OAI211_X1 port map( C1 => n1784, C2 => n22634, A => n22626, B => 
                           n22625, ZN => boothmul_pipelined_i_mux_out_1_14_port
                           );
   U1858 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n22628);
   U1859 : NAND2_X1 port map( A1 => n22631, A2 => n9048, ZN => n22627);
   U1860 : OAI211_X1 port map( C1 => n1783, C2 => n22634, A => n22628, B => 
                           n22627, ZN => boothmul_pipelined_i_mux_out_1_15_port
                           );
   U1861 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n22630);
   U1862 : NAND2_X1 port map( A1 => n22631, A2 => n9045, ZN => n22629);
   U1863 : OAI211_X1 port map( C1 => n1782, C2 => n22634, A => n22630, B => 
                           n22629, ZN => boothmul_pipelined_i_mux_out_1_16_port
                           );
   U1864 : AOI22_X1 port map( A1 => n22637, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n22633);
   U1865 : NAND2_X1 port map( A1 => n22631, A2 => data1_mul_15_port, ZN => 
                           n22632);
   U1866 : OAI211_X1 port map( C1 => n1781, C2 => n22634, A => n22633, B => 
                           n22632, ZN => boothmul_pipelined_i_mux_out_1_17_port
                           );
   U1867 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n22635, ZN => 
                           n22640);
   U1868 : AOI22_X1 port map( A1 => n22637, A2 => n18051, B1 => n22636, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n22638);
   U1869 : OAI21_X1 port map( B1 => n22640, B2 => n22639, A => n22638, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1870 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n22927);
   U1871 : OR2_X1 port map( A1 => n22927, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n14252);
   U1872 : AOI22_X1 port map( A1 => n21214, A2 => n19413, B1 => n9084, B2 => 
                           n19200, ZN => n22641);
   U1873 : OAI221_X1 port map( B1 => n1796, B2 => n19365, C1 => n1796, C2 => 
                           n19252, A => n22641, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1874 : AOI22_X1 port map( A1 => n21214, A2 => n19145, B1 => n9081, B2 => 
                           n19200, ZN => n22643);
   U1875 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n19413, ZN => n22642);
   U1876 : OAI211_X1 port map( C1 => n19252, C2 => n1795, A => n22643, B => 
                           n22642, ZN => boothmul_pipelined_i_mux_out_2_6_port)
                           ;
   U1877 : AOI22_X1 port map( A1 => n9078, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n19413, ZN => n22645);
   U1878 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n19145, ZN => n22644);
   U1879 : OAI211_X1 port map( C1 => n19252, C2 => n1794, A => n22645, B => 
                           n22644, ZN => boothmul_pipelined_i_mux_out_2_7_port)
                           ;
   U1880 : AOI22_X1 port map( A1 => n9075, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n19413, ZN => n22647);
   U1881 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n19145, ZN => n22646);
   U1882 : OAI211_X1 port map( C1 => n19252, C2 => n1793, A => n22647, B => 
                           n22646, ZN => boothmul_pipelined_i_mux_out_2_8_port)
                           ;
   U1883 : AOI22_X1 port map( A1 => n9072, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n19413, ZN => n22649);
   U1884 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n19145, ZN => n22648);
   U1885 : OAI211_X1 port map( C1 => n19252, C2 => n1792, A => n22649, B => 
                           n22648, ZN => boothmul_pipelined_i_mux_out_2_9_port)
                           ;
   U1886 : AOI22_X1 port map( A1 => n9069, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n19413, ZN => n22651);
   U1887 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n19145, ZN => n22650);
   U1888 : OAI211_X1 port map( C1 => n19252, C2 => n1790, A => n22651, B => 
                           n22650, ZN => boothmul_pipelined_i_mux_out_2_10_port
                           );
   U1889 : AOI22_X1 port map( A1 => n9066, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n19413, ZN => n22653);
   U1890 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n19145, ZN => n22652);
   U1891 : OAI211_X1 port map( C1 => n19252, C2 => n1789, A => n22653, B => 
                           n22652, ZN => boothmul_pipelined_i_mux_out_2_11_port
                           );
   U1892 : AOI22_X1 port map( A1 => n9063, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n19413, ZN => n22655);
   U1893 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n19145, ZN => n22654);
   U1894 : OAI211_X1 port map( C1 => n19252, C2 => n1788, A => n22655, B => 
                           n22654, ZN => boothmul_pipelined_i_mux_out_2_12_port
                           );
   U1895 : AOI22_X1 port map( A1 => n9060, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n19413, ZN => n22657);
   U1896 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n19145, ZN => n22656);
   U1897 : OAI211_X1 port map( C1 => n19252, C2 => n1787, A => n22657, B => 
                           n22656, ZN => boothmul_pipelined_i_mux_out_2_13_port
                           );
   U1898 : AOI22_X1 port map( A1 => n9057, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n19413, ZN => n22659);
   U1899 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n19145, ZN => n22658);
   U1900 : OAI211_X1 port map( C1 => n19252, C2 => n1786, A => n22659, B => 
                           n22658, ZN => boothmul_pipelined_i_mux_out_2_14_port
                           );
   U1901 : AOI22_X1 port map( A1 => n9054, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n19413, ZN => n22661);
   U1902 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n19145, ZN => n22660);
   U1903 : OAI211_X1 port map( C1 => n19252, C2 => n1785, A => n22661, B => 
                           n22660, ZN => boothmul_pipelined_i_mux_out_2_15_port
                           );
   U1904 : AOI22_X1 port map( A1 => n9051, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n19413, ZN => n22663);
   U1905 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n19145, ZN => n22662);
   U1906 : OAI211_X1 port map( C1 => n19252, C2 => n1784, A => n22663, B => 
                           n22662, ZN => boothmul_pipelined_i_mux_out_2_16_port
                           );
   U1907 : AOI22_X1 port map( A1 => n9048, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n19413, ZN => n22665);
   U1908 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n19145, ZN => n22664);
   U1909 : OAI211_X1 port map( C1 => n19252, C2 => n1783, A => n22665, B => 
                           n22664, ZN => boothmul_pipelined_i_mux_out_2_17_port
                           );
   U1910 : AOI22_X1 port map( A1 => n9045, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n19413, ZN => n22667);
   U1911 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n19145, ZN => n22666);
   U1912 : OAI211_X1 port map( C1 => n19252, C2 => n1782, A => n22667, B => 
                           n22666, ZN => boothmul_pipelined_i_mux_out_2_18_port
                           );
   U1913 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n19200, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n19413, ZN => n22669);
   U1914 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n19145, ZN => n22668);
   U1915 : OAI211_X1 port map( C1 => n19252, C2 => n1781, A => n22669, B => 
                           n22668, ZN => boothmul_pipelined_i_mux_out_2_19_port
                           );
   U1916 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN 
                           => n22763);
   U1917 : OAI222_X1 port map( A1 => n22763, A2 => n19365, B1 => n1780, B2 => 
                           n19201, C1 => n19290, C2 => n22762, ZN => n13855);
   U1918 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4295, ZN => n22670);
   U1919 : NAND2_X1 port map( A1 => n7769, A2 => n22670, ZN => n14251);
   U1920 : AOI22_X1 port map( A1 => n21214, A2 => n19217, B1 => n9084, B2 => 
                           n19279, ZN => n22671);
   U1921 : OAI221_X1 port map( B1 => n1796, B2 => n19251, C1 => n1796, C2 => 
                           n19215, A => n22671, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1922 : OAI22_X1 port map( A1 => n19251, A2 => n21213, B1 => n19215, B2 => 
                           n1795, ZN => n22672);
   U1923 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           B2 => n19217, A => n22672, ZN => n22673);
   U1924 : OAI21_X1 port map( B1 => n19411, B2 => n1794, A => n22673, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1925 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN 
                           => n22841);
   U1926 : OAI22_X1 port map( A1 => n19215, A2 => n1794, B1 => n19411, B2 => 
                           n1793, ZN => n22674);
   U1927 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           B2 => n19217, A => n22674, ZN => n22675);
   U1928 : OAI21_X1 port map( B1 => n19251, B2 => n22841, A => n22675, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1929 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN 
                           => n22842);
   U1930 : OAI22_X1 port map( A1 => n19251, A2 => n22842, B1 => n19411, B2 => 
                           n1792, ZN => n22676);
   U1931 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           B2 => n19217, A => n22676, ZN => n22677);
   U1932 : OAI21_X1 port map( B1 => n19215, B2 => n1793, A => n22677, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1933 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN 
                           => n22843);
   U1934 : OAI22_X1 port map( A1 => n19251, A2 => n22843, B1 => n19411, B2 => 
                           n1790, ZN => n22678);
   U1935 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           B2 => n19217, A => n22678, ZN => n22679);
   U1936 : OAI21_X1 port map( B1 => n19215, B2 => n1792, A => n22679, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1937 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN 
                           => n22844);
   U1938 : OAI22_X1 port map( A1 => n19251, A2 => n22844, B1 => n19411, B2 => 
                           n1789, ZN => n22680);
   U1939 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           B2 => n19217, A => n22680, ZN => n22681);
   U1940 : OAI21_X1 port map( B1 => n19215, B2 => n1790, A => n22681, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1941 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN 
                           => n22845);
   U1942 : OAI22_X1 port map( A1 => n19251, A2 => n22845, B1 => n19411, B2 => 
                           n1788, ZN => n22682);
   U1943 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           B2 => n19217, A => n22682, ZN => n22683);
   U1944 : OAI21_X1 port map( B1 => n19215, B2 => n1789, A => n22683, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1945 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN 
                           => n22846);
   U1946 : OAI22_X1 port map( A1 => n19251, A2 => n22846, B1 => n19411, B2 => 
                           n1787, ZN => n22684);
   U1947 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           B2 => n19217, A => n22684, ZN => n22685);
   U1948 : OAI21_X1 port map( B1 => n19215, B2 => n1788, A => n22685, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U1949 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN 
                           => n22847);
   U1950 : OAI22_X1 port map( A1 => n19251, A2 => n22847, B1 => n19411, B2 => 
                           n1786, ZN => n22686);
   U1951 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           B2 => n19217, A => n22686, ZN => n22687);
   U1952 : OAI21_X1 port map( B1 => n19215, B2 => n1787, A => n22687, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U1953 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN 
                           => n22848);
   U1954 : OAI22_X1 port map( A1 => n19251, A2 => n22848, B1 => n19411, B2 => 
                           n1785, ZN => n22688);
   U1955 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           B2 => n19217, A => n22688, ZN => n22689);
   U1956 : OAI21_X1 port map( B1 => n19215, B2 => n1786, A => n22689, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U1957 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN 
                           => n22849);
   U1958 : OAI22_X1 port map( A1 => n19251, A2 => n22849, B1 => n19411, B2 => 
                           n1784, ZN => n22690);
   U1959 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           B2 => n19217, A => n22690, ZN => n22691);
   U1960 : OAI21_X1 port map( B1 => n19215, B2 => n1785, A => n22691, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U1961 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN 
                           => n22850);
   U1962 : OAI22_X1 port map( A1 => n19251, A2 => n22850, B1 => n19411, B2 => 
                           n1783, ZN => n22692);
   U1963 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           B2 => n19217, A => n22692, ZN => n22693);
   U1964 : OAI21_X1 port map( B1 => n19215, B2 => n1784, A => n22693, ZN => 
                           n14145);
   U1965 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN 
                           => n22851);
   U1966 : OAI22_X1 port map( A1 => n19251, A2 => n22851, B1 => n19411, B2 => 
                           n1782, ZN => n22694);
   U1967 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           B2 => n19217, A => n22694, ZN => n22695);
   U1968 : OAI21_X1 port map( B1 => n19215, B2 => n1783, A => n22695, ZN => 
                           n14144);
   U1969 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN 
                           => n22853);
   U1970 : OAI22_X1 port map( A1 => n19251, A2 => n22853, B1 => n19411, B2 => 
                           n1781, ZN => n22696);
   U1971 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           B2 => n19217, A => n22696, ZN => n22697);
   U1972 : OAI21_X1 port map( B1 => n19215, B2 => n1782, A => n22697, ZN => 
                           n14143);
   U1973 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN 
                           => n22855);
   U1974 : OAI22_X1 port map( A1 => n19251, A2 => n22855, B1 => n19411, B2 => 
                           n1780, ZN => n22698);
   U1975 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           B2 => n19217, A => n22698, ZN => n22699);
   U1976 : OAI21_X1 port map( B1 => n19215, B2 => n1781, A => n22699, ZN => 
                           n14142);
   U1977 : OAI222_X1 port map( A1 => n22763, A2 => n19251, B1 => n1780, B2 => 
                           n19278, C1 => n19358, C2 => n22762, ZN => n13854);
   U1978 : OR2_X1 port map( A1 => n4302, A2 => n22700, ZN => n14141);
   U1979 : AOI22_X1 port map( A1 => n21214, A2 => n19280, B1 => n9084, B2 => 
                           n19219, ZN => n22701);
   U1980 : OAI221_X1 port map( B1 => n1796, B2 => n19160, C1 => n1796, C2 => 
                           n19218, A => n22701, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U1981 : AOI22_X1 port map( A1 => n21214, A2 => n19410, B1 => n9081, B2 => 
                           n19219, ZN => n22703);
   U1982 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n19280, ZN => n22702);
   U1983 : OAI211_X1 port map( C1 => n19160, C2 => n1795, A => n22703, B => 
                           n22702, ZN => boothmul_pipelined_i_mux_out_4_10_port
                           );
   U1984 : AOI22_X1 port map( A1 => n9078, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n19280, ZN => n22705);
   U1985 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n19410, ZN => n22704);
   U1986 : OAI211_X1 port map( C1 => n19160, C2 => n1794, A => n22705, B => 
                           n22704, ZN => boothmul_pipelined_i_mux_out_4_11_port
                           );
   U1987 : AOI22_X1 port map( A1 => n9075, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n19280, ZN => n22707);
   U1988 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n19410, ZN => n22706);
   U1989 : OAI211_X1 port map( C1 => n19160, C2 => n1793, A => n22707, B => 
                           n22706, ZN => boothmul_pipelined_i_mux_out_4_12_port
                           );
   U1990 : AOI22_X1 port map( A1 => n9072, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n19280, ZN => n22709);
   U1991 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n19410, ZN => n22708);
   U1992 : OAI211_X1 port map( C1 => n19160, C2 => n1792, A => n22709, B => 
                           n22708, ZN => boothmul_pipelined_i_mux_out_4_13_port
                           );
   U1993 : AOI22_X1 port map( A1 => n9069, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n19280, ZN => n22711);
   U1994 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n19410, ZN => n22710);
   U1995 : OAI211_X1 port map( C1 => n19160, C2 => n1790, A => n22711, B => 
                           n22710, ZN => boothmul_pipelined_i_mux_out_4_14_port
                           );
   U1996 : AOI22_X1 port map( A1 => n9066, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n19280, ZN => n22713);
   U1997 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n19410, ZN => n22712);
   U1998 : OAI211_X1 port map( C1 => n19160, C2 => n1789, A => n22713, B => 
                           n22712, ZN => boothmul_pipelined_i_mux_out_4_15_port
                           );
   U1999 : AOI22_X1 port map( A1 => n9063, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n19280, ZN => n22715);
   U2000 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n19410, ZN => n22714);
   U2001 : OAI211_X1 port map( C1 => n19160, C2 => n1788, A => n22715, B => 
                           n22714, ZN => n8928);
   U2002 : AOI22_X1 port map( A1 => n9060, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n19280, ZN => n22717);
   U2003 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n19410, ZN => n22716);
   U2004 : OAI211_X1 port map( C1 => n19160, C2 => n1787, A => n22717, B => 
                           n22716, ZN => n13904);
   U2005 : AOI22_X1 port map( A1 => n9057, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n19280, ZN => n22719);
   U2006 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n19410, ZN => n22718);
   U2007 : OAI211_X1 port map( C1 => n19160, C2 => n1786, A => n22719, B => 
                           n22718, ZN => n13903);
   U2008 : AOI22_X1 port map( A1 => n9054, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n19280, ZN => n22721);
   U2009 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n19410, ZN => n22720);
   U2010 : OAI211_X1 port map( C1 => n19160, C2 => n1785, A => n22721, B => 
                           n22720, ZN => n13902);
   U2011 : AOI22_X1 port map( A1 => n9051, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n19280, ZN => n22723);
   U2012 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n19410, ZN => n22722);
   U2013 : OAI211_X1 port map( C1 => n19160, C2 => n1784, A => n22723, B => 
                           n22722, ZN => n13901);
   U2014 : AOI22_X1 port map( A1 => n9048, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n19280, ZN => n22725);
   U2015 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n19410, ZN => n22724);
   U2016 : OAI211_X1 port map( C1 => n19160, C2 => n1783, A => n22725, B => 
                           n22724, ZN => n13900);
   U2017 : AOI22_X1 port map( A1 => n9045, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n19280, ZN => n22727);
   U2018 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n19410, ZN => n22726);
   U2019 : OAI211_X1 port map( C1 => n19160, C2 => n1782, A => n22727, B => 
                           n22726, ZN => n13899);
   U2020 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n19219, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n19280, ZN => n22729);
   U2021 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n19410, ZN => n22728);
   U2022 : OAI211_X1 port map( C1 => n19160, C2 => n1781, A => n22729, B => 
                           n22728, ZN => n13898);
   U2023 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n19410, B1 => n19280, B2 => n18051, ZN => 
                           n22730);
   U2024 : OAI221_X1 port map( B1 => n1780, B2 => n19160, C1 => n1780, C2 => 
                           n19357, A => n22730, ZN => n13861);
   U2025 : NOR2_X1 port map( A1 => n4302, A2 => n14286, ZN => n22731);
   U2026 : NAND2_X1 port map( A1 => n14287, A2 => n22731, ZN => n17968);
   U2027 : AOI22_X1 port map( A1 => n21214, A2 => n19249, B1 => n9084, B2 => 
                           n19291, ZN => n22732);
   U2028 : OAI221_X1 port map( B1 => n1796, B2 => n19250, C1 => n1796, C2 => 
                           n19159, A => n22732, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2029 : OAI22_X1 port map( A1 => n19250, A2 => n21213, B1 => n19159, B2 => 
                           n1795, ZN => n22733);
   U2030 : AOI21_X1 port map( B1 => n9081, B2 => n19291, A => n22733, ZN => 
                           n22734);
   U2031 : OAI21_X1 port map( B1 => n19415, B2 => n22841, A => n22734, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2032 : OAI22_X1 port map( A1 => n19415, A2 => n22842, B1 => n19159, B2 => 
                           n1794, ZN => n22735);
   U2033 : AOI21_X1 port map( B1 => n9078, B2 => n19291, A => n22735, ZN => 
                           n22736);
   U2034 : OAI21_X1 port map( B1 => n19250, B2 => n22841, A => n22736, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2035 : OAI22_X1 port map( A1 => n19415, A2 => n22843, B1 => n19250, B2 => 
                           n22842, ZN => n22737);
   U2036 : AOI21_X1 port map( B1 => n9075, B2 => n19291, A => n22737, ZN => 
                           n22738);
   U2037 : OAI21_X1 port map( B1 => n19159, B2 => n1793, A => n22738, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2038 : OAI22_X1 port map( A1 => n19415, A2 => n22844, B1 => n19250, B2 => 
                           n22843, ZN => n22739);
   U2039 : AOI21_X1 port map( B1 => n9072, B2 => n19291, A => n22739, ZN => 
                           n22740);
   U2040 : OAI21_X1 port map( B1 => n19159, B2 => n1792, A => n22740, ZN => 
                           n14249);
   U2041 : OAI22_X1 port map( A1 => n19415, A2 => n22845, B1 => n19250, B2 => 
                           n22844, ZN => n22741);
   U2042 : AOI21_X1 port map( B1 => n9069, B2 => n19291, A => n22741, ZN => 
                           n22742);
   U2043 : OAI21_X1 port map( B1 => n19159, B2 => n1790, A => n22742, ZN => 
                           n14248);
   U2044 : OAI22_X1 port map( A1 => n19415, A2 => n22846, B1 => n19250, B2 => 
                           n22845, ZN => n22743);
   U2045 : AOI21_X1 port map( B1 => n9066, B2 => n19291, A => n22743, ZN => 
                           n22744);
   U2046 : OAI21_X1 port map( B1 => n19159, B2 => n1789, A => n22744, ZN => 
                           n14247);
   U2047 : OAI22_X1 port map( A1 => n19415, A2 => n22847, B1 => n19250, B2 => 
                           n22846, ZN => n22745);
   U2048 : AOI21_X1 port map( B1 => n9063, B2 => n19291, A => n22745, ZN => 
                           n22746);
   U2049 : OAI21_X1 port map( B1 => n19159, B2 => n1788, A => n22746, ZN => 
                           n14246);
   U2050 : OAI22_X1 port map( A1 => n19415, A2 => n22848, B1 => n19250, B2 => 
                           n22847, ZN => n22747);
   U2051 : AOI21_X1 port map( B1 => n9060, B2 => n19291, A => n22747, ZN => 
                           n22748);
   U2052 : OAI21_X1 port map( B1 => n19159, B2 => n1787, A => n22748, ZN => 
                           n14245);
   U2053 : OAI22_X1 port map( A1 => n19415, A2 => n22849, B1 => n19250, B2 => 
                           n22848, ZN => n22749);
   U2054 : AOI21_X1 port map( B1 => n9057, B2 => n19291, A => n22749, ZN => 
                           n22750);
   U2055 : OAI21_X1 port map( B1 => n19159, B2 => n1786, A => n22750, ZN => 
                           n14244);
   U2056 : OAI22_X1 port map( A1 => n19415, A2 => n22850, B1 => n19250, B2 => 
                           n22849, ZN => n22751);
   U2057 : AOI21_X1 port map( B1 => n9054, B2 => n19291, A => n22751, ZN => 
                           n22752);
   U2058 : OAI21_X1 port map( B1 => n19159, B2 => n1785, A => n22752, ZN => 
                           n14243);
   U2059 : OAI22_X1 port map( A1 => n19415, A2 => n22851, B1 => n19250, B2 => 
                           n22850, ZN => n22753);
   U2060 : AOI21_X1 port map( B1 => n9051, B2 => n19291, A => n22753, ZN => 
                           n22754);
   U2061 : OAI21_X1 port map( B1 => n19159, B2 => n1784, A => n22754, ZN => 
                           n14242);
   U2062 : OAI22_X1 port map( A1 => n19415, A2 => n22853, B1 => n19250, B2 => 
                           n22851, ZN => n22755);
   U2063 : AOI21_X1 port map( B1 => n9048, B2 => n19291, A => n22755, ZN => 
                           n22756);
   U2064 : OAI21_X1 port map( B1 => n19159, B2 => n1783, A => n22756, ZN => 
                           n14241);
   U2065 : OAI22_X1 port map( A1 => n19415, A2 => n22855, B1 => n19250, B2 => 
                           n22853, ZN => n22757);
   U2066 : AOI21_X1 port map( B1 => n9045, B2 => n19291, A => n22757, ZN => 
                           n22758);
   U2067 : OAI21_X1 port map( B1 => n19159, B2 => n1782, A => n22758, ZN => 
                           n14240);
   U2068 : OAI22_X1 port map( A1 => n19415, A2 => n22763, B1 => n19250, B2 => 
                           n22855, ZN => n22759);
   U2069 : AOI21_X1 port map( B1 => data1_mul_15_port, B2 => n19291, A => 
                           n22759, ZN => n22760);
   U2070 : OAI21_X1 port map( B1 => n19159, B2 => n1781, A => n22760, ZN => 
                           n13897);
   U2071 : NOR2_X1 port map( A1 => n14287, A2 => n22761, ZN => n21162);
   U2072 : NOR2_X1 port map( A1 => n14287, A2 => n17932, ZN => n17965);
   U2073 : NOR2_X1 port map( A1 => n17965, A2 => n21162, ZN => n17966);
   U2074 : OAI222_X1 port map( A1 => n22763, A2 => n19250, B1 => n1780, B2 => 
                           n19248, C1 => n19415, C2 => n22762, ZN => n13860);
   U2075 : NAND3_X1 port map( A1 => n21161, A2 => n19292, A3 => n21158, ZN => 
                           n22800);
   U2076 : NOR2_X1 port map( A1 => n19292, A2 => n21161, ZN => n22764);
   U2077 : NAND2_X1 port map( A1 => n22764, A2 => n19293, ZN => n22767);
   U2078 : AOI22_X1 port map( A1 => n21214, A2 => n22797, B1 => n9084, B2 => 
                           n22796, ZN => n22766);
   U2079 : OAI221_X1 port map( B1 => n1796, B2 => n22800, C1 => n1796, C2 => 
                           n22767, A => n22766, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2080 : INV_X1 port map( A => n22767, ZN => n22798);
   U2081 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n22797, B1 => n21214, B2 => n22798, ZN => 
                           n22769);
   U2082 : NAND2_X1 port map( A1 => n9081, A2 => n22796, ZN => n22768);
   U2083 : OAI211_X1 port map( C1 => n22800, C2 => n1795, A => n22769, B => 
                           n22768, ZN => boothmul_pipelined_i_mux_out_6_14_port
                           );
   U2084 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n22797, ZN => n22771);
   U2085 : NAND2_X1 port map( A1 => n9078, A2 => n22796, ZN => n22770);
   U2086 : OAI211_X1 port map( C1 => n22800, C2 => n1794, A => n22771, B => 
                           n22770, ZN => boothmul_pipelined_i_mux_out_6_15_port
                           );
   U2087 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n22797, ZN => n22773);
   U2088 : NAND2_X1 port map( A1 => n9075, A2 => n22796, ZN => n22772);
   U2089 : OAI211_X1 port map( C1 => n22800, C2 => n1793, A => n22773, B => 
                           n22772, ZN => boothmul_pipelined_i_mux_out_6_16_port
                           );
   U2090 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n22797, ZN => n22775);
   U2091 : NAND2_X1 port map( A1 => n9072, A2 => n22796, ZN => n22774);
   U2092 : OAI211_X1 port map( C1 => n22800, C2 => n1792, A => n22775, B => 
                           n22774, ZN => boothmul_pipelined_i_mux_out_6_17_port
                           );
   U2093 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n22797, ZN => n22777);
   U2094 : NAND2_X1 port map( A1 => n9069, A2 => n22796, ZN => n22776);
   U2095 : OAI211_X1 port map( C1 => n22800, C2 => n1790, A => n22777, B => 
                           n22776, ZN => boothmul_pipelined_i_mux_out_6_18_port
                           );
   U2096 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n22797, ZN => n22779);
   U2097 : NAND2_X1 port map( A1 => n9066, A2 => n22796, ZN => n22778);
   U2098 : OAI211_X1 port map( C1 => n22800, C2 => n1789, A => n22779, B => 
                           n22778, ZN => boothmul_pipelined_i_mux_out_6_19_port
                           );
   U2099 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n22797, ZN => n22781);
   U2100 : NAND2_X1 port map( A1 => n9063, A2 => n22796, ZN => n22780);
   U2101 : OAI211_X1 port map( C1 => n22800, C2 => n1788, A => n22781, B => 
                           n22780, ZN => boothmul_pipelined_i_mux_out_6_20_port
                           );
   U2102 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n22797, ZN => n22783);
   U2103 : NAND2_X1 port map( A1 => n9060, A2 => n22796, ZN => n22782);
   U2104 : OAI211_X1 port map( C1 => n22800, C2 => n1787, A => n22783, B => 
                           n22782, ZN => boothmul_pipelined_i_mux_out_6_21_port
                           );
   U2105 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n22797, ZN => n22785);
   U2106 : NAND2_X1 port map( A1 => n9057, A2 => n22796, ZN => n22784);
   U2107 : OAI211_X1 port map( C1 => n22800, C2 => n1786, A => n22785, B => 
                           n22784, ZN => boothmul_pipelined_i_mux_out_6_22_port
                           );
   U2108 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n22797, ZN => n22787);
   U2109 : NAND2_X1 port map( A1 => n9054, A2 => n22796, ZN => n22786);
   U2110 : OAI211_X1 port map( C1 => n22800, C2 => n1785, A => n22787, B => 
                           n22786, ZN => boothmul_pipelined_i_mux_out_6_23_port
                           );
   U2111 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n22797, ZN => n22789);
   U2112 : NAND2_X1 port map( A1 => n9051, A2 => n22796, ZN => n22788);
   U2113 : OAI211_X1 port map( C1 => n22800, C2 => n1784, A => n22789, B => 
                           n22788, ZN => boothmul_pipelined_i_mux_out_6_24_port
                           );
   U2114 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n22797, ZN => n22791);
   U2115 : NAND2_X1 port map( A1 => n9048, A2 => n22796, ZN => n22790);
   U2116 : OAI211_X1 port map( C1 => n22800, C2 => n1783, A => n22791, B => 
                           n22790, ZN => n14239);
   U2117 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n22797, ZN => n22793);
   U2118 : NAND2_X1 port map( A1 => n9045, A2 => n22796, ZN => n22792);
   U2119 : OAI211_X1 port map( C1 => n22800, C2 => n1782, A => n22793, B => 
                           n22792, ZN => n14238);
   U2120 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n22798, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n22797, ZN => n22795);
   U2121 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n22796, ZN => 
                           n22794);
   U2122 : OAI211_X1 port map( C1 => n22800, C2 => n1781, A => n22795, B => 
                           n22794, ZN => n13896);
   U2123 : INV_X1 port map( A => n22796, ZN => n22801);
   U2124 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n22798, B1 => n22797, B2 => n18051, ZN => 
                           n22799);
   U2125 : OAI221_X1 port map( B1 => n1780, B2 => n22801, C1 => n1780, C2 => 
                           n22800, A => n22799, ZN => n13859);
   U2126 : NAND3_X1 port map( A1 => n21166, A2 => n21159, A3 => n19294, ZN => 
                           n22805);
   U2127 : INV_X1 port map( A => n22837, ZN => n22804);
   U2128 : AOI22_X1 port map( A1 => n22835, A2 => n19349, B1 => n22836, B2 => 
                           n19369, ZN => n22803);
   U2129 : OAI221_X1 port map( B1 => n19440, B2 => n22805, C1 => n19440, C2 => 
                           n22804, A => n22803, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2130 : INV_X1 port map( A => n22805, ZN => n22834);
   U2131 : AOI22_X1 port map( A1 => n19349, A2 => n22834, B1 => n22837, B2 => 
                           n19369, ZN => n22807);
   U2132 : AOI22_X1 port map( A1 => n22835, A2 => n19348, B1 => n22836, B2 => 
                           n19370, ZN => n22806);
   U2133 : NAND2_X1 port map( A1 => n22807, A2 => n22806, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2134 : AOI22_X1 port map( A1 => n22834, A2 => n19348, B1 => n22837, B2 => 
                           n19370, ZN => n22809);
   U2135 : AOI22_X1 port map( A1 => n22835, A2 => n19347, B1 => n22836, B2 => 
                           n19371, ZN => n22808);
   U2136 : NAND2_X1 port map( A1 => n22809, A2 => n22808, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2137 : AOI22_X1 port map( A1 => n22834, A2 => n19347, B1 => n22837, B2 => 
                           n19371, ZN => n22811);
   U2138 : AOI22_X1 port map( A1 => n22835, A2 => n19346, B1 => n22836, B2 => 
                           n19372, ZN => n22810);
   U2139 : NAND2_X1 port map( A1 => n22811, A2 => n22810, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2140 : AOI22_X1 port map( A1 => n22834, A2 => n19346, B1 => n22837, B2 => 
                           n19372, ZN => n22813);
   U2141 : AOI22_X1 port map( A1 => n22835, A2 => n19345, B1 => n22836, B2 => 
                           n19373, ZN => n22812);
   U2142 : NAND2_X1 port map( A1 => n22813, A2 => n22812, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2143 : AOI22_X1 port map( A1 => n22834, A2 => n19345, B1 => n22837, B2 => 
                           n19373, ZN => n22815);
   U2144 : AOI22_X1 port map( A1 => n22835, A2 => n19344, B1 => n22836, B2 => 
                           n19374, ZN => n22814);
   U2145 : NAND2_X1 port map( A1 => n22815, A2 => n22814, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2146 : AOI22_X1 port map( A1 => n22834, A2 => n19344, B1 => n22837, B2 => 
                           n19374, ZN => n22817);
   U2147 : AOI22_X1 port map( A1 => n22835, A2 => n19343, B1 => n22836, B2 => 
                           n19375, ZN => n22816);
   U2148 : NAND2_X1 port map( A1 => n22817, A2 => n22816, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2149 : AOI22_X1 port map( A1 => n22834, A2 => n19343, B1 => n22837, B2 => 
                           n19375, ZN => n22819);
   U2150 : AOI22_X1 port map( A1 => n22835, A2 => n19342, B1 => n22836, B2 => 
                           n19376, ZN => n22818);
   U2151 : NAND2_X1 port map( A1 => n22819, A2 => n22818, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2152 : AOI22_X1 port map( A1 => n22834, A2 => n19342, B1 => n22837, B2 => 
                           n19376, ZN => n22821);
   U2153 : AOI22_X1 port map( A1 => n22835, A2 => n19341, B1 => n22836, B2 => 
                           n19377, ZN => n22820);
   U2154 : NAND2_X1 port map( A1 => n22821, A2 => n22820, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2155 : AOI22_X1 port map( A1 => n22834, A2 => n19341, B1 => n22837, B2 => 
                           n19377, ZN => n22823);
   U2156 : AOI22_X1 port map( A1 => n22835, A2 => n19340, B1 => n22836, B2 => 
                           n19378, ZN => n22822);
   U2157 : NAND2_X1 port map( A1 => n22823, A2 => n22822, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2158 : AOI22_X1 port map( A1 => n22834, A2 => n19340, B1 => n22837, B2 => 
                           n19378, ZN => n22825);
   U2159 : AOI22_X1 port map( A1 => n22835, A2 => n19339, B1 => n22836, B2 => 
                           n19379, ZN => n22824);
   U2160 : NAND2_X1 port map( A1 => n22825, A2 => n22824, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2161 : AOI22_X1 port map( A1 => n22834, A2 => n19339, B1 => n22837, B2 => 
                           n19379, ZN => n22827);
   U2162 : AOI22_X1 port map( A1 => n22835, A2 => n19338, B1 => n22836, B2 => 
                           n19380, ZN => n22826);
   U2163 : NAND2_X1 port map( A1 => n22827, A2 => n22826, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2164 : AOI22_X1 port map( A1 => n22834, A2 => n19338, B1 => n22837, B2 => 
                           n19380, ZN => n22829);
   U2165 : AOI22_X1 port map( A1 => n22835, A2 => n19337, B1 => n22836, B2 => 
                           n19381, ZN => n22828);
   U2166 : NAND2_X1 port map( A1 => n22829, A2 => n22828, ZN => n14237);
   U2167 : AOI22_X1 port map( A1 => n22834, A2 => n19337, B1 => n22837, B2 => 
                           n19381, ZN => n22831);
   U2168 : AOI22_X1 port map( A1 => n22835, A2 => n19336, B1 => n22836, B2 => 
                           n19382, ZN => n22830);
   U2169 : NAND2_X1 port map( A1 => n22831, A2 => n22830, ZN => n14236);
   U2170 : AOI22_X1 port map( A1 => n22834, A2 => n19336, B1 => n22837, B2 => 
                           n19382, ZN => n22833);
   U2171 : AOI22_X1 port map( A1 => n22835, A2 => n21181, B1 => n22836, B2 => 
                           n19383, ZN => n22832);
   U2172 : NAND2_X1 port map( A1 => n22833, A2 => n22832, ZN => n14235);
   U2173 : OAI21_X1 port map( B1 => n22835, B2 => n22834, A => n21181, ZN => 
                           n22839);
   U2174 : AOI22_X1 port map( A1 => n22837, A2 => n19383, B1 => n22836, B2 => 
                           n19352, ZN => n22838);
   U2175 : NAND2_X1 port map( A1 => n22839, A2 => n22838, ZN => n14234);
   U2176 : INV_X1 port map( A => n22840, ZN => n22860);
   U2177 : OAI222_X1 port map( A1 => n1796, A2 => n22852, B1 => n21213, B2 => 
                           n22854, C1 => n22860, C2 => n1795, ZN => n13848);
   U2178 : OAI222_X1 port map( A1 => n22841, A2 => n22852, B1 => n22842, B2 => 
                           n22854, C1 => n1793, C2 => n22860, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2179 : OAI222_X1 port map( A1 => n1792, A2 => n22860, B1 => n22843, B2 => 
                           n22854, C1 => n22842, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2180 : OAI222_X1 port map( A1 => n1790, A2 => n22860, B1 => n22844, B2 => 
                           n22854, C1 => n22843, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2181 : OAI222_X1 port map( A1 => n1789, A2 => n22860, B1 => n22845, B2 => 
                           n22854, C1 => n22844, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2182 : OAI222_X1 port map( A1 => n1788, A2 => n22860, B1 => n22846, B2 => 
                           n22854, C1 => n22845, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2183 : OAI222_X1 port map( A1 => n1787, A2 => n22860, B1 => n22847, B2 => 
                           n22854, C1 => n22846, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2184 : OAI222_X1 port map( A1 => n1786, A2 => n22860, B1 => n22848, B2 => 
                           n22854, C1 => n22847, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2185 : OAI222_X1 port map( A1 => n1785, A2 => n22860, B1 => n22849, B2 => 
                           n22854, C1 => n22848, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2186 : OAI222_X1 port map( A1 => n1784, A2 => n22860, B1 => n22850, B2 => 
                           n22854, C1 => n22849, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2187 : OAI222_X1 port map( A1 => n1783, A2 => n22860, B1 => n22851, B2 => 
                           n22854, C1 => n22850, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2188 : OAI222_X1 port map( A1 => n1782, A2 => n22860, B1 => n22853, B2 => 
                           n22854, C1 => n22851, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2189 : OAI222_X1 port map( A1 => n1781, A2 => n22860, B1 => n22855, B2 => 
                           n22854, C1 => n22853, C2 => n22852, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2190 : AOI22_X1 port map( A1 => n22858, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n22857, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n22856);
   U2191 : OAI21_X1 port map( B1 => n22860, B2 => n1780, A => n22856, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2192 : AOI22_X1 port map( A1 => n22858, A2 => n18051, B1 => n22857, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n22859);
   U2193 : OAI21_X1 port map( B1 => n22860, B2 => n1780, A => n22859, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U2194 : XNOR2_X1 port map( A => n22862, B => n22861, ZN => n14140);
   U2195 : INV_X1 port map( A => n22863, ZN => n22867);
   U2196 : OAI22_X1 port map( A1 => n22867, A2 => n22866, B1 => n22865, B2 => 
                           n22864, ZN => n22871);
   U2197 : OAI22_X1 port map( A1 => n22874, A2 => n22869, B1 => n22868, B2 => 
                           n22948, ZN => n22870);
   U2198 : AOI211_X1 port map( C1 => n22873, C2 => n22872, A => n22871, B => 
                           n22870, ZN => n1871);
   U2199 : NOR2_X1 port map( A1 => n1814, A2 => n22874, ZN => n22888);
   U2200 : OAI22_X1 port map( A1 => n22878, A2 => n22877, B1 => n22876, B2 => 
                           n22875, ZN => n22879);
   U2201 : AOI22_X1 port map( A1 => n22880, A2 => n22879, B1 => n22998, B2 => 
                           n18867, ZN => n22884);
   U2202 : OAI221_X1 port map( B1 => n22882, B2 => n22881, C1 => n22882, C2 => 
                           n19298, A => DATA2(6), ZN => n22883);
   U2203 : OAI211_X1 port map( C1 => n22958, C2 => n22885, A => n22884, B => 
                           n22883, ZN => n22886);
   U2204 : AOI21_X1 port map( B1 => n22888, B2 => n22887, A => n22886, ZN => 
                           n18133);
   U2205 : OAI22_X1 port map( A1 => n19394, A2 => n22890, B1 => n19212, B2 => 
                           n22889, ZN => n22891);
   U2206 : INV_X1 port map( A => n22891, ZN => n22892);
   U2207 : OAI211_X1 port map( C1 => n22892, C2 => n22983, A => n18882, B => 
                           n19270, ZN => OUTALU(6));
   U2208 : INV_X1 port map( A => n22893, ZN => n22895);
   U2209 : AOI22_X1 port map( A1 => n1835, A2 => n22894, B1 => n1894, B2 => 
                           n22895, ZN => n14432);
   U2210 : AOI22_X1 port map( A1 => n1843, A2 => n22896, B1 => n13151, B2 => 
                           n22895, ZN => n14431);
   U2211 : NOR3_X1 port map( A1 => n22899, A2 => n22898, A3 => n22897, ZN => 
                           n22906);
   U2212 : AOI221_X1 port map( B1 => n22904, B2 => n22903, C1 => n22902, C2 => 
                           n22901, A => n22900, ZN => n22905);
   U2213 : AOI211_X1 port map( C1 => n22908, C2 => n22907, A => n22906, B => 
                           n22905, ZN => n14416);
   U2214 : AOI22_X1 port map( A1 => n22912, A2 => n22911, B1 => n22910, B2 => 
                           n22909, ZN => n14452);
   U2215 : NAND2_X1 port map( A1 => n22915, A2 => n18195, ZN => n21157);
   U2216 : NAND4_X1 port map( A1 => DATA2(2), A2 => DATA2(4), A3 => n22922, A4 
                           => n22933, ZN => n21160);
   U2217 : OR2_X1 port map( A1 => n1798, A2 => n4302, ZN => n21163);
   U2218 : NOR2_X1 port map( A1 => n22913, A2 => n22920, ZN => n22921);
   U2219 : NAND3_X1 port map( A1 => DATA2(2), A2 => n22921, A3 => n22933, ZN =>
                           n21170);
   U2220 : NAND4_X1 port map( A1 => n22922, A2 => n22934, A3 => n22933, A4 => 
                           n1834, ZN => n21171);
   U2221 : NAND2_X1 port map( A1 => DATA2(4), A2 => DATA2(2), ZN => n22914);
   U2222 : NOR4_X1 port map( A1 => DATA2(3), A2 => DATA2(0), A3 => n22919, A4 
                           => n22914, ZN => n21172);
   U2223 : NOR2_X1 port map( A1 => DATA2(2), A2 => DATA2(1), ZN => n22932);
   U2224 : NOR4_X1 port map( A1 => n22915, A2 => n22932, A3 => n22921, A4 => 
                           n1840, ZN => n21174);
   U2225 : NAND3_X1 port map( A1 => DATA2(2), A2 => n22929, A3 => n22922, ZN =>
                           n21175);
   U2226 : INV_X1 port map( A => n22918, ZN => n22916);
   U2227 : NAND2_X1 port map( A1 => n22917, A2 => n22916, ZN => n21176);
   U2228 : NOR2_X1 port map( A1 => n22919, A2 => n22918, ZN => n21177);
   U2229 : NOR3_X1 port map( A1 => DATA2(2), A2 => n22920, A3 => n22931, ZN => 
                           n21178);
   U2230 : NAND3_X1 port map( A1 => n22921, A2 => n22934, A3 => n22933, ZN => 
                           n21179);
   U2231 : NAND2_X1 port map( A1 => n22922, A2 => n22934, ZN => n22923);
   U2232 : NOR2_X1 port map( A1 => n22931, A2 => n22923, ZN => n21180);
   U2233 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n22924);
   U2234 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n22924, ZN => n21183);
   U2235 : INV_X1 port map( A => n1800, ZN => n22925);
   U2236 : NAND2_X1 port map( A1 => n7769, A2 => n22925, ZN => n21186);
   U2237 : NOR3_X1 port map( A1 => n7769, A2 => n8978, A3 => n22926, ZN => 
                           n21187);
   U2238 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n22927, ZN => n14132);
   U2239 : NOR2_X1 port map( A1 => n22928, A2 => n14132, ZN => n21188);
   U2240 : OAI21_X1 port map( B1 => DATA2(2), B2 => n22930, A => n22929, ZN => 
                           n1847);
   U2241 : NOR2_X1 port map( A1 => n22932, A2 => n22931, ZN => n1845);
   U2242 : NAND2_X1 port map( A1 => n22934, A2 => n22933, ZN => n22935);
   U2243 : OAI21_X1 port map( B1 => n22936, B2 => n22935, A => n1834, ZN => 
                           n1844);
   U2244 : INV_X1 port map( A => n14407, ZN => n22937);
   U2245 : AOI22_X1 port map( A1 => n13151, A2 => n22937, B1 => n1894, B2 => 
                           n1826, ZN => n1827);
   U2246 : AOI22_X1 port map( A1 => n22941, A2 => n22940, B1 => n22939, B2 => 
                           n22938, ZN => n22947);
   U2247 : AOI22_X1 port map( A1 => n22945, A2 => n22944, B1 => n22943, B2 => 
                           n22942, ZN => n22946);
   U2248 : OAI211_X1 port map( C1 => n22949, C2 => n22948, A => n22947, B => 
                           n22946, ZN => n1822);
   U2249 : INV_X1 port map( A => n14003, ZN => n22951);
   U2250 : OAI22_X1 port map( A1 => n22951, A2 => n22997, B1 => n22950, B2 => 
                           n1836, ZN => n1820);
   U2251 : AOI22_X1 port map( A1 => n13151, A2 => n1826, B1 => n22953, B2 => 
                           n22952, ZN => n1818);
   U2252 : NOR2_X1 port map( A1 => n22955, A2 => n22954, ZN => n22957);
   U2253 : NAND2_X1 port map( A1 => n22998, A2 => n19055, ZN => n22956);
   U2254 : OAI21_X1 port map( B1 => n22958, B2 => n22957, A => n22956, ZN => 
                           n1812);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n30042, n30044, n30046, n30048, n30053, n30054, n30055, n30056, 
      n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, 
      n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, 
      n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, 
      n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, 
      n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, 
      n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, 
      n30112, n30113, n30115, n30116, n30117, n30118, n30120, n30121, n30123, 
      n30124, n31164, n31166, n31167, n31168, n31169, n31170, n31171, n35769, 
      n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, 
      n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, 
      n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, 
      n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, 
      n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, 
      n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, 
      n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, 
      n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, 
      n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, 
      n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, 
      n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, 
      n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, 
      n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, 
      n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, 
      n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, 
      n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, 
      n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, 
      n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, 
      n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, 
      n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, 
      n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, 
      n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, 
      n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, 
      n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, 
      n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, 
      n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, 
      n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, 
      n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, 
      n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, 
      n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, 
      n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, 
      n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, 
      n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, 
      n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, 
      n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, 
      n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, 
      n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, 
      n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, 
      n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, 
      n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, 
      n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, 
      n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, 
      n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, 
      n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, 
      n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, 
      n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, 
      n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, 
      n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, 
      n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, 
      n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, 
      n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, 
      n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, 
      n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, 
      n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, 
      n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, 
      n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, 
      n36275, n36276, n36277, n36278, n36279, n36281, n36283, n36284, n36285, 
      n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, 
      n36295, n36297, n36298, n36299, n36300, n36301, n36302, n36304, n36305, 
      n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, 
      n36316, n36317, n36318, n36319, n36320, n36322, n36323, n36324, n36325, 
      n36326, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, 
      n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, 
      n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, 
      n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, 
      n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, 
      n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, 
      n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, 
      n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36399, 
      n36400, n36401, n36402, n36404, n36405, n36406, n36407, n36408, n36409, 
      n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, 
      n36419, n36421, n36423, n36424, n36426, n36428, n36430, n36432, n36434, 
      n36435, n36436, n36437, n36438, n36439, n36440, n36442, n36443, n36444, 
      n36445, n36446, n36447, n36448, n36450, n36451, n36452, n36453, n36455, 
      n36456, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, 
      n36466, n36467, n36468, n36470, n36471, n36473, n36474, n36475, n36476, 
      n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36486, n36488, 
      n36490, n36491, n36492, n36494, n36495, n36496, n36497, n36498, n36499, 
      n36500, n36501, n36502, n36504, n36506, n36507, n36509, n36510, n36512, 
      n36513, n36516, n36517, n36518, n36520, n36521, n36523, n36524, n36526, 
      n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36536, 
      n36537, n36539, n36540, n36541, n36542, n36544, n36545, n36546, n36547, 
      n36548, n36549, n36551, n36552, n36553, n36554, n36555, n36556, n36557, 
      n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, 
      n36567, n36568, n36569, n36570, n36571, n36573, n36574, n36575, n36576, 
      n36577, n36578, n36580, n36581, n36582, n36583, n36585, n36587, n36588, 
      n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, 
      n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36607, 
      n36608, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, 
      n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, 
      n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, 
      n36637, n36639, n36640, n36641, n36642, n36644, n36645, n36646, n36647, 
      n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, 
      n36657, n36658, n36659, n36660, n36661, n36663, n36664, n36665, n36666, 
      n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36675, n36678, 
      n36679, n36680, n36681, n36682, n36684, n36685, n36686, n36688, n36689, 
      n36690, n36691, n36693, n36695, n36697, n36699, n36702, n36704, n36706, 
      n36707, n36709, n36711, n36713, n36716, n36719, n36720, n36721, n36722, 
      n36723, n36724, n36725, n36727, n36728, n36729, n36731, n36732, n36733, 
      n36734, n36735, n36737, n36738, n36739, n36740, n36741, n36742, n36743, 
      n36744, n36745, n36746, n36747, n36749, n36750, n36752, n36753, n36754, 
      n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, 
      n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, 
      n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, 
      n36782, n36784, n36785, n36786, n36787, n36789, n36790, n36791, n36792, 
      n36793, n36794, n36795, n36796, n36797, n36798, n36800, n36802, n36804, 
      n36806, n36808, n36809, n36810, n36812, n36814, n36815, n36816, n36817, 
      n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, 
      n36827, n36828, n36829, n36830, n36831, n36832, n36834, n36836, n36837, 
      n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, 
      n36847, n36848, n36849, n36850, n36852, n36853, n36854, n36856, n36858, 
      n36859, n36860, n36861, n36862, n36864, n36865, n36867, n36868, n36869, 
      n36871, n36873, n36874, n36876, n36877, n36879, n36881, n36883, n36885, 
      n36886, n36888, n36890, n36893, n36895, n36897, n40552, n40553, n40554, 
      n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, 
      n40565, n40568, n40571, n40574, n40576, n40577, n40580, n40581, n40582, 
      n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40591, n40592, 
      n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612, 
      n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620, n40621, 
      n40622, n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630, 
      n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639, 
      n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648, 
      n40649, n40654, n40655, n40656, n40657, n40658, n40660, n40662, n40663, 
      n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672, 
      n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681, 
      n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690, 
      n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699, 
      n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708, 
      n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717, 
      n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726, 
      n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735, 
      n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744, 
      n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753, 
      n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762, 
      n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771, 
      n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780, 
      n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789, 
      n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798, 
      n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807, 
      n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816, 
      n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825, 
      n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834, 
      n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843, 
      n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852, 
      n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861, 
      n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870, 
      n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879, 
      n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888, 
      n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897, 
      n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906, 
      n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915, 
      n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924, 
      n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933, 
      n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942, 
      n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951, 
      n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960, 
      n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969, 
      n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978, 
      n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987, 
      n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996, 
      n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005, 
      n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014, 
      n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023, 
      n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032, 
      n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041, 
      n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050, 
      n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059, 
      n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068, 
      n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077, 
      n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086, 
      n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095, 
      n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104, 
      n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113, 
      n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122, 
      n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131, 
      n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140, 
      n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149, 
      n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158, 
      n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, 
      n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, 
      n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185, 
      n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194, 
      n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203, 
      n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212, 
      n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221, 
      n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230, 
      n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239, 
      n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248, 
      n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257, 
      n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266, 
      n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275, 
      n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, 
      n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293, 
      n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302, 
      n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311, 
      n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320, 
      n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329, 
      n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338, 
      n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347, 
      n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356, 
      n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365, 
      n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374, 
      n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383, 
      n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392, 
      n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401, 
      n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410, 
      n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419, 
      n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428, 
      n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437, 
      n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446, 
      n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455, 
      n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464, 
      n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473, 
      n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482, 
      n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491, 
      n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500, 
      n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509, 
      n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518, 
      n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527, 
      n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536, 
      n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545, 
      n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554, 
      n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563, 
      n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572, 
      n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581, 
      n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590, 
      n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599, 
      n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608, 
      n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617, 
      n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626, 
      n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635, 
      n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644, 
      n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, 
      n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, 
      n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, 
      n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, 
      n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689, 
      n41690, n41691, n41692, n41693, n41694, n41697, n41698, n41699, n41700, 
      n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709, 
      n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718, 
      n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727, 
      n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736, 
      n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, 
      n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, 
      n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, 
      n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772, 
      n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780, n41781, 
      n41782, n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790, 
      n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799, 
      n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808, 
      n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817, 
      n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826, 
      n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835, 
      n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844, 
      n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852, n41853, 
      n41854, n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862, 
      n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871, 
      n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880, 
      n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889, 
      n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898, 
      n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907, 
      n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916, 
      n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924, n41925, 
      n41926, n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934, 
      n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943, 
      n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952, 
      n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961, 
      n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970, 
      n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979, 
      n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988, 
      n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996, n41997, 
      n41998, n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006, 
      n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014, n42015, 
      n42016, n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024, 
      n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033, 
      n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042, 
      n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051, 
      n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060, 
      n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068, n42069, 
      n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078, 
      n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086, n42087, 
      n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096, 
      n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105, 
      n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114, 
      n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123, 
      n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132, 
      n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141, 
      n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150, 
      n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158, n42159, 
      n42160, n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168, 
      n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177, 
      n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186, 
      n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195, 
      n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204, 
      n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212, n42213, 
      n42214, n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222, 
      n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230, n42231, 
      n42232, n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240, 
      n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249, 
      n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258, 
      n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267, 
      n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276, 
      n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285, 
      n42286, n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294, 
      n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302, n42303, 
      n42304, n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312, 
      n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321, 
      n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330, 
      n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339, 
      n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348, 
      n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356, n42357, 
      n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366, 
      n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374, n42375, 
      n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384, 
      n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393, 
      n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402, 
      n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411, 
      n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420, 
      n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429, 
      n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438, 
      n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446, n42447, 
      n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456, 
      n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465, 
      n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474, 
      n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483, 
      n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492, 
      n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501, 
      n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510, 
      n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518, n42519, 
      n42520, n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528, 
      n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537, 
      n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546, 
      n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555, 
      n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564, 
      n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573, 
      n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582, 
      n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591, 
      n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600, 
      n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609, 
      n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618, 
      n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627, 
      n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636, 
      n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645, 
      n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654, 
      n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663, 
      n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, 
      n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, 
      n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690, 
      n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699, 
      n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708, 
      n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717, 
      n42718, n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726, 
      n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735, 
      n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744, 
      n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753, 
      n42754, n42755, n42756, n42757, n42758, n42760, n47428, n47429, n47430, 
      n47431, n47432, n47446, n47447, n47449, n47453, n47493, n47494, n47495, 
      n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504, 
      n47505, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514, 
      n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523, 
      n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531, n47532, 
      n47533, n47534, n47535, n47536, n47537, n47538, n47539, n47540, n47541, 
      n47542, n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550, 
      n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558, n47559, 
      n47560, n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568, 
      n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577, 
      n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586, 
      n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595, 
      n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603, n47604, 
      n47605, n47606, n47607, n47608, n47609, n47610, n47611, n47612, n47613, 
      n47614, n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622, 
      n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630, n47631, 
      n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640, 
      n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649, 
      n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658, 
      n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667, 
      n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676, 
      n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47685, 
      n47686, n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694, 
      n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702, n47703, 
      n47704, n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712, 
      n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721, 
      n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730, 
      n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739, 
      n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747, n47748, 
      n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756, n47757, 
      n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766, 
      n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774, n47775, 
      n47776, n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784, 
      n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793, 
      n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802, 
      n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811, 
      n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819, n47820, 
      n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828, n47829, 
      n47830, n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838, 
      n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846, n47847, 
      n47848, n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856, 
      n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865, 
      n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874, 
      n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883, 
      n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891, n47892, 
      n47893, n47894, n47895, n47896, n47897, n47898, n47899, n47900, n47901, 
      n47902, n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910, 
      n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919, 
      n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928, 
      n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937, 
      n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946, 
      n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955, 
      n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964, 
      n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973, 
      n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982, 
      n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991, 
      n47992, n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000, 
      n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009, 
      n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018, 
      n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027, 
      n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036, 
      n48037, n48038, n48039, n48040, n48041, n48042, n48043, n48044, n48045, 
      n48046, n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054, 
      n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062, n48063, 
      n48064, n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072, 
      n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081, 
      n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090, 
      n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099, 
      n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108, 
      n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48116, n48117, 
      n48118, n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126, 
      n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135, 
      n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144, 
      n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153, 
      n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162, 
      n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171, 
      n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179, n48180, 
      n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188, n48189, 
      n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198, 
      n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206, n48207, 
      n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216, 
      n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225, 
      n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234, 
      n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243, 
      n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252, 
      n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261, 
      n48262, n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270, 
      n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279, 
      n48280, n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288, 
      n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297, 
      n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306, 
      n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315, 
      n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323, n48324, 
      n48325, n48326, n48327, n48328, n48329, n48330, n48331, n48332, n48333, 
      n48334, n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342, 
      n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350, n48351, 
      n48352, n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360, 
      n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369, 
      n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378, 
      n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387, 
      n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396, 
      n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404, n48405, 
      n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414, 
      n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422, n48423, 
      n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432, 
      n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440, n48441, 
      n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450, 
      n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459, 
      n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468, 
      n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477, 
      n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486, 
      n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495, 
      n48496, n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504, 
      n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513, 
      n48514, n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522, 
      n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531, 
      n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539, n48540, 
      n48541, n48542, n48543, n48544, n48545, n48546, n48547, n48548, n48549, 
      n48550, n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558, 
      n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567, 
      n48568, n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576, 
      n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584, n48585, 
      n48586, n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594, 
      n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603, 
      n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611, n48612, 
      n48613, n48614, n48615, n48616, n48617, n48618, n48619, n48620, n48621, 
      n48622, n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630, 
      n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638, n48639, 
      n48640, n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648, 
      n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656, n48657, 
      n48658, n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666, 
      n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675, 
      n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683, n48684, 
      n48685, n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693, 
      n48694, n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702, 
      n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710, n48711, 
      n48712, n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720, 
      n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728, n48729, 
      n48730, n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738, 
      n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747, 
      n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755, n48756, 
      n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764, n48765, 
      n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774, 
      n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782, n48783, 
      n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792, 
      n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801, 
      n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810, 
      n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819, 
      n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828, 
      n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837, 
      n48838, n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846, 
      n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855, 
      n48856, n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864, 
      n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872, n48873, 
      n48874, n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882, 
      n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891, 
      n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900, 
      n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908, n48909, 
      n48910, n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918, 
      n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926, n48927, 
      n48928, n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936, 
      n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944, n48945, 
      n48946, n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954, 
      n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963, 
      n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972, 
      n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980, n48981, 
      n48982, n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990, 
      n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998, n48999, 
      n49000, n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008, 
      n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016, n49017, 
      n49018, n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026, 
      n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035, 
      n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043, n49044, 
      n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052, n49053, 
      n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062, 
      n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49071, 
      n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080, 
      n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088, n49089, 
      n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, 
      n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, 
      n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, 
      n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, 
      n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, 
      n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, 
      n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, 
      n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, 
      n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, 
      n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, 
      n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, 
      n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, 
      n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, 
      n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, 
      n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, 
      n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, 
      n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, 
      n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, 
      n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, 
      n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, 
      n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, 
      n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, 
      n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, 
      n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, 
      n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, 
      n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, 
      n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, 
      n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, 
      n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, 
      n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, 
      n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, 
      n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, 
      n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, 
      n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, 
      n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, 
      n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, 
      n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, 
      n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, 
      n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, 
      n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, 
      n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, 
      n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, 
      n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, 
      n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, 
      n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, 
      n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, 
      n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, 
      n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, 
      n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, 
      n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, 
      n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, 
      n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, 
      n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, 
      n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, 
      n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, 
      n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, 
      n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, 
      n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, 
      n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, 
      n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, 
      n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, 
      n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, 
      n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, 
      n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, 
      n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, 
      n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, 
      n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, 
      n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, 
      n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, 
      n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, 
      n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, 
      n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, 
      n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, 
      n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, 
      n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, 
      n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, 
      n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, 
      n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, 
      n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, 
      n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, 
      n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, 
      n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, 
      n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, 
      n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, 
      n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, 
      n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, 
      n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, 
      n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, 
      n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, 
      n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, 
      n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, 
      n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, 
      n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, 
      n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, 
      n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, 
      n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, 
      n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, 
      n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, 
      n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, 
      n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, 
      n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, 
      n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, 
      n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, 
      n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, 
      n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, 
      n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, 
      n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, 
      n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, 
      n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, 
      n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, 
      n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, 
      n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, 
      n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, 
      n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, 
      n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, 
      n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, 
      n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, 
      n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, 
      n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, 
      n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, 
      n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, 
      n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, 
      n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, 
      n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, 
      n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, 
      n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, 
      n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, 
      n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, 
      n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, 
      n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, 
      n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, 
      n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, 
      n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, 
      n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, 
      n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, 
      n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, 
      n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, 
      n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, 
      n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, 
      n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, 
      n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, 
      n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, 
      n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, 
      n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, 
      n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, 
      n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, 
      n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, 
      n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, 
      n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, 
      n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, 
      n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, 
      n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, 
      n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, 
      n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, 
      n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, 
      n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, 
      n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, 
      n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, 
      n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, 
      n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, 
      n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, 
      n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, 
      n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, 
      n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, 
      n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, 
      n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, 
      n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, 
      n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, 
      n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, 
      n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, 
      n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, 
      n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, 
      n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, 
      n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, 
      n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, 
      n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, 
      n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, 
      n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, 
      n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, 
      n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, 
      n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, 
      n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, 
      n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, 
      n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, 
      n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, 
      n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, 
      n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, 
      n_3776, n_3777, n_3778, n_3779, n_3780, n_3781 : std_logic;

begin
   
   clk_r_REG13379_S2 : DFFR_X1 port map( D => ENABLE, CK => CLK, RN => 
                           RESET_BAR, Q => n42760, QN => n_1579);
   clk_r_REG13412_S2 : DFFR_X1 port map( D => RD1, CK => CLK, RN => RESET_BAR, 
                           Q => n42758, QN => n_1580);
   clk_r_REG13420_S2 : DFFR_X1 port map( D => RD2, CK => CLK, RN => RESET_BAR, 
                           Q => n42757, QN => n_1581);
   clk_r_REG13499_S7 : DFFR_X1 port map( D => ADD_RD1(4), CK => CLK, RN => 
                           RESET_BAR, Q => n42756, QN => n_1582);
   clk_r_REG13624_S7 : DFFR_X1 port map( D => ADD_RD2(4), CK => CLK, RN => 
                           RESET_BAR, Q => n42755, QN => n_1583);
   clk_r_REG10366_S6 : DFFR_X1 port map( D => DATAIN(31), CK => CLK, RN => 
                           RESET_BAR, Q => n42754, QN => n_1584);
   clk_r_REG10376_S5 : DFFR_X1 port map( D => DATAIN(30), CK => CLK, RN => 
                           n47506, Q => n42753, QN => n_1585);
   clk_r_REG10357_S6 : DFFR_X1 port map( D => DATAIN(29), CK => CLK, RN => 
                           RESET_BAR, Q => n42752, QN => n_1586);
   clk_r_REG10469_S6 : DFFR_X1 port map( D => DATAIN(28), CK => CLK, RN => 
                           RESET_BAR, Q => n42751, QN => n_1587);
   clk_r_REG10462_S6 : DFFR_X1 port map( D => DATAIN(27), CK => CLK, RN => 
                           RESET_BAR, Q => n42750, QN => n_1588);
   clk_r_REG10455_S6 : DFFR_X1 port map( D => DATAIN(26), CK => CLK, RN => 
                           RESET_BAR, Q => n42749, QN => n_1589);
   clk_r_REG10448_S6 : DFFR_X1 port map( D => DATAIN(25), CK => CLK, RN => 
                           RESET_BAR, Q => n42748, QN => n_1590);
   clk_r_REG10439_S12 : DFFR_X1 port map( D => DATAIN(24), CK => CLK, RN => 
                           RESET_BAR, Q => n42747, QN => n_1591);
   clk_r_REG10403_S6 : DFFR_X1 port map( D => DATAIN(23), CK => CLK, RN => 
                           RESET_BAR, Q => n42746, QN => n_1592);
   clk_r_REG10396_S6 : DFFR_X1 port map( D => DATAIN(22), CK => CLK, RN => 
                           RESET_BAR, Q => n42745, QN => n_1593);
   clk_r_REG10389_S5 : DFFR_X1 port map( D => DATAIN(21), CK => CLK, RN => 
                           RESET_BAR, Q => n42744, QN => n_1594);
   clk_r_REG10487_S6 : DFFR_X1 port map( D => DATAIN(20), CK => CLK, RN => 
                           RESET_BAR, Q => n42743, QN => n_1595);
   clk_r_REG10307_S6 : DFFR_X1 port map( D => DATAIN(19), CK => CLK, RN => 
                           RESET_BAR, Q => n42742, QN => n_1596);
   clk_r_REG10480_S5 : DFFR_X1 port map( D => DATAIN(18), CK => CLK, RN => 
                           RESET_BAR, Q => n42741, QN => n_1597);
   clk_r_REG10349_S6 : DFFR_X1 port map( D => DATAIN(17), CK => CLK, RN => 
                           RESET_BAR, Q => n42740, QN => n_1598);
   clk_r_REG10342_S12 : DFFR_X1 port map( D => DATAIN(16), CK => CLK, RN => 
                           RESET_BAR, Q => n42739, QN => n_1599);
   clk_r_REG10618_S12 : DFFR_X1 port map( D => DATAIN(15), CK => CLK, RN => 
                           RESET_BAR, Q => n42738, QN => n_1600);
   clk_r_REG10634_S5 : DFFR_X1 port map( D => DATAIN(14), CK => CLK, RN => 
                           RESET_BAR, Q => n42737, QN => n_1601);
   clk_r_REG10540_S12 : DFFR_X1 port map( D => DATAIN(13), CK => CLK, RN => 
                           RESET_BAR, Q => n42736, QN => n_1602);
   clk_r_REG10521_S5 : DFFR_X1 port map( D => DATAIN(12), CK => CLK, RN => 
                           RESET_BAR, Q => n42735, QN => n_1603);
   clk_r_REG10710_S12 : DFFR_X1 port map( D => DATAIN(11), CK => CLK, RN => 
                           RESET_BAR, Q => n42734, QN => n_1604);
   clk_r_REG10775_S12 : DFFR_X1 port map( D => DATAIN(10), CK => CLK, RN => 
                           RESET_BAR, Q => n42733, QN => n_1605);
   clk_r_REG10838_S12 : DFFR_X1 port map( D => DATAIN(9), CK => CLK, RN => 
                           RESET_BAR, Q => n42732, QN => n_1606);
   clk_r_REG10877_S12 : DFFR_X1 port map( D => DATAIN(8), CK => CLK, RN => 
                           RESET_BAR, Q => n42731, QN => n_1607);
   clk_r_REG10824_S5 : DFFR_X1 port map( D => DATAIN(7), CK => CLK, RN => 
                           RESET_BAR, Q => n42730, QN => n_1608);
   clk_r_REG10415_S5 : DFFR_X1 port map( D => DATAIN(6), CK => CLK, RN => 
                           RESET_BAR, Q => n42729, QN => n_1609);
   clk_r_REG10805_S12 : DFFR_X1 port map( D => DATAIN(5), CK => CLK, RN => 
                           RESET_BAR, Q => n42728, QN => n_1610);
   clk_r_REG10864_S5 : DFFR_X1 port map( D => DATAIN(4), CK => CLK, RN => 
                           RESET_BAR, Q => n42727, QN => n_1611);
   clk_r_REG10791_S5 : DFFR_X1 port map( D => DATAIN(3), CK => CLK, RN => 
                           RESET_BAR, Q => n42726, QN => n_1612);
   clk_r_REG10762_S5 : DFFR_X1 port map( D => DATAIN(2), CK => CLK, RN => 
                           RESET_BAR, Q => n42725, QN => n_1613);
   clk_r_REG10694_S5 : DFFR_X1 port map( D => DATAIN(1), CK => CLK, RN => 
                           RESET_BAR, Q => n42724, QN => n_1614);
   clk_r_REG10321_S8 : DFFR_X1 port map( D => DATAIN(0), CK => CLK, RN => 
                           RESET_BAR, Q => n42723, QN => n_1615);
   clk_r_REG13518_S7 : DFFR_X1 port map( D => ADD_RD1(3), CK => CLK, RN => 
                           RESET_BAR, Q => n_1616, QN => n42722);
   clk_r_REG13620_S7 : DFFR_X1 port map( D => ADD_RD2(3), CK => CLK, RN => 
                           n47506, Q => n_1617, QN => n42721);
   clk_r_REG12000_S1 : DFF_X1 port map( D => n35769, CK => CLK, Q => n_1618, QN
                           => n42720);
   clk_r_REG11933_S1 : DFF_X1 port map( D => n35770, CK => CLK, Q => n_1619, QN
                           => n42719);
   clk_r_REG12702_S1 : DFF_X1 port map( D => n35771, CK => CLK, Q => n_1620, QN
                           => n42718);
   clk_r_REG11788_S1 : DFF_X1 port map( D => n35772, CK => CLK, Q => n_1621, QN
                           => n42717);
   clk_r_REG11913_S1 : DFF_X1 port map( D => n35773, CK => CLK, Q => n_1622, QN
                           => n42716);
   clk_r_REG11856_S1 : DFF_X1 port map( D => n35774, CK => CLK, Q => n_1623, QN
                           => n42715);
   clk_r_REG11911_S1 : DFF_X1 port map( D => n35775, CK => CLK, Q => n_1624, QN
                           => n42714);
   clk_r_REG11349_S1 : DFF_X1 port map( D => n35776, CK => CLK, Q => n_1625, QN
                           => n42713);
   clk_r_REG11568_S1 : DFF_X1 port map( D => n35777, CK => CLK, Q => n_1626, QN
                           => n42712);
   clk_r_REG11347_S1 : DFF_X1 port map( D => n35778, CK => CLK, Q => n_1627, QN
                           => n42711);
   clk_r_REG11548_S1 : DFF_X1 port map( D => n35779, CK => CLK, Q => n_1628, QN
                           => n42710);
   clk_r_REG11786_S1 : DFF_X1 port map( D => n35780, CK => CLK, Q => n_1629, QN
                           => n42709);
   clk_r_REG11327_S1 : DFF_X1 port map( D => n35781, CK => CLK, Q => n_1630, QN
                           => n42708);
   clk_r_REG11325_S1 : DFF_X1 port map( D => n35782, CK => CLK, Q => n_1631, QN
                           => n42707);
   clk_r_REG12700_S1 : DFF_X1 port map( D => n35783, CK => CLK, Q => n_1632, QN
                           => n42706);
   clk_r_REG11646_S1 : DFF_X1 port map( D => n35784, CK => CLK, Q => n_1633, QN
                           => n42705);
   clk_r_REG13364_S1 : DFF_X1 port map( D => n35785, CK => CLK, Q => n_1634, QN
                           => n42704);
   clk_r_REG12698_S1 : DFF_X1 port map( D => n35786, CK => CLK, Q => n_1635, QN
                           => n42703);
   clk_r_REG11766_S1 : DFF_X1 port map( D => n35787, CK => CLK, Q => n_1636, QN
                           => n42702);
   clk_r_REG11626_S1 : DFF_X1 port map( D => n35788, CK => CLK, Q => n_1637, QN
                           => n42701);
   clk_r_REG13275_S1 : DFF_X1 port map( D => n35789, CK => CLK, Q => n_1638, QN
                           => n42700);
   clk_r_REG11546_S1 : DFF_X1 port map( D => n35790, CK => CLK, Q => n_1639, QN
                           => n42699);
   clk_r_REG11909_S1 : DFF_X1 port map( D => n35791, CK => CLK, Q => n_1640, QN
                           => n42698);
   clk_r_REG11624_S1 : DFF_X1 port map( D => n35792, CK => CLK, Q => n_1641, QN
                           => n42697);
   clk_r_REG11764_S1 : DFF_X1 port map( D => n35793, CK => CLK, Q => n_1642, QN
                           => n42696);
   clk_r_REG12320_S1 : DFF_X1 port map( D => n35794, CK => CLK, Q => n_1643, QN
                           => n42695);
   clk_r_REG13273_S1 : DFF_X1 port map( D => n35795, CK => CLK, Q => n_1644, QN
                           => n42694);
   clk_r_REG11714_S1 : DFF_X1 port map( D => n35796, CK => CLK, Q => n_1645, QN
                           => n42693);
   clk_r_REG11437_S1 : DFF_X1 port map( D => n35797, CK => CLK, Q => n_1646, QN
                           => n42692);
   clk_r_REG11712_S1 : DFF_X1 port map( D => n35798, CK => CLK, Q => n_1647, QN
                           => n42691);
   clk_r_REG12129_S1 : DFF_X1 port map( D => n35799, CK => CLK, Q => n_1648, QN
                           => n42690);
   clk_r_REG10951_S1 : DFF_X1 port map( D => n35800, CK => CLK, Q => n_1649, QN
                           => n42689);
   clk_r_REG11854_S1 : DFF_X1 port map( D => n35801, CK => CLK, Q => n_1650, QN
                           => n42688);
   clk_r_REG11544_S1 : DFF_X1 port map( D => n35802, CK => CLK, Q => n_1651, QN
                           => n42687);
   clk_r_REG12127_S1 : DFF_X1 port map( D => n35803, CK => CLK, Q => n_1652, QN
                           => n42686);
   clk_r_REG11852_S1 : DFF_X1 port map( D => n35804, CK => CLK, Q => n_1653, QN
                           => n42685);
   clk_r_REG12193_S1 : DFF_X1 port map( D => n35805, CK => CLK, Q => n_1654, QN
                           => n42684);
   clk_r_REG12893_S1 : DFF_X1 port map( D => n35806, CK => CLK, Q => n_1655, QN
                           => n42683);
   clk_r_REG13209_S1 : DFF_X1 port map( D => n35807, CK => CLK, Q => n_1656, QN
                           => n42682);
   clk_r_REG11998_S1 : DFF_X1 port map( D => n35808, CK => CLK, Q => n_1657, QN
                           => n42681);
   clk_r_REG12125_S1 : DFF_X1 port map( D => n35809, CK => CLK, Q => n_1658, QN
                           => n42680);
   clk_r_REG12123_S1 : DFF_X1 port map( D => n35810, CK => CLK, Q => n_1659, QN
                           => n42679);
   clk_r_REG13362_S1 : DFF_X1 port map( D => n35811, CK => CLK, Q => n_1660, QN
                           => n42678);
   clk_r_REG12318_S1 : DFF_X1 port map( D => n35812, CK => CLK, Q => n_1661, QN
                           => n42677);
   clk_r_REG13360_S1 : DFF_X1 port map( D => n35813, CK => CLK, Q => n_1662, QN
                           => n42676);
   clk_r_REG12696_S1 : DFF_X1 port map( D => n35814, CK => CLK, Q => n_1663, QN
                           => n42675);
   clk_r_REG11542_S1 : DFF_X1 port map( D => n35815, CK => CLK, Q => n_1664, QN
                           => n42674);
   clk_r_REG13358_S1 : DFF_X1 port map( D => n35816, CK => CLK, Q => n_1665, QN
                           => n42673);
   clk_r_REG11850_S1 : DFF_X1 port map( D => n35817, CK => CLK, Q => n_1666, QN
                           => n42672);
   clk_r_REG11622_S1 : DFF_X1 port map( D => n35818, CK => CLK, Q => n_1667, QN
                           => n42671);
   clk_r_REG13207_S1 : DFF_X1 port map( D => n35819, CK => CLK, Q => n_1668, QN
                           => n42670);
   clk_r_REG12694_S1 : DFF_X1 port map( D => n35820, CK => CLK, Q => n_1669, QN
                           => n42669);
   clk_r_REG13271_S1 : DFF_X1 port map( D => n35821, CK => CLK, Q => n_1670, QN
                           => n42668);
   clk_r_REG10949_S1 : DFF_X1 port map( D => n35822, CK => CLK, Q => n_1671, QN
                           => n42667);
   clk_r_REG12891_S1 : DFF_X1 port map( D => n35823, CK => CLK, Q => n_1672, QN
                           => n42666);
   clk_r_REG13356_S1 : DFF_X1 port map( D => n35824, CK => CLK, Q => n_1673, QN
                           => n42665);
   clk_r_REG12316_S1 : DFF_X1 port map( D => n35825, CK => CLK, Q => n_1674, QN
                           => n42664);
   clk_r_REG13145_S1 : DFF_X1 port map( D => n35826, CK => CLK, Q => n_1675, QN
                           => n42663);
   clk_r_REG10947_S1 : DFF_X1 port map( D => n35827, CK => CLK, Q => n_1676, QN
                           => n42662);
   clk_r_REG11848_S1 : DFF_X1 port map( D => n35828, CK => CLK, Q => n_1677, QN
                           => n42661);
   clk_r_REG11435_S1 : DFF_X1 port map( D => n35829, CK => CLK, Q => n_1678, QN
                           => n42660);
   clk_r_REG13143_S1 : DFF_X1 port map( D => n35830, CK => CLK, Q => n_1679, QN
                           => n42659);
   clk_r_REG10945_S1 : DFF_X1 port map( D => n35831, CK => CLK, Q => n_1680, QN
                           => n42658);
   clk_r_REG13205_S1 : DFF_X1 port map( D => n35832, CK => CLK, Q => n_1681, QN
                           => n42657);
   clk_r_REG11996_S1 : DFF_X1 port map( D => n35833, CK => CLK, Q => n_1682, QN
                           => n42656);
   clk_r_REG12121_S1 : DFF_X1 port map( D => n35834, CK => CLK, Q => n_1683, QN
                           => n42655);
   clk_r_REG12191_S1 : DFF_X1 port map( D => n35835, CK => CLK, Q => n_1684, QN
                           => n42654);
   clk_r_REG12314_S1 : DFF_X1 port map( D => n35836, CK => CLK, Q => n_1685, QN
                           => n42653);
   clk_r_REG12065_S1 : DFF_X1 port map( D => n35837, CK => CLK, Q => n_1686, QN
                           => n42652);
   clk_r_REG13354_S1 : DFF_X1 port map( D => n35838, CK => CLK, Q => n_1687, QN
                           => n42651);
   clk_r_REG11907_S1 : DFF_X1 port map( D => n35839, CK => CLK, Q => n_1688, QN
                           => n42650);
   clk_r_REG12189_S1 : DFF_X1 port map( D => n35840, CK => CLK, Q => n_1689, QN
                           => n42649);
   clk_r_REG11644_S1 : DFF_X1 port map( D => n35841, CK => CLK, Q => n_1690, QN
                           => n42648);
   clk_r_REG12889_S1 : DFF_X1 port map( D => n35842, CK => CLK, Q => n_1691, QN
                           => n42647);
   clk_r_REG11846_S1 : DFF_X1 port map( D => n35843, CK => CLK, Q => n_1692, QN
                           => n42646);
   clk_r_REG11976_S1 : DFF_X1 port map( D => n35844, CK => CLK, Q => n_1693, QN
                           => n42645);
   clk_r_REG12119_S1 : DFF_X1 port map( D => n35845, CK => CLK, Q => n_1694, QN
                           => n42644);
   clk_r_REG11762_S1 : DFF_X1 port map( D => n35846, CK => CLK, Q => n_1695, QN
                           => n42643);
   clk_r_REG13187_S1 : DFF_X1 port map( D => n35847, CK => CLK, Q => n_1696, QN
                           => n42642);
   clk_r_REG11323_S1 : DFF_X1 port map( D => n35848, CK => CLK, Q => n_1697, QN
                           => n42641);
   clk_r_REG10923_S1 : DFF_X1 port map( D => n35849, CK => CLK, Q => n_1698, QN
                           => n42640);
   clk_r_REG12063_S1 : DFF_X1 port map( D => n35850, CK => CLK, Q => n_1699, QN
                           => n42639);
   clk_r_REG10921_S1 : DFF_X1 port map( D => n35851, CK => CLK, Q => n_1700, QN
                           => n42638);
   clk_r_REG11433_S1 : DFF_X1 port map( D => n35852, CK => CLK, Q => n_1701, QN
                           => n42637);
   clk_r_REG11824_S1 : DFF_X1 port map( D => n35853, CK => CLK, Q => n_1702, QN
                           => n42636);
   clk_r_REG12169_S1 : DFF_X1 port map( D => n35854, CK => CLK, Q => n_1703, QN
                           => n42635);
   clk_r_REG12103_S1 : DFF_X1 port map( D => n35855, CK => CLK, Q => n_1704, QN
                           => n42634);
   clk_r_REG11974_S1 : DFF_X1 port map( D => n35856, CK => CLK, Q => n_1705, QN
                           => n42633);
   clk_r_REG13141_S1 : DFF_X1 port map( D => n35857, CK => CLK, Q => n_1706, QN
                           => n42632);
   clk_r_REG12061_S1 : DFF_X1 port map( D => n35858, CK => CLK, Q => n_1707, QN
                           => n42631);
   clk_r_REG13185_S1 : DFF_X1 port map( D => n35859, CK => CLK, Q => n_1708, QN
                           => n42630);
   clk_r_REG13139_S1 : DFF_X1 port map( D => n35860, CK => CLK, Q => n_1709, QN
                           => n42629);
   clk_r_REG12294_S1 : DFF_X1 port map( D => n35861, CK => CLK, Q => n_1710, QN
                           => n42628);
   clk_r_REG13336_S1 : DFF_X1 port map( D => n35862, CK => CLK, Q => n_1711, QN
                           => n42627);
   clk_r_REG12059_S1 : DFF_X1 port map( D => n35863, CK => CLK, Q => n_1712, QN
                           => n42626);
   clk_r_REG13137_S1 : DFF_X1 port map( D => n35864, CK => CLK, Q => n_1713, QN
                           => n42625);
   clk_r_REG11972_S1 : DFF_X1 port map( D => n35865, CK => CLK, Q => n_1714, QN
                           => n42624);
   clk_r_REG12101_S1 : DFF_X1 port map( D => n35866, CK => CLK, Q => n_1715, QN
                           => n42623);
   clk_r_REG11822_S1 : DFF_X1 port map( D => n35867, CK => CLK, Q => n_1716, QN
                           => n42622);
   clk_r_REG12292_S1 : DFF_X1 port map( D => n35868, CK => CLK, Q => n_1717, QN
                           => n42621);
   clk_r_REG11431_S1 : DFF_X1 port map( D => n35869, CK => CLK, Q => n_1718, QN
                           => n42620);
   clk_r_REG12869_S1 : DFF_X1 port map( D => n35870, CK => CLK, Q => n_1719, QN
                           => n42619);
   clk_r_REG13269_S1 : DFF_X1 port map( D => n35871, CK => CLK, Q => n_1720, QN
                           => n42618);
   clk_r_REG12057_S1 : DFF_X1 port map( D => n35872, CK => CLK, Q => n_1721, QN
                           => n42617);
   clk_r_REG11994_S1 : DFF_X1 port map( D => n35873, CK => CLK, Q => n_1722, QN
                           => n42616);
   clk_r_REG12117_S1 : DFF_X1 port map( D => n35874, CK => CLK, Q => n_1723, QN
                           => n42615);
   clk_r_REG12187_S1 : DFF_X1 port map( D => n35875, CK => CLK, Q => n_1724, QN
                           => n42614);
   clk_r_REG10943_S1 : DFF_X1 port map( D => n35876, CK => CLK, Q => n_1725, QN
                           => n42613);
   clk_r_REG11429_S1 : DFF_X1 port map( D => n35877, CK => CLK, Q => n_1726, QN
                           => n42612);
   clk_r_REG11844_S1 : DFF_X1 port map( D => n35878, CK => CLK, Q => n_1727, QN
                           => n42611);
   clk_r_REG11427_S1 : DFF_X1 port map( D => n35879, CK => CLK, Q => n_1728, QN
                           => n42610);
   clk_r_REG10941_S1 : DFF_X1 port map( D => n35880, CK => CLK, Q => n_1729, QN
                           => n42609);
   clk_r_REG11842_S1 : DFF_X1 port map( D => n35881, CK => CLK, Q => n_1730, QN
                           => n42608);
   clk_r_REG12185_S1 : DFF_X1 port map( D => n35882, CK => CLK, Q => n_1731, QN
                           => n42607);
   clk_r_REG12115_S1 : DFF_X1 port map( D => n35883, CK => CLK, Q => n_1732, QN
                           => n42606);
   clk_r_REG11992_S1 : DFF_X1 port map( D => n35884, CK => CLK, Q => n_1733, QN
                           => n42605);
   clk_r_REG12312_S1 : DFF_X1 port map( D => n35885, CK => CLK, Q => n_1734, QN
                           => n42604);
   clk_r_REG13352_S1 : DFF_X1 port map( D => n35886, CK => CLK, Q => n_1735, QN
                           => n42603);
   clk_r_REG12256_S1 : DFF_X1 port map( D => n35887, CK => CLK, Q => n_1736, QN
                           => n42602);
   clk_r_REG12829_S1 : DFF_X1 port map( D => n35888, CK => CLK, Q => n_1737, QN
                           => n42601);
   clk_r_REG12765_S1 : DFF_X1 port map( D => n35889, CK => CLK, Q => n_1738, QN
                           => n42600);
   clk_r_REG12867_S1 : DFF_X1 port map( D => n35890, CK => CLK, Q => n_1739, QN
                           => n42599);
   clk_r_REG12763_S1 : DFF_X1 port map( D => n35891, CK => CLK, Q => n_1740, QN
                           => n42598);
   clk_r_REG12827_S1 : DFF_X1 port map( D => n35892, CK => CLK, Q => n_1741, QN
                           => n42597);
   clk_r_REG12254_S1 : DFF_X1 port map( D => n35893, CK => CLK, Q => n_1742, QN
                           => n42596);
   clk_r_REG13350_S1 : DFF_X1 port map( D => n35894, CK => CLK, Q => n_1743, QN
                           => n42595);
   clk_r_REG12887_S1 : DFF_X1 port map( D => n35895, CK => CLK, Q => n_1744, QN
                           => n42594);
   clk_r_REG12885_S1 : DFF_X1 port map( D => n35896, CK => CLK, Q => n_1745, QN
                           => n42593);
   clk_r_REG12883_S1 : DFF_X1 port map( D => n35897, CK => CLK, Q => n_1746, QN
                           => n42592);
   clk_r_REG12881_S1 : DFF_X1 port map( D => n35898, CK => CLK, Q => n_1747, QN
                           => n42591);
   clk_r_REG12310_S1 : DFF_X1 port map( D => n35899, CK => CLK, Q => n_1748, QN
                           => n42590);
   clk_r_REG12055_S1 : DFF_X1 port map( D => n35900, CK => CLK, Q => n_1749, QN
                           => n42589);
   clk_r_REG11990_S1 : DFF_X1 port map( D => n35901, CK => CLK, Q => n_1750, QN
                           => n42588);
   clk_r_REG12099_S1 : DFF_X1 port map( D => n35902, CK => CLK, Q => n_1751, QN
                           => n42587);
   clk_r_REG12183_S1 : DFF_X1 port map( D => n35903, CK => CLK, Q => n_1752, QN
                           => n42586);
   clk_r_REG11840_S1 : DFF_X1 port map( D => n35904, CK => CLK, Q => n_1753, QN
                           => n42585);
   clk_r_REG13135_S1 : DFF_X1 port map( D => n35905, CK => CLK, Q => n_1754, QN
                           => n42584);
   clk_r_REG11321_S1 : DFF_X1 port map( D => n35906, CK => CLK, Q => n_1755, QN
                           => n42583);
   clk_r_REG11505_S1 : DFF_X1 port map( D => n35907, CK => CLK, Q => n_1756, QN
                           => n42582);
   clk_r_REG11620_S1 : DFF_X1 port map( D => n35908, CK => CLK, Q => n_1757, QN
                           => n42581);
   clk_r_REG11503_S1 : DFF_X1 port map( D => n35909, CK => CLK, Q => n_1758, QN
                           => n42580);
   clk_r_REG11540_S1 : DFF_X1 port map( D => n35910, CK => CLK, Q => n_1759, QN
                           => n42579);
   clk_r_REG11501_S1 : DFF_X1 port map( D => n35911, CK => CLK, Q => n_1760, QN
                           => n42578);
   clk_r_REG11905_S1 : DFF_X1 port map( D => n35912, CK => CLK, Q => n_1761, QN
                           => n42577);
   clk_r_REG12053_S1 : DFF_X1 port map( D => n35913, CK => CLK, Q => n_1762, QN
                           => n42576);
   clk_r_REG11618_S1 : DFF_X1 port map( D => n35914, CK => CLK, Q => n_1763, QN
                           => n42575);
   clk_r_REG12051_S1 : DFF_X1 port map( D => n35915, CK => CLK, Q => n_1764, QN
                           => n42574);
   clk_r_REG13133_S1 : DFF_X1 port map( D => n35916, CK => CLK, Q => n_1765, QN
                           => n42573);
   clk_r_REG11319_S1 : DFF_X1 port map( D => n35917, CK => CLK, Q => n_1766, QN
                           => n42572);
   clk_r_REG11903_S1 : DFF_X1 port map( D => n35918, CK => CLK, Q => n_1767, QN
                           => n42571);
   clk_r_REG11317_S1 : DFF_X1 port map( D => n35919, CK => CLK, Q => n_1768, QN
                           => n42570);
   clk_r_REG12692_S1 : DFF_X1 port map( D => n35920, CK => CLK, Q => n_1769, QN
                           => n42569);
   clk_r_REG12690_S1 : DFF_X1 port map( D => n35921, CK => CLK, Q => n_1770, QN
                           => n42568);
   clk_r_REG11901_S1 : DFF_X1 port map( D => n35922, CK => CLK, Q => n_1771, QN
                           => n42567);
   clk_r_REG11538_S1 : DFF_X1 port map( D => n35923, CK => CLK, Q => n_1772, QN
                           => n42566);
   clk_r_REG12688_S1 : DFF_X1 port map( D => n35924, CK => CLK, Q => n_1773, QN
                           => n42565);
   clk_r_REG11616_S1 : DFF_X1 port map( D => n35925, CK => CLK, Q => n_1774, QN
                           => n42564);
   clk_r_REG11536_S1 : DFF_X1 port map( D => n35926, CK => CLK, Q => n_1775, QN
                           => n42563);
   clk_r_REG13267_S1 : DFF_X1 port map( D => n35927, CK => CLK, Q => n_1776, QN
                           => n42562);
   clk_r_REG11760_S1 : DFF_X1 port map( D => n35928, CK => CLK, Q => n_1777, QN
                           => n42561);
   clk_r_REG13265_S1 : DFF_X1 port map( D => n35929, CK => CLK, Q => n_1778, QN
                           => n42560);
   clk_r_REG13263_S1 : DFF_X1 port map( D => n35930, CK => CLK, Q => n_1779, QN
                           => n42559);
   clk_r_REG13113_S1 : DFF_X1 port map( D => n35931, CK => CLK, Q => n_1780, QN
                           => n42558);
   clk_r_REG13111_S1 : DFF_X1 port map( D => n35932, CK => CLK, Q => n_1781, QN
                           => n42557);
   clk_r_REG11425_S1 : DFF_X1 port map( D => n35933, CK => CLK, Q => n_1782, QN
                           => n42556);
   clk_r_REG10919_S1 : DFF_X1 port map( D => n35934, CK => CLK, Q => n_1783, QN
                           => n42555);
   clk_r_REG13109_S1 : DFF_X1 port map( D => n35935, CK => CLK, Q => n_1784, QN
                           => n42554);
   clk_r_REG11614_S1 : DFF_X1 port map( D => n35936, CK => CLK, Q => n_1785, QN
                           => n42553);
   clk_r_REG11499_S1 : DFF_X1 port map( D => n35937, CK => CLK, Q => n_1786, QN
                           => n42552);
   clk_r_REG11758_S1 : DFF_X1 port map( D => n35938, CK => CLK, Q => n_1787, QN
                           => n42551);
   clk_r_REG12035_S1 : DFF_X1 port map( D => n35939, CK => CLK, Q => n_1788, QN
                           => n42550);
   clk_r_REG11534_S1 : DFF_X1 port map( D => n35940, CK => CLK, Q => n_1789, QN
                           => n42549);
   clk_r_REG12686_S1 : DFF_X1 port map( D => n35941, CK => CLK, Q => n_1790, QN
                           => n42548);
   clk_r_REG12252_S1 : DFF_X1 port map( D => n35942, CK => CLK, Q => n_1791, QN
                           => n42547);
   clk_r_REG13107_S1 : DFF_X1 port map( D => n35943, CK => CLK, Q => n_1792, QN
                           => n42546);
   clk_r_REG11315_S1 : DFF_X1 port map( D => n35944, CK => CLK, Q => n_1793, QN
                           => n42545);
   clk_r_REG11899_S1 : DFF_X1 port map( D => n35945, CK => CLK, Q => n_1794, QN
                           => n42544);
   clk_r_REG11756_S1 : DFF_X1 port map( D => n35946, CK => CLK, Q => n_1795, QN
                           => n42543);
   clk_r_REG13131_S1 : DFF_X1 port map( D => n35947, CK => CLK, Q => n_1796, QN
                           => n42542);
   clk_r_REG11497_S1 : DFF_X1 port map( D => n35948, CK => CLK, Q => n_1797, QN
                           => n42541);
   clk_r_REG11532_S1 : DFF_X1 port map( D => n35949, CK => CLK, Q => n_1798, QN
                           => n42540);
   clk_r_REG12250_S1 : DFF_X1 port map( D => n35950, CK => CLK, Q => n_1799, QN
                           => n42539);
   clk_r_REG11612_S1 : DFF_X1 port map( D => n35951, CK => CLK, Q => n_1800, QN
                           => n42538);
   clk_r_REG12684_S1 : DFF_X1 port map( D => n35952, CK => CLK, Q => n_1801, QN
                           => n42537);
   clk_r_REG11897_S1 : DFF_X1 port map( D => n35953, CK => CLK, Q => n_1802, QN
                           => n42536);
   clk_r_REG11313_S1 : DFF_X1 port map( D => n35954, CK => CLK, Q => n_1803, QN
                           => n42535);
   clk_r_REG12049_S1 : DFF_X1 port map( D => n35955, CK => CLK, Q => n_1804, QN
                           => n42534);
   clk_r_REG13129_S1 : DFF_X1 port map( D => n35956, CK => CLK, Q => n_1805, QN
                           => n42533);
   clk_r_REG11754_S1 : DFF_X1 port map( D => n35957, CK => CLK, Q => n_1806, QN
                           => n42532);
   clk_r_REG11752_S1 : DFF_X1 port map( D => n35958, CK => CLK, Q => n_1807, QN
                           => n42531);
   clk_r_REG13183_S1 : DFF_X1 port map( D => n35959, CK => CLK, Q => n_1808, QN
                           => n42530);
   clk_r_REG12290_S1 : DFF_X1 port map( D => n35960, CK => CLK, Q => n_1809, QN
                           => n42529);
   clk_r_REG13181_S1 : DFF_X1 port map( D => n35961, CK => CLK, Q => n_1810, QN
                           => n42528);
   clk_r_REG10917_S1 : DFF_X1 port map( D => n35962, CK => CLK, Q => n_1811, QN
                           => n42527);
   clk_r_REG11409_S1 : DFF_X1 port map( D => n35963, CK => CLK, Q => n_1812, QN
                           => n42526);
   clk_r_REG11970_S1 : DFF_X1 port map( D => n35964, CK => CLK, Q => n_1813, QN
                           => n42525);
   clk_r_REG10915_S1 : DFF_X1 port map( D => n35965, CK => CLK, Q => n_1814, QN
                           => n42524);
   clk_r_REG11968_S1 : DFF_X1 port map( D => n35966, CK => CLK, Q => n_1815, QN
                           => n42523);
   clk_r_REG12167_S1 : DFF_X1 port map( D => n35967, CK => CLK, Q => n_1816, QN
                           => n42522);
   clk_r_REG12165_S1 : DFF_X1 port map( D => n35968, CK => CLK, Q => n_1817, QN
                           => n42521);
   clk_r_REG11495_S1 : DFF_X1 port map( D => n35969, CK => CLK, Q => n_1818, QN
                           => n42520);
   clk_r_REG11493_S1 : DFF_X1 port map( D => n35970, CK => CLK, Q => n_1819, QN
                           => n42519);
   clk_r_REG13203_S1 : DFF_X1 port map( D => n35971, CK => CLK, Q => n_1820, QN
                           => n42518);
   clk_r_REG11491_S1 : DFF_X1 port map( D => n35972, CK => CLK, Q => n_1821, QN
                           => n42517);
   clk_r_REG11489_S1 : DFF_X1 port map( D => n35973, CK => CLK, Q => n_1822, QN
                           => n42516);
   clk_r_REG12761_S1 : DFF_X1 port map( D => n35974, CK => CLK, Q => n_1823, QN
                           => n42515);
   clk_r_REG12825_S1 : DFF_X1 port map( D => n35975, CK => CLK, Q => n_1824, QN
                           => n42514);
   clk_r_REG12759_S1 : DFF_X1 port map( D => n35976, CK => CLK, Q => n_1825, QN
                           => n42513);
   clk_r_REG12823_S1 : DFF_X1 port map( D => n35977, CK => CLK, Q => n_1826, QN
                           => n42512);
   clk_r_REG12757_S1 : DFF_X1 port map( D => n35978, CK => CLK, Q => n_1827, QN
                           => n42511);
   clk_r_REG12821_S1 : DFF_X1 port map( D => n35979, CK => CLK, Q => n_1828, QN
                           => n42510);
   clk_r_REG12755_S1 : DFF_X1 port map( D => n35980, CK => CLK, Q => n_1829, QN
                           => n42509);
   clk_r_REG12819_S1 : DFF_X1 port map( D => n35981, CK => CLK, Q => n_1830, QN
                           => n42508);
   clk_r_REG12817_S1 : DFF_X1 port map( D => n35982, CK => CLK, Q => n_1831, QN
                           => n42507);
   clk_r_REG12232_S1 : DFF_X1 port map( D => n35983, CK => CLK, Q => n_1832, QN
                           => n42506);
   clk_r_REG12815_S1 : DFF_X1 port map( D => n35984, CK => CLK, Q => n_1833, QN
                           => n42505);
   clk_r_REG12795_S1 : DFF_X1 port map( D => n35985, CK => CLK, Q => n_1834, QN
                           => n42504);
   clk_r_REG13179_S1 : DFF_X1 port map( D => n35986, CK => CLK, Q => n_1835, QN
                           => n42503);
   clk_r_REG13177_S1 : DFF_X1 port map( D => n35987, CK => CLK, Q => n_1836, QN
                           => n42502);
   clk_r_REG12230_S1 : DFF_X1 port map( D => n35988, CK => CLK, Q => n_1837, QN
                           => n42501);
   clk_r_REG13261_S1 : DFF_X1 port map( D => n35989, CK => CLK, Q => n_1838, QN
                           => n42500);
   clk_r_REG13259_S1 : DFF_X1 port map( D => n35990, CK => CLK, Q => n_1839, QN
                           => n42499);
   clk_r_REG13257_S1 : DFF_X1 port map( D => n35991, CK => CLK, Q => n_1840, QN
                           => n42498);
   clk_r_REG12228_S1 : DFF_X1 port map( D => n35992, CK => CLK, Q => n_1841, QN
                           => n42497);
   clk_r_REG11710_S1 : DFF_X1 port map( D => n35993, CK => CLK, Q => n_1842, QN
                           => n42496);
   clk_r_REG11708_S1 : DFF_X1 port map( D => n35994, CK => CLK, Q => n_1843, QN
                           => n42495);
   clk_r_REG12753_S1 : DFF_X1 port map( D => n35995, CK => CLK, Q => n_1844, QN
                           => n42494);
   clk_r_REG11706_S1 : DFF_X1 port map( D => n35996, CK => CLK, Q => n_1845, QN
                           => n42493);
   clk_r_REG12163_S1 : DFF_X1 port map( D => n35997, CK => CLK, Q => n_1846, QN
                           => n42492);
   clk_r_REG13255_S1 : DFF_X1 port map( D => n35998, CK => CLK, Q => n_1847, QN
                           => n42491);
   clk_r_REG11820_S1 : DFF_X1 port map( D => n35999, CK => CLK, Q => n_1848, QN
                           => n42490);
   clk_r_REG11487_S1 : DFF_X1 port map( D => n36000, CK => CLK, Q => n_1849, QN
                           => n42489);
   clk_r_REG12793_S1 : DFF_X1 port map( D => n36001, CK => CLK, Q => n_1850, QN
                           => n42488);
   clk_r_REG13175_S1 : DFF_X1 port map( D => n36002, CK => CLK, Q => n_1851, QN
                           => n42487);
   clk_r_REG12097_S1 : DFF_X1 port map( D => n36003, CK => CLK, Q => n_1852, QN
                           => n42486);
   clk_r_REG12226_S1 : DFF_X1 port map( D => n36004, CK => CLK, Q => n_1853, QN
                           => n42485);
   clk_r_REG12288_S1 : DFF_X1 port map( D => n36005, CK => CLK, Q => n_1854, QN
                           => n42484);
   clk_r_REG10913_S1 : DFF_X1 port map( D => n36006, CK => CLK, Q => n_1855, QN
                           => n42483);
   clk_r_REG12751_S1 : DFF_X1 port map( D => n36007, CK => CLK, Q => n_1856, QN
                           => n42482);
   clk_r_REG11407_S1 : DFF_X1 port map( D => n36008, CK => CLK, Q => n_1857, QN
                           => n42481);
   clk_r_REG11966_S1 : DFF_X1 port map( D => n36009, CK => CLK, Q => n_1858, QN
                           => n42480);
   clk_r_REG11964_S1 : DFF_X1 port map( D => n36010, CK => CLK, Q => n_1859, QN
                           => n42479);
   clk_r_REG12248_S1 : DFF_X1 port map( D => n36011, CK => CLK, Q => n_1860, QN
                           => n42478);
   clk_r_REG11962_S1 : DFF_X1 port map( D => n36012, CK => CLK, Q => n_1861, QN
                           => n42477);
   clk_r_REG12224_S1 : DFF_X1 port map( D => n36013, CK => CLK, Q => n_1862, QN
                           => n42476);
   clk_r_REG12749_S1 : DFF_X1 port map( D => n36014, CK => CLK, Q => n_1863, QN
                           => n42475);
   clk_r_REG12747_S1 : DFF_X1 port map( D => n36015, CK => CLK, Q => n_1864, QN
                           => n42474);
   clk_r_REG12745_S1 : DFF_X1 port map( D => n36016, CK => CLK, Q => n_1865, QN
                           => n42473);
   clk_r_REG12791_S1 : DFF_X1 port map( D => n36017, CK => CLK, Q => n_1866, QN
                           => n42472);
   clk_r_REG12743_S1 : DFF_X1 port map( D => n36018, CK => CLK, Q => n_1867, QN
                           => n42471);
   clk_r_REG12789_S1 : DFF_X1 port map( D => n36019, CK => CLK, Q => n_1868, QN
                           => n42470);
   clk_r_REG12787_S1 : DFF_X1 port map( D => n36020, CK => CLK, Q => n_1869, QN
                           => n42469);
   clk_r_REG12286_S1 : DFF_X1 port map( D => n36021, CK => CLK, Q => n_1870, QN
                           => n42468);
   clk_r_REG10911_S1 : DFF_X1 port map( D => n36022, CK => CLK, Q => n_1871, QN
                           => n42467);
   clk_r_REG13173_S1 : DFF_X1 port map( D => n36023, CK => CLK, Q => n_1872, QN
                           => n42466);
   clk_r_REG10909_S1 : DFF_X1 port map( D => n36024, CK => CLK, Q => n_1873, QN
                           => n42465);
   clk_r_REG11960_S1 : DFF_X1 port map( D => n36025, CK => CLK, Q => n_1874, QN
                           => n42464);
   clk_r_REG10907_S1 : DFF_X1 port map( D => n36026, CK => CLK, Q => n_1875, QN
                           => n42463);
   clk_r_REG12284_S1 : DFF_X1 port map( D => n36027, CK => CLK, Q => n_1876, QN
                           => n42462);
   clk_r_REG12222_S1 : DFF_X1 port map( D => n36028, CK => CLK, Q => n_1877, QN
                           => n42461);
   clk_r_REG12785_S1 : DFF_X1 port map( D => n36029, CK => CLK, Q => n_1878, QN
                           => n42460);
   clk_r_REG11405_S1 : DFF_X1 port map( D => n36030, CK => CLK, Q => n_1879, QN
                           => n42459);
   clk_r_REG12033_S1 : DFF_X1 port map( D => n36031, CK => CLK, Q => n_1880, QN
                           => n42458);
   clk_r_REG12813_S1 : DFF_X1 port map( D => n36032, CK => CLK, Q => n_1881, QN
                           => n42457);
   clk_r_REG11485_S1 : DFF_X1 port map( D => n36033, CK => CLK, Q => n_1882, QN
                           => n42456);
   clk_r_REG12682_S1 : DFF_X1 port map( D => n36034, CK => CLK, Q => n_1883, QN
                           => n42455);
   clk_r_REG12031_S1 : DFF_X1 port map( D => n36035, CK => CLK, Q => n_1884, QN
                           => n42454);
   clk_r_REG13253_S1 : DFF_X1 port map( D => n36036, CK => CLK, Q => n_1885, QN
                           => n42453);
   clk_r_REG11311_S1 : DFF_X1 port map( D => n36037, CK => CLK, Q => n_1886, QN
                           => n42452);
   clk_r_REG11895_S1 : DFF_X1 port map( D => n36038, CK => CLK, Q => n_1887, QN
                           => n42451);
   clk_r_REG11483_S1 : DFF_X1 port map( D => n36039, CK => CLK, Q => n_1888, QN
                           => n42450);
   clk_r_REG11784_S1 : DFF_X1 port map( D => n36040, CK => CLK, Q => n_1889, QN
                           => n42449);
   clk_r_REG11893_S1 : DFF_X1 port map( D => n36041, CK => CLK, Q => n_1890, QN
                           => n42448);
   clk_r_REG11309_S1 : DFF_X1 port map( D => n36042, CK => CLK, Q => n_1891, QN
                           => n42447);
   clk_r_REG11891_S1 : DFF_X1 port map( D => n36043, CK => CLK, Q => n_1892, QN
                           => n42446);
   clk_r_REG11704_S1 : DFF_X1 port map( D => n36044, CK => CLK, Q => n_1893, QN
                           => n42445);
   clk_r_REG12029_S1 : DFF_X1 port map( D => n36045, CK => CLK, Q => n_1894, QN
                           => n42444);
   clk_r_REG11530_S1 : DFF_X1 port map( D => n36046, CK => CLK, Q => n_1895, QN
                           => n42443);
   clk_r_REG11818_S1 : DFF_X1 port map( D => n36047, CK => CLK, Q => n_1896, QN
                           => n42442);
   clk_r_REG11610_S1 : DFF_X1 port map( D => n36048, CK => CLK, Q => n_1897, QN
                           => n42441);
   clk_r_REG11608_S1 : DFF_X1 port map( D => n36049, CK => CLK, Q => n_1898, QN
                           => n42440);
   clk_r_REG11606_S1 : DFF_X1 port map( D => n36050, CK => CLK, Q => n_1899, QN
                           => n42439);
   clk_r_REG11566_S1 : DFF_X1 port map( D => n36051, CK => CLK, Q => n_1900, QN
                           => n42438);
   clk_r_REG12246_S1 : DFF_X1 port map( D => n36052, CK => CLK, Q => n_1901, QN
                           => n42437);
   clk_r_REG11750_S1 : DFF_X1 port map( D => n36053, CK => CLK, Q => n_1902, QN
                           => n42436);
   clk_r_REG11307_S1 : DFF_X1 port map( D => n36054, CK => CLK, Q => n_1903, QN
                           => n42435);
   clk_r_REG13251_S1 : DFF_X1 port map( D => n36055, CK => CLK, Q => n_1904, QN
                           => n42434);
   clk_r_REG11642_S1 : DFF_X1 port map( D => n36056, CK => CLK, Q => n_1905, QN
                           => n42433);
   clk_r_REG11748_S1 : DFF_X1 port map( D => n36057, CK => CLK, Q => n_1906, QN
                           => n42432);
   clk_r_REG11816_S1 : DFF_X1 port map( D => n36058, CK => CLK, Q => n_1907, QN
                           => n42431);
   clk_r_REG13249_S1 : DFF_X1 port map( D => n36059, CK => CLK, Q => n_1908, QN
                           => n42430);
   clk_r_REG11889_S1 : DFF_X1 port map( D => n36060, CK => CLK, Q => n_1909, QN
                           => n42429);
   clk_r_REG11814_S1 : DFF_X1 port map( D => n36061, CK => CLK, Q => n_1910, QN
                           => n42428);
   clk_r_REG11931_S1 : DFF_X1 port map( D => n36062, CK => CLK, Q => n_1911, QN
                           => n42427);
   clk_r_REG11528_S1 : DFF_X1 port map( D => n36063, CK => CLK, Q => n_1912, QN
                           => n42426);
   clk_r_REG12161_S1 : DFF_X1 port map( D => n36064, CK => CLK, Q => n_1913, QN
                           => n42425);
   clk_r_REG11481_S1 : DFF_X1 port map( D => n36065, CK => CLK, Q => n_1914, QN
                           => n42424);
   clk_r_REG12159_S1 : DFF_X1 port map( D => n36066, CK => CLK, Q => n_1915, QN
                           => n42423);
   clk_r_REG11526_S1 : DFF_X1 port map( D => n36067, CK => CLK, Q => n_1916, QN
                           => n42422);
   clk_r_REG12095_S1 : DFF_X1 port map( D => n36068, CK => CLK, Q => n_1917, QN
                           => n42421);
   clk_r_REG12662_S1 : DFF_X1 port map( D => n36069, CK => CLK, Q => n_1918, QN
                           => n42420);
   clk_r_REG11564_S1 : DFF_X1 port map( D => n36070, CK => CLK, Q => n_1919, QN
                           => n42419);
   clk_r_REG12157_S1 : DFF_X1 port map( D => n36071, CK => CLK, Q => n_1920, QN
                           => n42418);
   clk_r_REG12680_S1 : DFF_X1 port map( D => n36072, CK => CLK, Q => n_1921, QN
                           => n42417);
   clk_r_REG11469_S1 : DFF_X1 port map( D => n36073, CK => CLK, Q => n_1922, QN
                           => n42416);
   clk_r_REG11782_S1 : DFF_X1 port map( D => n36074, CK => CLK, Q => n_1923, QN
                           => n42415);
   clk_r_REG11345_S1 : DFF_X1 port map( D => n36075, CK => CLK, Q => n_1924, QN
                           => n42414);
   clk_r_REG12113_S1 : DFF_X1 port map( D => n36076, CK => CLK, Q => n_1925, QN
                           => n42413);
   clk_r_REG11640_S1 : DFF_X1 port map( D => n36077, CK => CLK, Q => n_1926, QN
                           => n42412);
   clk_r_REG12678_S1 : DFF_X1 port map( D => n36078, CK => CLK, Q => n_1927, QN
                           => n42411);
   clk_r_REG11305_S1 : DFF_X1 port map( D => n36079, CK => CLK, Q => n_1928, QN
                           => n42410);
   clk_r_REG12093_S1 : DFF_X1 port map( D => n36080, CK => CLK, Q => n_1929, QN
                           => n42409);
   clk_r_REG11780_S1 : DFF_X1 port map( D => n36081, CK => CLK, Q => n_1930, QN
                           => n42408);
   clk_r_REG12676_S1 : DFF_X1 port map( D => n36082, CK => CLK, Q => n_1931, QN
                           => n42407);
   clk_r_REG13171_S1 : DFF_X1 port map( D => n36083, CK => CLK, Q => n_1932, QN
                           => n42406);
   clk_r_REG13169_S1 : DFF_X1 port map( D => n36084, CK => CLK, Q => n_1933, QN
                           => n42405);
   clk_r_REG13167_S1 : DFF_X1 port map( D => n36085, CK => CLK, Q => n_1934, QN
                           => n42404);
   clk_r_REG13165_S1 : DFF_X1 port map( D => n36086, CK => CLK, Q => n_1935, QN
                           => n42403);
   clk_r_REG13163_S1 : DFF_X1 port map( D => n36087, CK => CLK, Q => n_1936, QN
                           => n42402);
   clk_r_REG11812_S1 : DFF_X1 port map( D => n36088, CK => CLK, Q => n_1937, QN
                           => n42401);
   clk_r_REG13334_S1 : DFF_X1 port map( D => n36089, CK => CLK, Q => n_1938, QN
                           => n42400);
   clk_r_REG11810_S1 : DFF_X1 port map( D => n36090, CK => CLK, Q => n_1939, QN
                           => n42399);
   clk_r_REG11808_S1 : DFF_X1 port map( D => n36091, CK => CLK, Q => n_1940, QN
                           => n42398);
   clk_r_REG11838_S1 : DFF_X1 port map( D => n36092, CK => CLK, Q => n_1941, QN
                           => n42397);
   clk_r_REG11806_S1 : DFF_X1 port map( D => n36093, CK => CLK, Q => n_1942, QN
                           => n42396);
   clk_r_REG11836_S1 : DFF_X1 port map( D => n36094, CK => CLK, Q => n_1943, QN
                           => n42395);
   clk_r_REG13127_S1 : DFF_X1 port map( D => n36095, CK => CLK, Q => n_1944, QN
                           => n42394);
   clk_r_REG12155_S1 : DFF_X1 port map( D => n36096, CK => CLK, Q => n_1945, QN
                           => n42393);
   clk_r_REG12153_S1 : DFF_X1 port map( D => n36097, CK => CLK, Q => n_1946, QN
                           => n42392);
   clk_r_REG12151_S1 : DFF_X1 port map( D => n36098, CK => CLK, Q => n_1947, QN
                           => n42391);
   clk_r_REG12149_S1 : DFF_X1 port map( D => n36099, CK => CLK, Q => n_1948, QN
                           => n42390);
   clk_r_REG12282_S1 : DFF_X1 port map( D => n36100, CK => CLK, Q => n_1949, QN
                           => n42389);
   clk_r_REG12181_S1 : DFF_X1 port map( D => n36101, CK => CLK, Q => n_1950, QN
                           => n42388);
   clk_r_REG12091_S1 : DFF_X1 port map( D => n36102, CK => CLK, Q => n_1951, QN
                           => n42387);
   clk_r_REG12089_S1 : DFF_X1 port map( D => n36103, CK => CLK, Q => n_1952, QN
                           => n42386);
   clk_r_REG12087_S1 : DFF_X1 port map( D => n36104, CK => CLK, Q => n_1953, QN
                           => n42385);
   clk_r_REG12085_S1 : DFF_X1 port map( D => n36105, CK => CLK, Q => n_1954, QN
                           => n42384);
   clk_r_REG12083_S1 : DFF_X1 port map( D => n36106, CK => CLK, Q => n_1955, QN
                           => n42383);
   clk_r_REG11958_S1 : DFF_X1 port map( D => n36107, CK => CLK, Q => n_1956, QN
                           => n42382);
   clk_r_REG11988_S1 : DFF_X1 port map( D => n36108, CK => CLK, Q => n_1957, QN
                           => n42381);
   clk_r_REG12047_S1 : DFF_X1 port map( D => n36109, CK => CLK, Q => n_1958, QN
                           => n42380);
   clk_r_REG11956_S1 : DFF_X1 port map( D => n36110, CK => CLK, Q => n_1959, QN
                           => n42379);
   clk_r_REG11986_S1 : DFF_X1 port map( D => n36111, CK => CLK, Q => n_1960, QN
                           => n42378);
   clk_r_REG10939_S1 : DFF_X1 port map( D => n36112, CK => CLK, Q => n_1961, QN
                           => n42377);
   clk_r_REG10905_S1 : DFF_X1 port map( D => n36113, CK => CLK, Q => n_1962, QN
                           => n42376);
   clk_r_REG10903_S1 : DFF_X1 port map( D => n36114, CK => CLK, Q => n_1963, QN
                           => n42375);
   clk_r_REG10901_S1 : DFF_X1 port map( D => n36115, CK => CLK, Q => n_1964, QN
                           => n42374);
   clk_r_REG10937_S1 : DFF_X1 port map( D => n36116, CK => CLK, Q => n_1965, QN
                           => n42373);
   clk_r_REG10899_S1 : DFF_X1 port map( D => n36117, CK => CLK, Q => n_1966, QN
                           => n42372);
   clk_r_REG11403_S1 : DFF_X1 port map( D => n36118, CK => CLK, Q => n_1967, QN
                           => n42371);
   clk_r_REG11401_S1 : DFF_X1 port map( D => n36119, CK => CLK, Q => n_1968, QN
                           => n42370);
   clk_r_REG11399_S1 : DFF_X1 port map( D => n36120, CK => CLK, Q => n_1969, QN
                           => n42369);
   clk_r_REG11397_S1 : DFF_X1 port map( D => n36121, CK => CLK, Q => n_1970, QN
                           => n42368);
   clk_r_REG11423_S1 : DFF_X1 port map( D => n36122, CK => CLK, Q => n_1971, QN
                           => n42367);
   clk_r_REG11395_S1 : DFF_X1 port map( D => n36123, CK => CLK, Q => n_1972, QN
                           => n42366);
   clk_r_REG10935_S1 : DFF_X1 port map( D => n36124, CK => CLK, Q => n_1973, QN
                           => n42365);
   clk_r_REG11421_S1 : DFF_X1 port map( D => n36125, CK => CLK, Q => n_1974, QN
                           => n42364);
   clk_r_REG11804_S1 : DFF_X1 port map( D => n36126, CK => CLK, Q => n_1975, QN
                           => n42363);
   clk_r_REG12081_S1 : DFF_X1 port map( D => n36127, CK => CLK, Q => n_1976, QN
                           => n42362);
   clk_r_REG12879_S1 : DFF_X1 port map( D => n36128, CK => CLK, Q => n_1977, QN
                           => n42361);
   clk_r_REG13348_S1 : DFF_X1 port map( D => n36129, CK => CLK, Q => n_1978, QN
                           => n42360);
   clk_r_REG12308_S1 : DFF_X1 port map( D => n36130, CK => CLK, Q => n_1979, QN
                           => n42359);
   clk_r_REG13201_S1 : DFF_X1 port map( D => n36131, CK => CLK, Q => n_1980, QN
                           => n42358);
   clk_r_REG13125_S1 : DFF_X1 port map( D => n36132, CK => CLK, Q => n_1981, QN
                           => n42357);
   clk_r_REG13161_S1 : DFF_X1 port map( D => n36133, CK => CLK, Q => n_1982, QN
                           => n42356);
   clk_r_REG12027_S1 : DFF_X1 port map( D => n36134, CK => CLK, Q => n_1983, QN
                           => n42355);
   clk_r_REG11954_S1 : DFF_X1 port map( D => n36135, CK => CLK, Q => n_1984, QN
                           => n42354);
   clk_r_REG12079_S1 : DFF_X1 port map( D => n36136, CK => CLK, Q => n_1985, QN
                           => n42353);
   clk_r_REG11802_S1 : DFF_X1 port map( D => n36137, CK => CLK, Q => n_1986, QN
                           => n42352);
   clk_r_REG11393_S1 : DFF_X1 port map( D => n36138, CK => CLK, Q => n_1987, QN
                           => n42351);
   clk_r_REG10897_S1 : DFF_X1 port map( D => n36139, CK => CLK, Q => n_1988, QN
                           => n42350);
   clk_r_REG12865_S1 : DFF_X1 port map( D => n36140, CK => CLK, Q => n_1989, QN
                           => n42349);
   clk_r_REG13332_S1 : DFF_X1 port map( D => n36141, CK => CLK, Q => n_1990, QN
                           => n42348);
   clk_r_REG12280_S1 : DFF_X1 port map( D => n36142, CK => CLK, Q => n_1991, QN
                           => n42347);
   clk_r_REG13105_S1 : DFF_X1 port map( D => n36143, CK => CLK, Q => n_1992, QN
                           => n42346);
   clk_r_REG12025_S1 : DFF_X1 port map( D => n36144, CK => CLK, Q => n_1993, QN
                           => n42345);
   clk_r_REG12741_S1 : DFF_X1 port map( D => n36145, CK => CLK, Q => n_1994, QN
                           => n42344);
   clk_r_REG12783_S1 : DFF_X1 port map( D => n36146, CK => CLK, Q => n_1995, QN
                           => n42343);
   clk_r_REG12244_S1 : DFF_X1 port map( D => n36147, CK => CLK, Q => n_1996, QN
                           => n42342);
   clk_r_REG11467_S1 : DFF_X1 port map( D => n36148, CK => CLK, Q => n_1997, QN
                           => n42341);
   clk_r_REG12811_S1 : DFF_X1 port map( D => n36149, CK => CLK, Q => n_1998, QN
                           => n42340);
   clk_r_REG12242_S1 : DFF_X1 port map( D => n36150, CK => CLK, Q => n_1999, QN
                           => n42339);
   clk_r_REG12220_S1 : DFF_X1 port map( D => n36151, CK => CLK, Q => n_2000, QN
                           => n42338);
   clk_r_REG11465_S1 : DFF_X1 port map( D => n36152, CK => CLK, Q => n_2001, QN
                           => n42337);
   clk_r_REG11463_S1 : DFF_X1 port map( D => n36153, CK => CLK, Q => n_2002, QN
                           => n42336);
   clk_r_REG12809_S1 : DFF_X1 port map( D => n36154, CK => CLK, Q => n_2003, QN
                           => n42335);
   clk_r_REG12218_S1 : DFF_X1 port map( D => n36155, CK => CLK, Q => n_2004, QN
                           => n42334);
   clk_r_REG12216_S1 : DFF_X1 port map( D => n36156, CK => CLK, Q => n_2005, QN
                           => n42333);
   clk_r_REG12214_S1 : DFF_X1 port map( D => n36157, CK => CLK, Q => n_2006, QN
                           => n42332);
   clk_r_REG11694_S1 : DFF_X1 port map( D => n36158, CK => CLK, Q => n_2007, QN
                           => n42331);
   clk_r_REG11692_S1 : DFF_X1 port map( D => n36159, CK => CLK, Q => n_2008, QN
                           => n42330);
   clk_r_REG11461_S1 : DFF_X1 port map( D => n36160, CK => CLK, Q => n_2009, QN
                           => n42329);
   clk_r_REG12674_S1 : DFF_X1 port map( D => n36161, CK => CLK, Q => n_2010, QN
                           => n42328);
   clk_r_REG11459_S1 : DFF_X1 port map( D => n36162, CK => CLK, Q => n_2011, QN
                           => n42327);
   clk_r_REG11524_S1 : DFF_X1 port map( D => n36163, CK => CLK, Q => n_2012, QN
                           => n42326);
   clk_r_REG11303_S1 : DFF_X1 port map( D => n36164, CK => CLK, Q => n_2013, QN
                           => n42325);
   clk_r_REG11604_S1 : DFF_X1 port map( D => n36165, CK => CLK, Q => n_2014, QN
                           => n42324);
   clk_r_REG11746_S1 : DFF_X1 port map( D => n36166, CK => CLK, Q => n_2015, QN
                           => n42323);
   clk_r_REG11887_S1 : DFF_X1 port map( D => n36167, CK => CLK, Q => n_2016, QN
                           => n42322);
   clk_r_REG11744_S1 : DFF_X1 port map( D => n36168, CK => CLK, Q => n_2017, QN
                           => n42321);
   clk_r_REG11602_S1 : DFF_X1 port map( D => n36169, CK => CLK, Q => n_2018, QN
                           => n42320);
   clk_r_REG11301_S1 : DFF_X1 port map( D => n36170, CK => CLK, Q => n_2019, QN
                           => n42319);
   clk_r_REG11522_S1 : DFF_X1 port map( D => n36171, CK => CLK, Q => n_2020, QN
                           => n42318);
   clk_r_REG11885_S1 : DFF_X1 port map( D => n36172, CK => CLK, Q => n_2021, QN
                           => n42317);
   clk_r_REG11457_S1 : DFF_X1 port map( D => n36173, CK => CLK, Q => n_2022, QN
                           => n42316);
   clk_r_REG12660_S1 : DFF_X1 port map( D => n36174, CK => CLK, Q => n_2023, QN
                           => n42315);
   clk_r_REG11690_S1 : DFF_X1 port map( D => n36175, CK => CLK, Q => n_2024, QN
                           => n42314);
   clk_r_REG13247_S1 : DFF_X1 port map( D => n36176, CK => CLK, Q => n_2025, QN
                           => n42313);
   clk_r_REG13245_S1 : DFF_X1 port map( D => n36177, CK => CLK, Q => n_2026, QN
                           => n42312);
   clk_r_REG11702_S1 : DFF_X1 port map( D => n36178, CK => CLK, Q => n_2027, QN
                           => n42311);
   clk_r_REG13243_S1 : DFF_X1 port map( D => n36179, CK => CLK, Q => n_2028, QN
                           => n42310);
   clk_r_REG11700_S1 : DFF_X1 port map( D => n36180, CK => CLK, Q => n_2029, QN
                           => n42309);
   clk_r_REG13241_S1 : DFF_X1 port map( D => n36181, CK => CLK, Q => n_2030, QN
                           => n42308);
   clk_r_REG11698_S1 : DFF_X1 port map( D => n36182, CK => CLK, Q => n_2031, QN
                           => n42307);
   clk_r_REG13239_S1 : DFF_X1 port map( D => n36183, CK => CLK, Q => n_2032, QN
                           => n42306);
   clk_r_REG11696_S1 : DFF_X1 port map( D => n36185, CK => CLK, Q => n_2033, QN
                           => n42305);
   clk_r_REG13103_S1 : DFF_X1 port map( D => n36186, CK => CLK, Q => n_2034, QN
                           => n42304);
   clk_r_REG13123_S1 : DFF_X1 port map( D => n36187, CK => CLK, Q => n_2035, QN
                           => n42303);
   clk_r_REG11688_S1 : DFF_X1 port map( D => n36188, CK => CLK, Q => n_2036, QN
                           => n42302);
   clk_r_REG11455_S1 : DFF_X1 port map( D => n36189, CK => CLK, Q => n_2037, QN
                           => n42301);
   clk_r_REG11453_S1 : DFF_X1 port map( D => n36190, CK => CLK, Q => n_2038, QN
                           => n42300);
   clk_r_REG11883_S1 : DFF_X1 port map( D => n36191, CK => CLK, Q => n_2039, QN
                           => n42299);
   clk_r_REG13101_S1 : DFF_X1 port map( D => n36192, CK => CLK, Q => n_2040, QN
                           => n42298);
   clk_r_REG13159_S1 : DFF_X1 port map( D => n36193, CK => CLK, Q => n_2041, QN
                           => n42297);
   clk_r_REG11299_S1 : DFF_X1 port map( D => n36194, CK => CLK, Q => n_2042, QN
                           => n42296);
   clk_r_REG13099_S1 : DFF_X1 port map( D => n36195, CK => CLK, Q => n_2043, QN
                           => n42295);
   clk_r_REG11881_S1 : DFF_X1 port map( D => n36196, CK => CLK, Q => n_2044, QN
                           => n42294);
   clk_r_REG13097_S1 : DFF_X1 port map( D => n36197, CK => CLK, Q => n_2045, QN
                           => n42293);
   clk_r_REG11297_S1 : DFF_X1 port map( D => n36198, CK => CLK, Q => n_2046, QN
                           => n42292);
   clk_r_REG12807_S1 : DFF_X1 port map( D => n36199, CK => CLK, Q => n_2047, QN
                           => n42291);
   clk_r_REG11742_S1 : DFF_X1 port map( D => n36200, CK => CLK, Q => n_2048, QN
                           => n42290);
   clk_r_REG11952_S1 : DFF_X1 port map( D => n36201, CK => CLK, Q => n_2049, QN
                           => n42289);
   clk_r_REG11778_S1 : DFF_X1 port map( D => n36202, CK => CLK, Q => n_2050, QN
                           => n42288);
   clk_r_REG11929_S1 : DFF_X1 port map( D => n36203, CK => CLK, Q => n_2051, QN
                           => n42287);
   clk_r_REG11927_S1 : DFF_X1 port map( D => n36204, CK => CLK, Q => n_2052, QN
                           => n42286);
   clk_r_REG11879_S1 : DFF_X1 port map( D => n36205, CK => CLK, Q => n_2053, QN
                           => n42285);
   clk_r_REG11877_S1 : DFF_X1 port map( D => n36206, CK => CLK, Q => n_2054, QN
                           => n42284);
   clk_r_REG12658_S1 : DFF_X1 port map( D => n36207, CK => CLK, Q => n_2055, QN
                           => n42283);
   clk_r_REG11343_S1 : DFF_X1 port map( D => n36208, CK => CLK, Q => n_2056, QN
                           => n42282);
   clk_r_REG11600_S1 : DFF_X1 port map( D => n36209, CK => CLK, Q => n_2057, QN
                           => n42281);
   clk_r_REG11776_S1 : DFF_X1 port map( D => n36210, CK => CLK, Q => n_2058, QN
                           => n42280);
   clk_r_REG11740_S1 : DFF_X1 port map( D => n36211, CK => CLK, Q => n_2059, QN
                           => n42279);
   clk_r_REG11341_S1 : DFF_X1 port map( D => n36212, CK => CLK, Q => n_2060, QN
                           => n42278);
   clk_r_REG11295_S1 : DFF_X1 port map( D => n36213, CK => CLK, Q => n_2061, QN
                           => n42277);
   clk_r_REG11598_S1 : DFF_X1 port map( D => n36214, CK => CLK, Q => n_2062, QN
                           => n42276);
   clk_r_REG11596_S1 : DFF_X1 port map( D => n36215, CK => CLK, Q => n_2063, QN
                           => n42275);
   clk_r_REG11738_S1 : DFF_X1 port map( D => n36216, CK => CLK, Q => n_2064, QN
                           => n42274);
   clk_r_REG12739_S1 : DFF_X1 port map( D => n36217, CK => CLK, Q => n_2065, QN
                           => n42273);
   clk_r_REG11293_S1 : DFF_X1 port map( D => n36218, CK => CLK, Q => n_2066, QN
                           => n42272);
   clk_r_REG12023_S1 : DFF_X1 port map( D => n36219, CK => CLK, Q => n_2067, QN
                           => n42271);
   clk_r_REG11736_S1 : DFF_X1 port map( D => n36220, CK => CLK, Q => n_2068, QN
                           => n42270);
   clk_r_REG11594_S1 : DFF_X1 port map( D => n36221, CK => CLK, Q => n_2069, QN
                           => n42269);
   clk_r_REG12656_S1 : DFF_X1 port map( D => n36222, CK => CLK, Q => n_2070, QN
                           => n42268);
   clk_r_REG11520_S1 : DFF_X1 port map( D => n36223, CK => CLK, Q => n_2071, QN
                           => n42267);
   clk_r_REG11592_S1 : DFF_X1 port map( D => n36224, CK => CLK, Q => n_2072, QN
                           => n42266);
   clk_r_REG13237_S1 : DFF_X1 port map( D => n36225, CK => CLK, Q => n_2073, QN
                           => n42265);
   clk_r_REG13235_S1 : DFF_X1 port map( D => n36226, CK => CLK, Q => n_2074, QN
                           => n42264);
   clk_r_REG11590_S1 : DFF_X1 port map( D => n36227, CK => CLK, Q => n_2075, QN
                           => n42263);
   clk_r_REG11518_S1 : DFF_X1 port map( D => n36228, CK => CLK, Q => n_2076, QN
                           => n42262);
   clk_r_REG12021_S1 : DFF_X1 port map( D => n36229, CK => CLK, Q => n_2077, QN
                           => n42261);
   clk_r_REG12863_S1 : DFF_X1 port map( D => n36230, CK => CLK, Q => n_2078, QN
                           => n42260);
   clk_r_REG13330_S1 : DFF_X1 port map( D => n36231, CK => CLK, Q => n_2079, QN
                           => n42259);
   clk_r_REG12278_S1 : DFF_X1 port map( D => n36232, CK => CLK, Q => n_2080, QN
                           => n42258);
   clk_r_REG12276_S1 : DFF_X1 port map( D => n36233, CK => CLK, Q => n_2081, QN
                           => n42257);
   clk_r_REG12723_S1 : DFF_X1 port map( D => n36234, CK => CLK, Q => n_2082, QN
                           => n42256);
   clk_r_REG12274_S1 : DFF_X1 port map( D => n36235, CK => CLK, Q => n_2083, QN
                           => n42255);
   clk_r_REG12212_S1 : DFF_X1 port map( D => n36236, CK => CLK, Q => n_2084, QN
                           => n42254);
   clk_r_REG12210_S1 : DFF_X1 port map( D => n36237, CK => CLK, Q => n_2085, QN
                           => n42253);
   clk_r_REG12861_S1 : DFF_X1 port map( D => n36238, CK => CLK, Q => n_2086, QN
                           => n42252);
   clk_r_REG12859_S1 : DFF_X1 port map( D => n36239, CK => CLK, Q => n_2087, QN
                           => n42251);
   clk_r_REG11516_S1 : DFF_X1 port map( D => n36240, CK => CLK, Q => n_2088, QN
                           => n42250);
   clk_r_REG13346_S1 : DFF_X1 port map( D => n36241, CK => CLK, Q => n_2089, QN
                           => n42249);
   clk_r_REG12019_S1 : DFF_X1 port map( D => n36242, CK => CLK, Q => n_2090, QN
                           => n42248);
   clk_r_REG12045_S1 : DFF_X1 port map( D => n36243, CK => CLK, Q => n_2091, QN
                           => n42247);
   clk_r_REG12857_S1 : DFF_X1 port map( D => n36244, CK => CLK, Q => n_2092, QN
                           => n42246);
   clk_r_REG12654_S1 : DFF_X1 port map( D => n36245, CK => CLK, Q => n_2093, QN
                           => n42245);
   clk_r_REG12652_S1 : DFF_X1 port map( D => n36246, CK => CLK, Q => n_2094, QN
                           => n42244);
   clk_r_REG12672_S1 : DFF_X1 port map( D => n36247, CK => CLK, Q => n_2095, QN
                           => n42243);
   clk_r_REG12855_S1 : DFF_X1 port map( D => n36248, CK => CLK, Q => n_2096, QN
                           => n42242);
   clk_r_REG11562_S1 : DFF_X1 port map( D => n36249, CK => CLK, Q => n_2097, QN
                           => n42241);
   clk_r_REG11560_S1 : DFF_X1 port map( D => n36250, CK => CLK, Q => n_2098, QN
                           => n42240);
   clk_r_REG12737_S1 : DFF_X1 port map( D => n36251, CK => CLK, Q => n_2099, QN
                           => n42239);
   clk_r_REG12272_S1 : DFF_X1 port map( D => n36252, CK => CLK, Q => n_2100, QN
                           => n42238);
   clk_r_REG12270_S1 : DFF_X1 port map( D => n36253, CK => CLK, Q => n_2101, QN
                           => n42237);
   clk_r_REG12781_S1 : DFF_X1 port map( D => n36254, CK => CLK, Q => n_2102, QN
                           => n42236);
   clk_r_REG11514_S1 : DFF_X1 port map( D => n36255, CK => CLK, Q => n_2103, QN
                           => n42235);
   clk_r_REG12670_S1 : DFF_X1 port map( D => n36256, CK => CLK, Q => n_2104, QN
                           => n42234);
   clk_r_REG12735_S1 : DFF_X1 port map( D => n36257, CK => CLK, Q => n_2105, QN
                           => n42233);
   clk_r_REG12017_S1 : DFF_X1 port map( D => n36258, CK => CLK, Q => n_2106, QN
                           => n42232);
   clk_r_REG12111_S1 : DFF_X1 port map( D => n36259, CK => CLK, Q => n_2107, QN
                           => n42231);
   clk_r_REG11984_S1 : DFF_X1 port map( D => n36260, CK => CLK, Q => n_2108, QN
                           => n42230);
   clk_r_REG12015_S1 : DFF_X1 port map( D => n36261, CK => CLK, Q => n_2109, QN
                           => n42229);
   clk_r_REG12306_S1 : DFF_X1 port map( D => n36262, CK => CLK, Q => n_2110, QN
                           => n42228);
   clk_r_REG13344_S1 : DFF_X1 port map( D => n36263, CK => CLK, Q => n_2111, QN
                           => n42227);
   clk_r_REG12208_S1 : DFF_X1 port map( D => n36264, CK => CLK, Q => n_2112, QN
                           => n42226);
   clk_r_REG12779_S1 : DFF_X1 port map( D => n36265, CK => CLK, Q => n_2113, QN
                           => n42225);
   clk_r_REG11479_S1 : DFF_X1 port map( D => n36266, CK => CLK, Q => n_2114, QN
                           => n42224);
   clk_r_REG11477_S1 : DFF_X1 port map( D => n36267, CK => CLK, Q => n_2115, QN
                           => n42223);
   clk_r_REG12650_S1 : DFF_X1 port map( D => n36268, CK => CLK, Q => n_2116, QN
                           => n42222);
   clk_r_REG11475_S1 : DFF_X1 port map( D => n36269, CK => CLK, Q => n_2117, QN
                           => n42221);
   clk_r_REG11473_S1 : DFF_X1 port map( D => n36270, CK => CLK, Q => n_2118, QN
                           => n42220);
   clk_r_REG11291_S1 : DFF_X1 port map( D => n36271, CK => CLK, Q => n_2119, QN
                           => n42219);
   clk_r_REG11588_S1 : DFF_X1 port map( D => n36272, CK => CLK, Q => n_2120, QN
                           => n42218);
   clk_r_REG12668_S1 : DFF_X1 port map( D => n36273, CK => CLK, Q => n_2121, QN
                           => n42217);
   clk_r_REG11734_S1 : DFF_X1 port map( D => n36274, CK => CLK, Q => n_2122, QN
                           => n42216);
   clk_r_REG11774_S1 : DFF_X1 port map( D => n36275, CK => CLK, Q => n_2123, QN
                           => n42215);
   clk_r_REG11451_S1 : DFF_X1 port map( D => n36276, CK => CLK, Q => n_2124, QN
                           => n42214);
   clk_r_REG11772_S1 : DFF_X1 port map( D => n36277, CK => CLK, Q => n_2125, QN
                           => n42213);
   clk_r_REG11770_S1 : DFF_X1 port map( D => n36278, CK => CLK, Q => n_2126, QN
                           => n42212);
   clk_r_REG12666_S1 : DFF_X1 port map( D => n36279, CK => CLK, Q => n_2127, QN
                           => n42211);
   clk_r_REG12664_S1 : DFF_X1 port map( D => n36281, CK => CLK, Q => n_2128, QN
                           => n42210);
   clk_r_REG11768_S1 : DFF_X1 port map( D => n36283, CK => CLK, Q => n_2129, QN
                           => n42209);
   clk_r_REG11512_S1 : DFF_X1 port map( D => n36284, CK => CLK, Q => n_2130, QN
                           => n42208);
   clk_r_REG11449_S1 : DFF_X1 port map( D => n36285, CK => CLK, Q => n_2131, QN
                           => n42207);
   clk_r_REG12648_S1 : DFF_X1 port map( D => n36286, CK => CLK, Q => n_2132, QN
                           => n42206);
   clk_r_REG12646_S1 : DFF_X1 port map( D => n36287, CK => CLK, Q => n_2133, QN
                           => n42205);
   clk_r_REG12805_S1 : DFF_X1 port map( D => n36288, CK => CLK, Q => n_2134, QN
                           => n42204);
   clk_r_REG11558_S1 : DFF_X1 port map( D => n36289, CK => CLK, Q => n_2135, QN
                           => n42203);
   clk_r_REG11339_S1 : DFF_X1 port map( D => n36290, CK => CLK, Q => n_2136, QN
                           => n42202);
   clk_r_REG12644_S1 : DFF_X1 port map( D => n36291, CK => CLK, Q => n_2137, QN
                           => n42201);
   clk_r_REG12733_S1 : DFF_X1 port map( D => n36292, CK => CLK, Q => n_2138, QN
                           => n42200);
   clk_r_REG12803_S1 : DFF_X1 port map( D => n36293, CK => CLK, Q => n_2139, QN
                           => n42199);
   clk_r_REG11556_S1 : DFF_X1 port map( D => n36294, CK => CLK, Q => n_2140, QN
                           => n42198);
   clk_r_REG12731_S1 : DFF_X1 port map( D => n36295, CK => CLK, Q => n_2141, QN
                           => n42197);
   clk_r_REG11471_S1 : DFF_X1 port map( D => n36297, CK => CLK, Q => n_2142, QN
                           => n42196);
   clk_r_REG11638_S1 : DFF_X1 port map( D => n36298, CK => CLK, Q => n_2143, QN
                           => n42195);
   clk_r_REG11554_S1 : DFF_X1 port map( D => n36299, CK => CLK, Q => n_2144, QN
                           => n42194);
   clk_r_REG11552_S1 : DFF_X1 port map( D => n36300, CK => CLK, Q => n_2145, QN
                           => n42193);
   clk_r_REG11925_S1 : DFF_X1 port map( D => n36301, CK => CLK, Q => n_2146, QN
                           => n42192);
   clk_r_REG11923_S1 : DFF_X1 port map( D => n36302, CK => CLK, Q => n_2147, QN
                           => n42191);
   clk_r_REG11550_S1 : DFF_X1 port map( D => n36304, CK => CLK, Q => n_2148, QN
                           => n42190);
   clk_r_REG11337_S1 : DFF_X1 port map( D => n36305, CK => CLK, Q => n_2149, QN
                           => n42189);
   clk_r_REG11636_S1 : DFF_X1 port map( D => n36306, CK => CLK, Q => n_2150, QN
                           => n42188);
   clk_r_REG11732_S1 : DFF_X1 port map( D => n36307, CK => CLK, Q => n_2151, QN
                           => n42187);
   clk_r_REG11921_S1 : DFF_X1 port map( D => n36308, CK => CLK, Q => n_2152, QN
                           => n42186);
   clk_r_REG12206_S1 : DFF_X1 port map( D => n36309, CK => CLK, Q => n_2153, QN
                           => n42185);
   clk_r_REG11447_S1 : DFF_X1 port map( D => n36310, CK => CLK, Q => n_2154, QN
                           => n42184);
   clk_r_REG11510_S1 : DFF_X1 port map( D => n36311, CK => CLK, Q => n_2155, QN
                           => n42183);
   clk_r_REG11335_S1 : DFF_X1 port map( D => n36312, CK => CLK, Q => n_2156, QN
                           => n42182);
   clk_r_REG11333_S1 : DFF_X1 port map( D => n36313, CK => CLK, Q => n_2157, QN
                           => n42181);
   clk_r_REG11331_S1 : DFF_X1 port map( D => n36314, CK => CLK, Q => n_2158, QN
                           => n42180);
   clk_r_REG11329_S1 : DFF_X1 port map( D => n36316, CK => CLK, Q => n_2159, QN
                           => n42179);
   clk_r_REG11634_S1 : DFF_X1 port map( D => n36317, CK => CLK, Q => n_2160, QN
                           => n42178);
   clk_r_REG11632_S1 : DFF_X1 port map( D => n36318, CK => CLK, Q => n_2161, QN
                           => n42177);
   clk_r_REG11919_S1 : DFF_X1 port map( D => n36319, CK => CLK, Q => n_2162, QN
                           => n42176);
   clk_r_REG11917_S1 : DFF_X1 port map( D => n36320, CK => CLK, Q => n_2163, QN
                           => n42175);
   clk_r_REG11915_S1 : DFF_X1 port map( D => n36322, CK => CLK, Q => n_2164, QN
                           => n42174);
   clk_r_REG11630_S1 : DFF_X1 port map( D => n36323, CK => CLK, Q => n_2165, QN
                           => n42173);
   clk_r_REG11586_S1 : DFF_X1 port map( D => n36324, CK => CLK, Q => n_2166, QN
                           => n42172);
   clk_r_REG11730_S1 : DFF_X1 port map( D => n36325, CK => CLK, Q => n_2167, QN
                           => n42171);
   clk_r_REG11875_S1 : DFF_X1 port map( D => n36326, CK => CLK, Q => n_2168, QN
                           => n42170);
   clk_r_REG10792_S1 : DFF_X1 port map( D => n36328, CK => CLK, Q => n_2169, QN
                           => n42169);
   clk_r_REG11728_S1 : DFF_X1 port map( D => n36329, CK => CLK, Q => n_2170, QN
                           => n42168);
   clk_r_REG11873_S1 : DFF_X1 port map( D => n36330, CK => CLK, Q => n_2171, QN
                           => n42167);
   clk_r_REG11686_S1 : DFF_X1 port map( D => n36331, CK => CLK, Q => n_2172, QN
                           => n42166);
   clk_r_REG11508_S1 : DFF_X1 port map( D => n36332, CK => CLK, Q => n_2173, QN
                           => n42165);
   clk_r_REG11289_S1 : DFF_X1 port map( D => n36333, CK => CLK, Q => n_2174, QN
                           => n42164);
   clk_r_REG11445_S1 : DFF_X1 port map( D => n36334, CK => CLK, Q => n_2175, QN
                           => n42163);
   clk_r_REG12179_S1 : DFF_X1 port map( D => n36335, CK => CLK, Q => n_2176, QN
                           => n42162);
   clk_r_REG12642_S1 : DFF_X1 port map( D => n36336, CK => CLK, Q => n_2177, QN
                           => n42161);
   clk_r_REG13233_S1 : DFF_X1 port map( D => n36337, CK => CLK, Q => n_2178, QN
                           => n42160);
   clk_r_REG11950_S1 : DFF_X1 port map( D => n36338, CK => CLK, Q => n_2179, QN
                           => n42159);
   clk_r_REG12077_S1 : DFF_X1 port map( D => n36339, CK => CLK, Q => n_2180, QN
                           => n42158);
   clk_r_REG13199_S1 : DFF_X1 port map( D => n36340, CK => CLK, Q => n_2181, QN
                           => n42157);
   clk_r_REG12043_S1 : DFF_X1 port map( D => n36341, CK => CLK, Q => n_2182, QN
                           => n42156);
   clk_r_REG12268_S1 : DFF_X1 port map( D => n36342, CK => CLK, Q => n_2183, QN
                           => n42155);
   clk_r_REG13328_S1 : DFF_X1 port map( D => n36343, CK => CLK, Q => n_2184, QN
                           => n42154);
   clk_r_REG12204_S1 : DFF_X1 port map( D => n36344, CK => CLK, Q => n_2185, QN
                           => n42153);
   clk_r_REG12853_S1 : DFF_X1 port map( D => n36345, CK => CLK, Q => n_2186, QN
                           => n42152);
   clk_r_REG12777_S1 : DFF_X1 port map( D => n36346, CK => CLK, Q => n_2187, QN
                           => n42151);
   clk_r_REG12721_S1 : DFF_X1 port map( D => n36347, CK => CLK, Q => n_2188, QN
                           => n42150);
   clk_r_REG13197_S1 : DFF_X1 port map( D => n36348, CK => CLK, Q => n_2189, QN
                           => n42149);
   clk_r_REG13195_S1 : DFF_X1 port map( D => n36349, CK => CLK, Q => n_2190, QN
                           => n42148);
   clk_r_REG13121_S1 : DFF_X1 port map( D => n36350, CK => CLK, Q => n_2191, QN
                           => n42147);
   clk_r_REG13193_S1 : DFF_X1 port map( D => n36351, CK => CLK, Q => n_2192, QN
                           => n42146);
   clk_r_REG13157_S1 : DFF_X1 port map( D => n36352, CK => CLK, Q => n_2193, QN
                           => n42145);
   clk_r_REG13155_S1 : DFF_X1 port map( D => n36353, CK => CLK, Q => n_2194, QN
                           => n42144);
   clk_r_REG13153_S1 : DFF_X1 port map( D => n36354, CK => CLK, Q => n_2195, QN
                           => n42143);
   clk_r_REG13191_S1 : DFF_X1 port map( D => n36355, CK => CLK, Q => n_2196, QN
                           => n42142);
   clk_r_REG13119_S1 : DFF_X1 port map( D => n36356, CK => CLK, Q => n_2197, QN
                           => n42141);
   clk_r_REG13095_S1 : DFF_X1 port map( D => n36357, CK => CLK, Q => n_2198, QN
                           => n42140);
   clk_r_REG13093_S1 : DFF_X1 port map( D => n36358, CK => CLK, Q => n_2199, QN
                           => n42139);
   clk_r_REG13091_S1 : DFF_X1 port map( D => n36359, CK => CLK, Q => n_2200, QN
                           => n42138);
   clk_r_REG13089_S1 : DFF_X1 port map( D => n36360, CK => CLK, Q => n_2201, QN
                           => n42137);
   clk_r_REG13087_S1 : DFF_X1 port map( D => n36361, CK => CLK, Q => n_2202, QN
                           => n42136);
   clk_r_REG13085_S1 : DFF_X1 port map( D => n36362, CK => CLK, Q => n_2203, QN
                           => n42135);
   clk_r_REG11834_S1 : DFF_X1 port map( D => n36363, CK => CLK, Q => n_2204, QN
                           => n42134);
   clk_r_REG12240_S1 : DFF_X1 port map( D => n36364, CK => CLK, Q => n_2205, QN
                           => n42133);
   clk_r_REG12877_S1 : DFF_X1 port map( D => n36365, CK => CLK, Q => n_2206, QN
                           => n42132);
   clk_r_REG12875_S1 : DFF_X1 port map( D => n36366, CK => CLK, Q => n_2207, QN
                           => n42131);
   clk_r_REG12873_S1 : DFF_X1 port map( D => n36367, CK => CLK, Q => n_2208, QN
                           => n42130);
   clk_r_REG12851_S1 : DFF_X1 port map( D => n36368, CK => CLK, Q => n_2209, QN
                           => n42129);
   clk_r_REG12849_S1 : DFF_X1 port map( D => n36369, CK => CLK, Q => n_2210, QN
                           => n42128);
   clk_r_REG12847_S1 : DFF_X1 port map( D => n36370, CK => CLK, Q => n_2211, QN
                           => n42127);
   clk_r_REG12845_S1 : DFF_X1 port map( D => n36371, CK => CLK, Q => n_2212, QN
                           => n42126);
   clk_r_REG11684_S1 : DFF_X1 port map( D => n36372, CK => CLK, Q => n_2213, QN
                           => n42125);
   clk_r_REG11419_S1 : DFF_X1 port map( D => n36373, CK => CLK, Q => n_2214, QN
                           => n42124);
   clk_r_REG10933_S1 : DFF_X1 port map( D => n36374, CK => CLK, Q => n_2215, QN
                           => n42123);
   clk_r_REG11832_S1 : DFF_X1 port map( D => n36375, CK => CLK, Q => n_2216, QN
                           => n42122);
   clk_r_REG12177_S1 : DFF_X1 port map( D => n36376, CK => CLK, Q => n_2217, QN
                           => n42121);
   clk_r_REG12109_S1 : DFF_X1 port map( D => n36377, CK => CLK, Q => n_2218, QN
                           => n42120);
   clk_r_REG11982_S1 : DFF_X1 port map( D => n36378, CK => CLK, Q => n_2219, QN
                           => n42119);
   clk_r_REG12041_S1 : DFF_X1 port map( D => n36379, CK => CLK, Q => n_2220, QN
                           => n42118);
   clk_r_REG12304_S1 : DFF_X1 port map( D => n36380, CK => CLK, Q => n_2221, QN
                           => n42117);
   clk_r_REG13342_S1 : DFF_X1 port map( D => n36381, CK => CLK, Q => n_2222, QN
                           => n42116);
   clk_r_REG10931_S1 : DFF_X1 port map( D => n36382, CK => CLK, Q => n_2223, QN
                           => n42115);
   clk_r_REG11417_S1 : DFF_X1 port map( D => n36383, CK => CLK, Q => n_2224, QN
                           => n42114);
   clk_r_REG11682_S1 : DFF_X1 port map( D => n36384, CK => CLK, Q => n_2225, QN
                           => n42113);
   clk_r_REG11830_S1 : DFF_X1 port map( D => n36385, CK => CLK, Q => n_2226, QN
                           => n42112);
   clk_r_REG12175_S1 : DFF_X1 port map( D => n36386, CK => CLK, Q => n_2227, QN
                           => n42111);
   clk_r_REG12719_S1 : DFF_X1 port map( D => n36387, CK => CLK, Q => n_2228, QN
                           => n42110);
   clk_r_REG10929_S1 : DFF_X1 port map( D => n36388, CK => CLK, Q => n_2229, QN
                           => n42109);
   clk_r_REG11415_S1 : DFF_X1 port map( D => n36389, CK => CLK, Q => n_2230, QN
                           => n42108);
   clk_r_REG11828_S1 : DFF_X1 port map( D => n36390, CK => CLK, Q => n_2231, QN
                           => n42107);
   clk_r_REG11800_S1 : DFF_X1 port map( D => n36391, CK => CLK, Q => n_2232, QN
                           => n42106);
   clk_r_REG11798_S1 : DFF_X1 port map( D => n36392, CK => CLK, Q => n_2233, QN
                           => n42105);
   clk_r_REG11796_S1 : DFF_X1 port map( D => n36393, CK => CLK, Q => n_2234, QN
                           => n42104);
   clk_r_REG12173_S1 : DFF_X1 port map( D => n36394, CK => CLK, Q => n_2235, QN
                           => n42103);
   clk_r_REG12107_S1 : DFF_X1 port map( D => n36395, CK => CLK, Q => n_2236, QN
                           => n42102);
   clk_r_REG11980_S1 : DFF_X1 port map( D => n36396, CK => CLK, Q => n_2237, QN
                           => n42101);
   clk_r_REG12013_S1 : DFF_X1 port map( D => n36397, CK => CLK, Q => n_2238, QN
                           => n42100);
   clk_r_REG10350_S1 : DFF_X1 port map( D => n36399, CK => CLK, Q => n_2239, QN
                           => n42099);
   clk_r_REG12302_S1 : DFF_X1 port map( D => n36400, CK => CLK, Q => n_2240, QN
                           => n42098);
   clk_r_REG13340_S1 : DFF_X1 port map( D => n36401, CK => CLK, Q => n_2241, QN
                           => n42097);
   clk_r_REG12202_S1 : DFF_X1 port map( D => n36402, CK => CLK, Q => n_2242, QN
                           => n42096);
   clk_r_REG10763_S1 : DFF_X1 port map( D => n36404, CK => CLK, Q => n_2243, QN
                           => n42095);
   clk_r_REG11680_S1 : DFF_X1 port map( D => n36405, CK => CLK, Q => n_2244, QN
                           => n42094);
   clk_r_REG12775_S1 : DFF_X1 port map( D => n36406, CK => CLK, Q => n_2245, QN
                           => n42093);
   clk_r_REG12147_S1 : DFF_X1 port map( D => n36407, CK => CLK, Q => n_2246, QN
                           => n42092);
   clk_r_REG12145_S1 : DFF_X1 port map( D => n36408, CK => CLK, Q => n_2247, QN
                           => n42091);
   clk_r_REG12143_S1 : DFF_X1 port map( D => n36409, CK => CLK, Q => n_2248, QN
                           => n42090);
   clk_r_REG12717_S1 : DFF_X1 port map( D => n36410, CK => CLK, Q => n_2249, QN
                           => n42089);
   clk_r_REG12075_S1 : DFF_X1 port map( D => n36411, CK => CLK, Q => n_2250, QN
                           => n42088);
   clk_r_REG11678_S1 : DFF_X1 port map( D => n36412, CK => CLK, Q => n_2251, QN
                           => n42087);
   clk_r_REG12073_S1 : DFF_X1 port map( D => n36413, CK => CLK, Q => n_2252, QN
                           => n42086);
   clk_r_REG11676_S1 : DFF_X1 port map( D => n36414, CK => CLK, Q => n_2253, QN
                           => n42085);
   clk_r_REG11413_S1 : DFF_X1 port map( D => n36415, CK => CLK, Q => n_2254, QN
                           => n42084);
   clk_r_REG12071_S1 : DFF_X1 port map( D => n36416, CK => CLK, Q => n_2255, QN
                           => n42083);
   clk_r_REG10927_S1 : DFF_X1 port map( D => n36417, CK => CLK, Q => n_2256, QN
                           => n42082);
   clk_r_REG11391_S1 : DFF_X1 port map( D => n36418, CK => CLK, Q => n_2257, QN
                           => n42081);
   clk_r_REG11948_S1 : DFF_X1 port map( D => n36419, CK => CLK, Q => n_2258, QN
                           => n42080);
   clk_r_REG10925_S1 : DFF_X1 port map( D => n36421, CK => CLK, Q => n_2259, QN
                           => n42079);
   clk_r_REG11411_S1 : DFF_X1 port map( D => n36423, CK => CLK, Q => n_2260, QN
                           => n42078);
   clk_r_REG11674_S1 : DFF_X1 port map( D => n36424, CK => CLK, Q => n_2261, QN
                           => n42077);
   clk_r_REG10695_S1 : DFF_X1 port map( D => n36426, CK => CLK, Q => n_2262, QN
                           => n42076);
   clk_r_REG11826_S1 : DFF_X1 port map( D => n36428, CK => CLK, Q => n_2263, QN
                           => n42075);
   clk_r_REG12171_S1 : DFF_X1 port map( D => n36430, CK => CLK, Q => n_2264, QN
                           => n42074);
   clk_r_REG12105_S1 : DFF_X1 port map( D => n36432, CK => CLK, Q => n_2265, QN
                           => n42073);
   clk_r_REG11978_S1 : DFF_X1 port map( D => n36434, CK => CLK, Q => n_2266, QN
                           => n42072);
   clk_r_REG12011_S1 : DFF_X1 port map( D => n36435, CK => CLK, Q => n_2267, QN
                           => n42071);
   clk_r_REG12009_S1 : DFF_X1 port map( D => n36436, CK => CLK, Q => n_2268, QN
                           => n42070);
   clk_r_REG12007_S1 : DFF_X1 port map( D => n36437, CK => CLK, Q => n_2269, QN
                           => n42069);
   clk_r_REG12300_S1 : DFF_X1 port map( D => n36438, CK => CLK, Q => n_2270, QN
                           => n42068);
   clk_r_REG12005_S1 : DFF_X1 port map( D => n36439, CK => CLK, Q => n_2271, QN
                           => n42067);
   clk_r_REG11672_S1 : DFF_X1 port map( D => n36440, CK => CLK, Q => n_2272, QN
                           => n42066);
   clk_r_REG10865_S1 : DFF_X1 port map( D => n36442, CK => CLK, Q => n_2273, QN
                           => n42065);
   clk_r_REG11389_S1 : DFF_X1 port map( D => n36443, CK => CLK, Q => n_2274, QN
                           => n42064);
   clk_r_REG11387_S1 : DFF_X1 port map( D => n36444, CK => CLK, Q => n_2275, QN
                           => n42063);
   clk_r_REG11385_S1 : DFF_X1 port map( D => n36445, CK => CLK, Q => n_2276, QN
                           => n42062);
   clk_r_REG10895_S1 : DFF_X1 port map( D => n36446, CK => CLK, Q => n_2277, QN
                           => n42061);
   clk_r_REG10893_S1 : DFF_X1 port map( D => n36447, CK => CLK, Q => n_2278, QN
                           => n42060);
   clk_r_REG11670_S1 : DFF_X1 port map( D => n36448, CK => CLK, Q => n_2279, QN
                           => n42059);
   clk_r_REG10619_S1 : DFF_X1 port map( D => n36450, CK => CLK, Q => n_2280, QN
                           => n42058);
   clk_r_REG10891_S1 : DFF_X1 port map( D => n36451, CK => CLK, Q => n_2281, QN
                           => n42057);
   clk_r_REG12715_S1 : DFF_X1 port map( D => n36452, CK => CLK, Q => n_2282, QN
                           => n42056);
   clk_r_REG12773_S1 : DFF_X1 port map( D => n36453, CK => CLK, Q => n_2283, QN
                           => n42055);
   clk_r_REG10416_S1 : DFF_X1 port map( D => n36455, CK => CLK, Q => n_2284, QN
                           => n42054);
   clk_r_REG11946_S1 : DFF_X1 port map( D => n36456, CK => CLK, Q => n_2285, QN
                           => n42053);
   clk_r_REG10878_S1 : DFF_X1 port map( D => n36458, CK => CLK, Q => n_2286, QN
                           => n42052);
   clk_r_REG13338_S1 : DFF_X1 port map( D => n36459, CK => CLK, Q => n_2287, QN
                           => n42051);
   clk_r_REG12266_S1 : DFF_X1 port map( D => n36460, CK => CLK, Q => n_2288, QN
                           => n42050);
   clk_r_REG12200_S1 : DFF_X1 port map( D => n36461, CK => CLK, Q => n_2289, QN
                           => n42049);
   clk_r_REG12198_S1 : DFF_X1 port map( D => n36462, CK => CLK, Q => n_2290, QN
                           => n42048);
   clk_r_REG12196_S1 : DFF_X1 port map( D => n36463, CK => CLK, Q => n_2291, QN
                           => n42047);
   clk_r_REG13326_S1 : DFF_X1 port map( D => n36464, CK => CLK, Q => n_2292, QN
                           => n42046);
   clk_r_REG12069_S1 : DFF_X1 port map( D => n36465, CK => CLK, Q => n_2293, QN
                           => n42045);
   clk_r_REG13324_S1 : DFF_X1 port map( D => n36466, CK => CLK, Q => n_2294, QN
                           => n42044);
   clk_r_REG11944_S1 : DFF_X1 port map( D => n36467, CK => CLK, Q => n_2295, QN
                           => n42043);
   clk_r_REG12713_S1 : DFF_X1 port map( D => n36468, CK => CLK, Q => n_2296, QN
                           => n42042);
   clk_r_REG10806_S1 : DFF_X1 port map( D => n36470, CK => CLK, Q => n_2297, QN
                           => n42041);
   clk_r_REG12771_S1 : DFF_X1 port map( D => n36471, CK => CLK, Q => n_2298, QN
                           => n42040);
   clk_r_REG10488_S1 : DFF_X1 port map( D => n36473, CK => CLK, Q => n_2299, QN
                           => n42039);
   clk_r_REG12141_S1 : DFF_X1 port map( D => n36474, CK => CLK, Q => n_2300, QN
                           => n42038);
   clk_r_REG12769_S1 : DFF_X1 port map( D => n36475, CK => CLK, Q => n_2301, QN
                           => n42037);
   clk_r_REG11942_S1 : DFF_X1 port map( D => n36476, CK => CLK, Q => n_2302, QN
                           => n42036);
   clk_r_REG12871_S1 : DFF_X1 port map( D => n36478, CK => CLK, Q => n_2303, QN
                           => n42035);
   clk_r_REG12264_S1 : DFF_X1 port map( D => n36479, CK => CLK, Q => n_2304, QN
                           => n42034);
   clk_r_REG13322_S1 : DFF_X1 port map( D => n36480, CK => CLK, Q => n_2305, QN
                           => n42033);
   clk_r_REG12711_S1 : DFF_X1 port map( D => n36481, CK => CLK, Q => n_2306, QN
                           => n42032);
   clk_r_REG12262_S1 : DFF_X1 port map( D => n36482, CK => CLK, Q => n_2307, QN
                           => n42031);
   clk_r_REG12298_S1 : DFF_X1 port map( D => n36483, CK => CLK, Q => n_2308, QN
                           => n42030);
   clk_r_REG13151_S1 : DFF_X1 port map( D => n36484, CK => CLK, Q => n_2309, QN
                           => n42029);
   clk_r_REG10711_S1 : DFF_X1 port map( D => n36486, CK => CLK, Q => n_2310, QN
                           => n42028);
   clk_r_REG10397_S1 : DFF_X1 port map( D => n36488, CK => CLK, Q => n_2311, QN
                           => n42027);
   clk_r_REG11628_S1 : DFF_X1 port map( D => n36490, CK => CLK, Q => n_2312, QN
                           => n42026);
   clk_r_REG12709_S1 : DFF_X1 port map( D => n36491, CK => CLK, Q => n_2313, QN
                           => n42025);
   clk_r_REG13320_S1 : DFF_X1 port map( D => n36492, CK => CLK, Q => n_2314, QN
                           => n42024);
   clk_r_REG13231_S1 : DFF_X1 port map( D => n36494, CK => CLK, Q => n_2315, QN
                           => n42023);
   clk_r_REG13229_S1 : DFF_X1 port map( D => n36495, CK => CLK, Q => n_2316, QN
                           => n42022);
   clk_r_REG13227_S1 : DFF_X1 port map( D => n36496, CK => CLK, Q => n_2317, QN
                           => n42021);
   clk_r_REG13225_S1 : DFF_X1 port map( D => n36497, CK => CLK, Q => n_2318, QN
                           => n42020);
   clk_r_REG13223_S1 : DFF_X1 port map( D => n36498, CK => CLK, Q => n_2319, QN
                           => n42019);
   clk_r_REG13221_S1 : DFF_X1 port map( D => n36499, CK => CLK, Q => n_2320, QN
                           => n42018);
   clk_r_REG13219_S1 : DFF_X1 port map( D => n36500, CK => CLK, Q => n_2321, QN
                           => n42017);
   clk_r_REG13217_S1 : DFF_X1 port map( D => n36501, CK => CLK, Q => n_2322, QN
                           => n42016);
   clk_r_REG13215_S1 : DFF_X1 port map( D => n36502, CK => CLK, Q => n_2323, QN
                           => n42015);
   clk_r_REG10322_S1 : DFF_X1 port map( D => n36504, CK => CLK, Q => n_2324, QN
                           => n42014);
   clk_r_REG12955_S1 : DFF_X1 port map( D => n36506, CK => CLK, Q => n_2325, QN
                           => n42013);
   clk_r_REG12446_S1 : DFF_X1 port map( D => n36507, CK => CLK, Q => n_2326, QN
                           => n42012);
   clk_r_REG12574_S1 : DFF_X1 port map( D => n36509, CK => CLK, Q => n_2327, QN
                           => n42011);
   clk_r_REG12953_S1 : DFF_X1 port map( D => n36510, CK => CLK, Q => n_2328, QN
                           => n42010);
   clk_r_REG12444_S1 : DFF_X1 port map( D => n36512, CK => CLK, Q => n_2329, QN
                           => n42009);
   clk_r_REG12382_S1 : DFF_X1 port map( D => n36513, CK => CLK, Q => n_2330, QN
                           => n42008);
   clk_r_REG10825_S1 : DFF_X1 port map( D => n36516, CK => CLK, Q => n_2331, QN
                           => n42007);
   clk_r_REG12380_S1 : DFF_X1 port map( D => n36517, CK => CLK, Q => n_2332, QN
                           => n42006);
   clk_r_REG12378_S1 : DFF_X1 port map( D => n36518, CK => CLK, Q => n_2333, QN
                           => n42005);
   clk_r_REG12362_S1 : DFF_X1 port map( D => n36520, CK => CLK, Q => n_2334, QN
                           => n42004);
   clk_r_REG12843_S1 : DFF_X1 port map( D => n36521, CK => CLK, Q => n_2335, QN
                           => n42003);
   clk_r_REG12139_S1 : DFF_X1 port map( D => n36523, CK => CLK, Q => n_2336, QN
                           => n42002);
   clk_r_REG13017_S1 : DFF_X1 port map( D => n36524, CK => CLK, Q => n_2337, QN
                           => n42001);
   clk_r_REG12238_S1 : DFF_X1 port map( D => n36526, CK => CLK, Q => n_2338, QN
                           => n42000);
   clk_r_REG12554_S1 : DFF_X1 port map( D => n36527, CK => CLK, Q => n_2339, QN
                           => n41999);
   clk_r_REG12572_S1 : DFF_X1 port map( D => n36528, CK => CLK, Q => n_2340, QN
                           => n41998);
   clk_r_REG12570_S1 : DFF_X1 port map( D => n36529, CK => CLK, Q => n_2341, QN
                           => n41997);
   clk_r_REG12442_S1 : DFF_X1 port map( D => n36530, CK => CLK, Q => n_2342, QN
                           => n41996);
   clk_r_REG12638_S1 : DFF_X1 port map( D => n36531, CK => CLK, Q => n_2343, QN
                           => n41995);
   clk_r_REG12440_S1 : DFF_X1 port map( D => n36532, CK => CLK, Q => n_2344, QN
                           => n41994);
   clk_r_REG12510_S1 : DFF_X1 port map( D => n36533, CK => CLK, Q => n_2345, QN
                           => n41993);
   clk_r_REG13318_S1 : DFF_X1 port map( D => n36534, CK => CLK, Q => n_2346, QN
                           => n41992);
   clk_r_REG13081_S1 : DFF_X1 port map( D => n36536, CK => CLK, Q => n_2347, QN
                           => n41991);
   clk_r_REG13061_S1 : DFF_X1 port map( D => n36537, CK => CLK, Q => n_2348, QN
                           => n41990);
   clk_r_REG12236_S1 : DFF_X1 port map( D => n36539, CK => CLK, Q => n_2349, QN
                           => n41989);
   clk_r_REG12508_S1 : DFF_X1 port map( D => n36540, CK => CLK, Q => n_2350, QN
                           => n41988);
   clk_r_REG12636_S1 : DFF_X1 port map( D => n36541, CK => CLK, Q => n_2351, QN
                           => n41987);
   clk_r_REG12422_S1 : DFF_X1 port map( D => n36542, CK => CLK, Q => n_2352, QN
                           => n41986);
   clk_r_REG12552_S1 : DFF_X1 port map( D => n36544, CK => CLK, Q => n_2353, QN
                           => n41985);
   clk_r_REG12360_S1 : DFF_X1 port map( D => n36545, CK => CLK, Q => n_2354, QN
                           => n41984);
   clk_r_REG12935_S1 : DFF_X1 port map( D => n36546, CK => CLK, Q => n_2355, QN
                           => n41983);
   clk_r_REG12488_S1 : DFF_X1 port map( D => n36547, CK => CLK, Q => n_2356, QN
                           => n41982);
   clk_r_REG13059_S1 : DFF_X1 port map( D => n36548, CK => CLK, Q => n_2357, QN
                           => n41981);
   clk_r_REG12358_S1 : DFF_X1 port map( D => n36549, CK => CLK, Q => n_2358, QN
                           => n41980);
   clk_r_REG12550_S1 : DFF_X1 port map( D => n36551, CK => CLK, Q => n_2359, QN
                           => n41979);
   clk_r_REG13015_S1 : DFF_X1 port map( D => n36552, CK => CLK, Q => n_2360, QN
                           => n41978);
   clk_r_REG12951_S1 : DFF_X1 port map( D => n36553, CK => CLK, Q => n_2361, QN
                           => n41977);
   clk_r_REG12376_S1 : DFF_X1 port map( D => n36554, CK => CLK, Q => n_2362, QN
                           => n41976);
   clk_r_REG12420_S1 : DFF_X1 port map( D => n36555, CK => CLK, Q => n_2363, QN
                           => n41975);
   clk_r_REG12418_S1 : DFF_X1 port map( D => n36556, CK => CLK, Q => n_2364, QN
                           => n41974);
   clk_r_REG12356_S1 : DFF_X1 port map( D => n36557, CK => CLK, Q => n_2365, QN
                           => n41973);
   clk_r_REG12933_S1 : DFF_X1 port map( D => n36558, CK => CLK, Q => n_2366, QN
                           => n41972);
   clk_r_REG12707_S1 : DFF_X1 port map( D => n36559, CK => CLK, Q => n_2367, QN
                           => n41971);
   clk_r_REG12548_S1 : DFF_X1 port map( D => n36560, CK => CLK, Q => n_2368, QN
                           => n41970);
   clk_r_REG12546_S1 : DFF_X1 port map( D => n36561, CK => CLK, Q => n_2369, QN
                           => n41969);
   clk_r_REG12416_S1 : DFF_X1 port map( D => n36562, CK => CLK, Q => n_2370, QN
                           => n41968);
   clk_r_REG12354_S1 : DFF_X1 port map( D => n36563, CK => CLK, Q => n_2371, QN
                           => n41967);
   clk_r_REG12931_S1 : DFF_X1 port map( D => n36564, CK => CLK, Q => n_2372, QN
                           => n41966);
   clk_r_REG12137_S1 : DFF_X1 port map( D => n36565, CK => CLK, Q => n_2373, QN
                           => n41965);
   clk_r_REG12544_S1 : DFF_X1 port map( D => n36566, CK => CLK, Q => n_2374, QN
                           => n41964);
   clk_r_REG12414_S1 : DFF_X1 port map( D => n36567, CK => CLK, Q => n_2375, QN
                           => n41963);
   clk_r_REG12929_S1 : DFF_X1 port map( D => n36568, CK => CLK, Q => n_2376, QN
                           => n41962);
   clk_r_REG12352_S1 : DFF_X1 port map( D => n36569, CK => CLK, Q => n_2377, QN
                           => n41961);
   clk_r_REG12995_S1 : DFF_X1 port map( D => n36570, CK => CLK, Q => n_2378, QN
                           => n41960);
   clk_r_REG11668_S1 : DFF_X1 port map( D => n36571, CK => CLK, Q => n_2379, QN
                           => n41959);
   clk_r_REG12634_S1 : DFF_X1 port map( D => n36573, CK => CLK, Q => n_2380, QN
                           => n41958);
   clk_r_REG12927_S1 : DFF_X1 port map( D => n36574, CK => CLK, Q => n_2381, QN
                           => n41957);
   clk_r_REG12729_S1 : DFF_X1 port map( D => n36575, CK => CLK, Q => n_2382, QN
                           => n41956);
   clk_r_REG12632_S1 : DFF_X1 port map( D => n36576, CK => CLK, Q => n_2383, QN
                           => n41955);
   clk_r_REG12841_S1 : DFF_X1 port map( D => n36577, CK => CLK, Q => n_2384, QN
                           => n41954);
   clk_r_REG12630_S1 : DFF_X1 port map( D => n36578, CK => CLK, Q => n_2385, QN
                           => n41953);
   clk_r_REG13189_S1 : DFF_X1 port map( D => n36580, CK => CLK, Q => n_2386, QN
                           => n41952);
   clk_r_REG12542_S1 : DFF_X1 port map( D => n36581, CK => CLK, Q => n_2387, QN
                           => n41951);
   clk_r_REG12993_S1 : DFF_X1 port map( D => n36582, CK => CLK, Q => n_2388, QN
                           => n41950);
   clk_r_REG11666_S1 : DFF_X1 port map( D => n36583, CK => CLK, Q => n_2389, QN
                           => n41949);
   clk_r_REG12234_S1 : DFF_X1 port map( D => n36585, CK => CLK, Q => n_2390, QN
                           => n41948);
   clk_r_REG12925_S1 : DFF_X1 port map( D => n36587, CK => CLK, Q => n_2391, QN
                           => n41947);
   clk_r_REG12412_S1 : DFF_X1 port map( D => n36588, CK => CLK, Q => n_2392, QN
                           => n41946);
   clk_r_REG12486_S1 : DFF_X1 port map( D => n36589, CK => CLK, Q => n_2393, QN
                           => n41945);
   clk_r_REG13316_S1 : DFF_X1 port map( D => n36590, CK => CLK, Q => n_2394, QN
                           => n41944);
   clk_r_REG12484_S1 : DFF_X1 port map( D => n36591, CK => CLK, Q => n_2395, QN
                           => n41943);
   clk_r_REG12616_S1 : DFF_X1 port map( D => n36592, CK => CLK, Q => n_2396, QN
                           => n41942);
   clk_r_REG11664_S1 : DFF_X1 port map( D => n36593, CK => CLK, Q => n_2397, QN
                           => n41941);
   clk_r_REG12839_S1 : DFF_X1 port map( D => n36594, CK => CLK, Q => n_2398, QN
                           => n41940);
   clk_r_REG13057_S1 : DFF_X1 port map( D => n36595, CK => CLK, Q => n_2399, QN
                           => n41939);
   clk_r_REG12540_S1 : DFF_X1 port map( D => n36596, CK => CLK, Q => n_2400, QN
                           => n41938);
   clk_r_REG12991_S1 : DFF_X1 port map( D => n36597, CK => CLK, Q => n_2401, QN
                           => n41937);
   clk_r_REG12614_S1 : DFF_X1 port map( D => n36598, CK => CLK, Q => n_2402, QN
                           => n41936);
   clk_r_REG12837_S1 : DFF_X1 port map( D => n36599, CK => CLK, Q => n_2403, QN
                           => n41935);
   clk_r_REG11662_S1 : DFF_X1 port map( D => n36600, CK => CLK, Q => n_2404, QN
                           => n41934);
   clk_r_REG12612_S1 : DFF_X1 port map( D => n36601, CK => CLK, Q => n_2405, QN
                           => n41933);
   clk_r_REG13149_S1 : DFF_X1 port map( D => n36602, CK => CLK, Q => n_2406, QN
                           => n41932);
   clk_r_REG12482_S1 : DFF_X1 port map( D => n36603, CK => CLK, Q => n_2407, QN
                           => n41931);
   clk_r_REG12350_S1 : DFF_X1 port map( D => n36604, CK => CLK, Q => n_2408, QN
                           => n41930);
   clk_r_REG12989_S1 : DFF_X1 port map( D => n36605, CK => CLK, Q => n_2409, QN
                           => n41929);
   clk_r_REG12610_S1 : DFF_X1 port map( D => n36607, CK => CLK, Q => n_2410, QN
                           => n41928);
   clk_r_REG13055_S1 : DFF_X1 port map( D => n36608, CK => CLK, Q => n_2411, QN
                           => n41927);
   clk_r_REG12608_S1 : DFF_X1 port map( D => n36610, CK => CLK, Q => n_2412, QN
                           => n41926);
   clk_r_REG11383_S1 : DFF_X1 port map( D => n36611, CK => CLK, Q => n_2413, QN
                           => n41925);
   clk_r_REG12480_S1 : DFF_X1 port map( D => n36612, CK => CLK, Q => n_2414, QN
                           => n41924);
   clk_r_REG13117_S1 : DFF_X1 port map( D => n36613, CK => CLK, Q => n_2415, QN
                           => n41923);
   clk_r_REG12478_S1 : DFF_X1 port map( D => n36614, CK => CLK, Q => n_2416, QN
                           => n41922);
   clk_r_REG13053_S1 : DFF_X1 port map( D => n36615, CK => CLK, Q => n_2417, QN
                           => n41921);
   clk_r_REG13051_S1 : DFF_X1 port map( D => n36616, CK => CLK, Q => n_2418, QN
                           => n41920);
   clk_r_REG12260_S1 : DFF_X1 port map( D => n36617, CK => CLK, Q => n_2419, QN
                           => n41919);
   clk_r_REG13115_S1 : DFF_X1 port map( D => n36619, CK => CLK, Q => n_2420, QN
                           => n41918);
   clk_r_REG12606_S1 : DFF_X1 port map( D => n36620, CK => CLK, Q => n_2421, QN
                           => n41917);
   clk_r_REG12987_S1 : DFF_X1 port map( D => n36621, CK => CLK, Q => n_2422, QN
                           => n41916);
   clk_r_REG11660_S1 : DFF_X1 port map( D => n36622, CK => CLK, Q => n_2423, QN
                           => n41915);
   clk_r_REG11658_S1 : DFF_X1 port map( D => n36623, CK => CLK, Q => n_2424, QN
                           => n41914);
   clk_r_REG12985_S1 : DFF_X1 port map( D => n36624, CK => CLK, Q => n_2425, QN
                           => n41913);
   clk_r_REG11656_S1 : DFF_X1 port map( D => n36625, CK => CLK, Q => n_2426, QN
                           => n41912);
   clk_r_REG11654_S1 : DFF_X1 port map( D => n36626, CK => CLK, Q => n_2427, QN
                           => n41911);
   clk_r_REG13049_S1 : DFF_X1 port map( D => n36627, CK => CLK, Q => n_2428, QN
                           => n41910);
   clk_r_REG12538_S1 : DFF_X1 port map( D => n36628, CK => CLK, Q => n_2429, QN
                           => n41909);
   clk_r_REG12835_S1 : DFF_X1 port map( D => n36629, CK => CLK, Q => n_2430, QN
                           => n41908);
   clk_r_REG12536_S1 : DFF_X1 port map( D => n36630, CK => CLK, Q => n_2431, QN
                           => n41907);
   clk_r_REG12534_S1 : DFF_X1 port map( D => n36631, CK => CLK, Q => n_2432, QN
                           => n41906);
   clk_r_REG12506_S1 : DFF_X1 port map( D => n36632, CK => CLK, Q => n_2433, QN
                           => n41905);
   clk_r_REG12348_S1 : DFF_X1 port map( D => n36633, CK => CLK, Q => n_2434, QN
                           => n41904);
   clk_r_REG12983_S1 : DFF_X1 port map( D => n36634, CK => CLK, Q => n_2435, QN
                           => n41903);
   clk_r_REG12532_S1 : DFF_X1 port map( D => n36635, CK => CLK, Q => n_2436, QN
                           => n41902);
   clk_r_REG13079_S1 : DFF_X1 port map( D => n36636, CK => CLK, Q => n_2437, QN
                           => n41901);
   clk_r_REG12504_S1 : DFF_X1 port map( D => n36637, CK => CLK, Q => n_2438, QN
                           => n41900);
   clk_r_REG12981_S1 : DFF_X1 port map( D => n36639, CK => CLK, Q => n_2439, QN
                           => n41899);
   clk_r_REG13013_S1 : DFF_X1 port map( D => n36640, CK => CLK, Q => n_2440, QN
                           => n41898);
   clk_r_REG12923_S1 : DFF_X1 port map( D => n36641, CK => CLK, Q => n_2441, QN
                           => n41897);
   clk_r_REG13077_S1 : DFF_X1 port map( D => n36642, CK => CLK, Q => n_2442, QN
                           => n41896);
   clk_r_REG10776_S1 : DFF_X1 port map( D => n36644, CK => CLK, Q => n_2443, QN
                           => n41895);
   clk_r_REG12346_S1 : DFF_X1 port map( D => n36645, CK => CLK, Q => n_2444, QN
                           => n41894);
   clk_r_REG13314_S1 : DFF_X1 port map( D => n36646, CK => CLK, Q => n_2445, QN
                           => n41893);
   clk_r_REG12410_S1 : DFF_X1 port map( D => n36647, CK => CLK, Q => n_2446, QN
                           => n41892);
   clk_r_REG12604_S1 : DFF_X1 port map( D => n36648, CK => CLK, Q => n_2447, QN
                           => n41891);
   clk_r_REG13011_S1 : DFF_X1 port map( D => n36649, CK => CLK, Q => n_2448, QN
                           => n41890);
   clk_r_REG13009_S1 : DFF_X1 port map( D => n36650, CK => CLK, Q => n_2449, QN
                           => n41889);
   clk_r_REG13007_S1 : DFF_X1 port map( D => n36651, CK => CLK, Q => n_2450, QN
                           => n41888);
   clk_r_REG12602_S1 : DFF_X1 port map( D => n36652, CK => CLK, Q => n_2451, QN
                           => n41887);
   clk_r_REG13312_S1 : DFF_X1 port map( D => n36653, CK => CLK, Q => n_2452, QN
                           => n41886);
   clk_r_REG11381_S1 : DFF_X1 port map( D => n36654, CK => CLK, Q => n_2453, QN
                           => n41885);
   clk_r_REG12502_S1 : DFF_X1 port map( D => n36655, CK => CLK, Q => n_2454, QN
                           => n41884);
   clk_r_REG12344_S1 : DFF_X1 port map( D => n36656, CK => CLK, Q => n_2455, QN
                           => n41883);
   clk_r_REG12342_S1 : DFF_X1 port map( D => n36657, CK => CLK, Q => n_2456, QN
                           => n41882);
   clk_r_REG12979_S1 : DFF_X1 port map( D => n36658, CK => CLK, Q => n_2457, QN
                           => n41881);
   clk_r_REG12500_S1 : DFF_X1 port map( D => n36659, CK => CLK, Q => n_2458, QN
                           => n41880);
   clk_r_REG12498_S1 : DFF_X1 port map( D => n36660, CK => CLK, Q => n_2459, QN
                           => n41879);
   clk_r_REG11379_S1 : DFF_X1 port map( D => n36661, CK => CLK, Q => n_2460, QN
                           => n41878);
   clk_r_REG10481_S1 : DFF_X1 port map( D => n36663, CK => CLK, Q => n_2461, QN
                           => n41877);
   clk_r_REG12600_S1 : DFF_X1 port map( D => n36664, CK => CLK, Q => n_2462, QN
                           => n41876);
   clk_r_REG12476_S1 : DFF_X1 port map( D => n36665, CK => CLK, Q => n_2463, QN
                           => n41875);
   clk_r_REG12039_S1 : DFF_X1 port map( D => n36666, CK => CLK, Q => n_2464, QN
                           => n41874);
   clk_r_REG12949_S1 : DFF_X1 port map( D => n36667, CK => CLK, Q => n_2465, QN
                           => n41873);
   clk_r_REG11377_S1 : DFF_X1 port map( D => n36668, CK => CLK, Q => n_2466, QN
                           => n41872);
   clk_r_REG12921_S1 : DFF_X1 port map( D => n36669, CK => CLK, Q => n_2467, QN
                           => n41871);
   clk_r_REG13310_S1 : DFF_X1 port map( D => n36670, CK => CLK, Q => n_2468, QN
                           => n41870);
   clk_r_REG12408_S1 : DFF_X1 port map( D => n36671, CK => CLK, Q => n_2469, QN
                           => n41869);
   clk_r_REG12919_S1 : DFF_X1 port map( D => n36672, CK => CLK, Q => n_2470, QN
                           => n41868);
   clk_r_REG13075_S1 : DFF_X1 port map( D => n36673, CK => CLK, Q => n_2471, QN
                           => n41867);
   clk_r_REG10839_S1 : DFF_X1 port map( D => n36675, CK => CLK, Q => n_2472, QN
                           => n41866);
   clk_r_REG12037_S1 : DFF_X1 port map( D => n36678, CK => CLK, Q => n_2473, QN
                           => n41865);
   clk_r_REG12496_S1 : DFF_X1 port map( D => n36679, CK => CLK, Q => n_2474, QN
                           => n41864);
   clk_r_REG12598_S1 : DFF_X1 port map( D => n36680, CK => CLK, Q => n_2475, QN
                           => n41863);
   clk_r_REG12406_S1 : DFF_X1 port map( D => n36681, CK => CLK, Q => n_2476, QN
                           => n41862);
   clk_r_REG12404_S1 : DFF_X1 port map( D => n36682, CK => CLK, Q => n_2477, QN
                           => n41861);
   clk_r_REG10343_S1 : DFF_X1 port map( D => n36684, CK => CLK, Q => n_2478, QN
                           => n41860);
   clk_r_REG12833_S1 : DFF_X1 port map( D => n36685, CK => CLK, Q => n_2479, QN
                           => n41859);
   clk_r_REG12402_S1 : DFF_X1 port map( D => n36686, CK => CLK, Q => n_2480, QN
                           => n41858);
   clk_r_REG13047_S1 : DFF_X1 port map( D => n36688, CK => CLK, Q => n_2481, QN
                           => n41857);
   clk_r_REG13045_S1 : DFF_X1 port map( D => n36689, CK => CLK, Q => n_2482, QN
                           => n41856);
   clk_r_REG12917_S1 : DFF_X1 port map( D => n36690, CK => CLK, Q => n_2483, QN
                           => n41855);
   clk_r_REG12705_S1 : DFF_X1 port map( D => n36691, CK => CLK, Q => n_2484, QN
                           => n41854);
   clk_r_REG12296_S1 : DFF_X1 port map( D => n36693, CK => CLK, Q => n_2485, QN
                           => n41853);
   clk_r_REG12915_S1 : DFF_X1 port map( D => n36695, CK => CLK, Q => n_2486, QN
                           => n41852);
   clk_r_REG13043_S1 : DFF_X1 port map( D => n36697, CK => CLK, Q => n_2487, QN
                           => n41851);
   clk_r_REG13041_S1 : DFF_X1 port map( D => n36699, CK => CLK, Q => n_2488, QN
                           => n41850);
   clk_r_REG10301_S1 : DFF_X1 port map( D => n36702, CK => CLK, Q => n_2489, QN
                           => n41849);
   clk_r_REG12596_S1 : DFF_X1 port map( D => n36704, CK => CLK, Q => n_2490, QN
                           => n41848);
   clk_r_REG13308_S1 : DFF_X1 port map( D => n36706, CK => CLK, Q => n_2491, QN
                           => n41847);
   clk_r_REG12135_S1 : DFF_X1 port map( D => n36707, CK => CLK, Q => n_2492, QN
                           => n41846);
   clk_r_REG13306_S1 : DFF_X1 port map( D => n36709, CK => CLK, Q => n_2493, QN
                           => n41845);
   clk_r_REG12977_S1 : DFF_X1 port map( D => n36711, CK => CLK, Q => n_2494, QN
                           => n41844);
   clk_r_REG10541_S1 : DFF_X1 port map( D => n36713, CK => CLK, Q => n_2495, QN
                           => n41843);
   clk_r_REG10390_S1 : DFF_X1 port map( D => n36716, CK => CLK, Q => n_2496, QN
                           => n41842);
   clk_r_REG10308_S1 : DFF_X1 port map( D => n36719, CK => CLK, Q => n_2497, QN
                           => n41841);
   clk_r_REG12594_S1 : DFF_X1 port map( D => n36720, CK => CLK, Q => n_2498, QN
                           => n41840);
   clk_r_REG12374_S1 : DFF_X1 port map( D => n36721, CK => CLK, Q => n_2499, QN
                           => n41839);
   clk_r_REG12372_S1 : DFF_X1 port map( D => n36722, CK => CLK, Q => n_2500, QN
                           => n41838);
   clk_r_REG12628_S1 : DFF_X1 port map( D => n36723, CK => CLK, Q => n_2501, QN
                           => n41837);
   clk_r_REG12370_S1 : DFF_X1 port map( D => n36724, CK => CLK, Q => n_2502, QN
                           => n41836);
   clk_r_REG12530_S1 : DFF_X1 port map( D => n36725, CK => CLK, Q => n_2503, QN
                           => n41835);
   clk_r_REG12592_S1 : DFF_X1 port map( D => n36727, CK => CLK, Q => n_2504, QN
                           => n41834);
   clk_r_REG12801_S1 : DFF_X1 port map( D => n36728, CK => CLK, Q => n_2505, QN
                           => n41833);
   clk_r_REG12590_S1 : DFF_X1 port map( D => n36729, CK => CLK, Q => n_2506, QN
                           => n41832);
   clk_r_REG10404_S1 : DFF_X1 port map( D => n36731, CK => CLK, Q => n_2507, QN
                           => n41831);
   clk_r_REG13039_S1 : DFF_X1 port map( D => n36732, CK => CLK, Q => n_2508, QN
                           => n41830);
   clk_r_REG12947_S1 : DFF_X1 port map( D => n36733, CK => CLK, Q => n_2509, QN
                           => n41829);
   clk_r_REG12799_S1 : DFF_X1 port map( D => n36734, CK => CLK, Q => n_2510, QN
                           => n41828);
   clk_r_REG12438_S1 : DFF_X1 port map( D => n36735, CK => CLK, Q => n_2511, QN
                           => n41827);
   clk_r_REG12975_S1 : DFF_X1 port map( D => n36737, CK => CLK, Q => n_2512, QN
                           => n41826);
   clk_r_REG13037_S1 : DFF_X1 port map( D => n36738, CK => CLK, Q => n_2513, QN
                           => n41825);
   clk_r_REG12474_S1 : DFF_X1 port map( D => n36739, CK => CLK, Q => n_2514, QN
                           => n41824);
   clk_r_REG13035_S1 : DFF_X1 port map( D => n36740, CK => CLK, Q => n_2515, QN
                           => n41823);
   clk_r_REG13033_S1 : DFF_X1 port map( D => n36741, CK => CLK, Q => n_2516, QN
                           => n41822);
   clk_r_REG12472_S1 : DFF_X1 port map( D => n36742, CK => CLK, Q => n_2517, QN
                           => n41821);
   clk_r_REG12528_S1 : DFF_X1 port map( D => n36743, CK => CLK, Q => n_2518, QN
                           => n41820);
   clk_r_REG13031_S1 : DFF_X1 port map( D => n36744, CK => CLK, Q => n_2519, QN
                           => n41819);
   clk_r_REG12470_S1 : DFF_X1 port map( D => n36745, CK => CLK, Q => n_2520, QN
                           => n41818);
   clk_r_REG12626_S1 : DFF_X1 port map( D => n36746, CK => CLK, Q => n_2521, QN
                           => n41817);
   clk_r_REG11940_S1 : DFF_X1 port map( D => n36747, CK => CLK, Q => n_2522, QN
                           => n41816);
   clk_r_REG10635_S1 : DFF_X1 port map( D => n36749, CK => CLK, Q => n_2523, QN
                           => n41815);
   clk_r_REG12727_S1 : DFF_X1 port map( D => n36750, CK => CLK, Q => n_2524, QN
                           => n41814);
   clk_r_REG12725_S1 : DFF_X1 port map( D => n36752, CK => CLK, Q => n_2525, QN
                           => n41813);
   clk_r_REG12436_S1 : DFF_X1 port map( D => n36753, CK => CLK, Q => n_2526, QN
                           => n41812);
   clk_r_REG12973_S1 : DFF_X1 port map( D => n36754, CK => CLK, Q => n_2527, QN
                           => n41811);
   clk_r_REG12568_S1 : DFF_X1 port map( D => n36755, CK => CLK, Q => n_2528, QN
                           => n41810);
   clk_r_REG12133_S1 : DFF_X1 port map( D => n36756, CK => CLK, Q => n_2529, QN
                           => n41809);
   clk_r_REG12468_S1 : DFF_X1 port map( D => n36757, CK => CLK, Q => n_2530, QN
                           => n41808);
   clk_r_REG12434_S1 : DFF_X1 port map( D => n36758, CK => CLK, Q => n_2531, QN
                           => n41807);
   clk_r_REG12588_S1 : DFF_X1 port map( D => n36759, CK => CLK, Q => n_2532, QN
                           => n41806);
   clk_r_REG13029_S1 : DFF_X1 port map( D => n36760, CK => CLK, Q => n_2533, QN
                           => n41805);
   clk_r_REG12566_S1 : DFF_X1 port map( D => n36761, CK => CLK, Q => n_2534, QN
                           => n41804);
   clk_r_REG13005_S1 : DFF_X1 port map( D => n36762, CK => CLK, Q => n_2535, QN
                           => n41803);
   clk_r_REG12432_S1 : DFF_X1 port map( D => n36763, CK => CLK, Q => n_2536, QN
                           => n41802);
   clk_r_REG12564_S1 : DFF_X1 port map( D => n36764, CK => CLK, Q => n_2537, QN
                           => n41801);
   clk_r_REG12466_S1 : DFF_X1 port map( D => n36765, CK => CLK, Q => n_2538, QN
                           => n41800);
   clk_r_REG12464_S1 : DFF_X1 port map( D => n36766, CK => CLK, Q => n_2539, QN
                           => n41799);
   clk_r_REG13003_S1 : DFF_X1 port map( D => n36767, CK => CLK, Q => n_2540, QN
                           => n41798);
   clk_r_REG12971_S1 : DFF_X1 port map( D => n36768, CK => CLK, Q => n_2541, QN
                           => n41797);
   clk_r_REG12945_S1 : DFF_X1 port map( D => n36769, CK => CLK, Q => n_2542, QN
                           => n41796);
   clk_r_REG12913_S1 : DFF_X1 port map( D => n36770, CK => CLK, Q => n_2543, QN
                           => n41795);
   clk_r_REG12911_S1 : DFF_X1 port map( D => n36771, CK => CLK, Q => n_2544, QN
                           => n41794);
   clk_r_REG13027_S1 : DFF_X1 port map( D => n36772, CK => CLK, Q => n_2545, QN
                           => n41793);
   clk_r_REG13025_S1 : DFF_X1 port map( D => n36773, CK => CLK, Q => n_2546, QN
                           => n41792);
   clk_r_REG12462_S1 : DFF_X1 port map( D => n36774, CK => CLK, Q => n_2547, QN
                           => n41791);
   clk_r_REG12494_S1 : DFF_X1 port map( D => n36775, CK => CLK, Q => n_2548, QN
                           => n41790);
   clk_r_REG12562_S1 : DFF_X1 port map( D => n36776, CK => CLK, Q => n_2549, QN
                           => n41789);
   clk_r_REG12969_S1 : DFF_X1 port map( D => n36777, CK => CLK, Q => n_2550, QN
                           => n41788);
   clk_r_REG12340_S1 : DFF_X1 port map( D => n36778, CK => CLK, Q => n_2551, QN
                           => n41787);
   clk_r_REG12430_S1 : DFF_X1 port map( D => n36779, CK => CLK, Q => n_2552, QN
                           => n41786);
   clk_r_REG12967_S1 : DFF_X1 port map( D => n36780, CK => CLK, Q => n_2553, QN
                           => n41785);
   clk_r_REG12428_S1 : DFF_X1 port map( D => n36781, CK => CLK, Q => n_2554, QN
                           => n41784);
   clk_r_REG12338_S1 : DFF_X1 port map( D => n36782, CK => CLK, Q => n_2555, QN
                           => n41783);
   clk_r_REG10522_S1 : DFF_X1 port map( D => n36784, CK => CLK, Q => n_2556, QN
                           => n41782);
   clk_r_REG12368_S1 : DFF_X1 port map( D => n36785, CK => CLK, Q => n_2557, QN
                           => n41781);
   clk_r_REG12336_S1 : DFF_X1 port map( D => n36786, CK => CLK, Q => n_2558, QN
                           => n41780);
   clk_r_REG12909_S1 : DFF_X1 port map( D => n36787, CK => CLK, Q => n_2559, QN
                           => n41779);
   clk_r_REG12797_S1 : DFF_X1 port map( D => n36789, CK => CLK, Q => n_2560, QN
                           => n41778);
   clk_r_REG12943_S1 : DFF_X1 port map( D => n36790, CK => CLK, Q => n_2561, QN
                           => n41777);
   clk_r_REG12586_S1 : DFF_X1 port map( D => n36791, CK => CLK, Q => n_2562, QN
                           => n41776);
   clk_r_REG12334_S1 : DFF_X1 port map( D => n36792, CK => CLK, Q => n_2563, QN
                           => n41775);
   clk_r_REG12941_S1 : DFF_X1 port map( D => n36793, CK => CLK, Q => n_2564, QN
                           => n41774);
   clk_r_REG12526_S1 : DFF_X1 port map( D => n36794, CK => CLK, Q => n_2565, QN
                           => n41773);
   clk_r_REG12426_S1 : DFF_X1 port map( D => n36795, CK => CLK, Q => n_2566, QN
                           => n41772);
   clk_r_REG12400_S1 : DFF_X1 port map( D => n36796, CK => CLK, Q => n_2567, QN
                           => n41771);
   clk_r_REG12560_S1 : DFF_X1 port map( D => n36797, CK => CLK, Q => n_2568, QN
                           => n41770);
   clk_r_REG12939_S1 : DFF_X1 port map( D => n36798, CK => CLK, Q => n_2569, QN
                           => n41769);
   clk_r_REG12584_S1 : DFF_X1 port map( D => n36800, CK => CLK, Q => n_2570, QN
                           => n41768);
   clk_r_REG13073_S1 : DFF_X1 port map( D => n36802, CK => CLK, Q => n_2571, QN
                           => n41767);
   clk_r_REG13071_S1 : DFF_X1 port map( D => n36804, CK => CLK, Q => n_2572, QN
                           => n41766);
   clk_r_REG13069_S1 : DFF_X1 port map( D => n36806, CK => CLK, Q => n_2573, QN
                           => n41765);
   clk_r_REG13023_S1 : DFF_X1 port map( D => n36808, CK => CLK, Q => n_2574, QN
                           => n41764);
   clk_r_REG12460_S1 : DFF_X1 port map( D => n36809, CK => CLK, Q => n_2575, QN
                           => n41763);
   clk_r_REG12458_S1 : DFF_X1 port map( D => n36810, CK => CLK, Q => n_2576, QN
                           => n41762);
   clk_r_REG12332_S1 : DFF_X1 port map( D => n36812, CK => CLK, Q => n_2577, QN
                           => n41761);
   clk_r_REG12456_S1 : DFF_X1 port map( D => n36814, CK => CLK, Q => n_2578, QN
                           => n41760);
   clk_r_REG12330_S1 : DFF_X1 port map( D => n36815, CK => CLK, Q => n_2579, QN
                           => n41759);
   clk_r_REG12454_S1 : DFF_X1 port map( D => n36816, CK => CLK, Q => n_2580, QN
                           => n41758);
   clk_r_REG13021_S1 : DFF_X1 port map( D => n36817, CK => CLK, Q => n_2581, QN
                           => n41757);
   clk_r_REG12398_S1 : DFF_X1 port map( D => n36818, CK => CLK, Q => n_2582, QN
                           => n41756);
   clk_r_REG12396_S1 : DFF_X1 port map( D => n36819, CK => CLK, Q => n_2583, QN
                           => n41755);
   clk_r_REG12907_S1 : DFF_X1 port map( D => n36820, CK => CLK, Q => n_2584, QN
                           => n41754);
   clk_r_REG12905_S1 : DFF_X1 port map( D => n36821, CK => CLK, Q => n_2585, QN
                           => n41753);
   clk_r_REG12328_S1 : DFF_X1 port map( D => n36822, CK => CLK, Q => n_2586, QN
                           => n41752);
   clk_r_REG12326_S1 : DFF_X1 port map( D => n36823, CK => CLK, Q => n_2587, QN
                           => n41751);
   clk_r_REG12394_S1 : DFF_X1 port map( D => n36824, CK => CLK, Q => n_2588, QN
                           => n41750);
   clk_r_REG12392_S1 : DFF_X1 port map( D => n36825, CK => CLK, Q => n_2589, QN
                           => n41749);
   clk_r_REG12324_S1 : DFF_X1 port map( D => n36826, CK => CLK, Q => n_2590, QN
                           => n41748);
   clk_r_REG12903_S1 : DFF_X1 port map( D => n36827, CK => CLK, Q => n_2591, QN
                           => n41747);
   clk_r_REG12901_S1 : DFF_X1 port map( D => n36828, CK => CLK, Q => n_2592, QN
                           => n41746);
   clk_r_REG12524_S1 : DFF_X1 port map( D => n36829, CK => CLK, Q => n_2593, QN
                           => n41745);
   clk_r_REG12899_S1 : DFF_X1 port map( D => n36830, CK => CLK, Q => n_2594, QN
                           => n41744);
   clk_r_REG12390_S1 : DFF_X1 port map( D => n36831, CK => CLK, Q => n_2595, QN
                           => n41743);
   clk_r_REG12965_S1 : DFF_X1 port map( D => n36832, CK => CLK, Q => n_2596, QN
                           => n41742);
   clk_r_REG12582_S1 : DFF_X1 port map( D => n36834, CK => CLK, Q => n_2597, QN
                           => n41741);
   clk_r_REG12897_S1 : DFF_X1 port map( D => n36836, CK => CLK, Q => n_2598, QN
                           => n41740);
   clk_r_REG13067_S1 : DFF_X1 port map( D => n36837, CK => CLK, Q => n_2599, QN
                           => n41739);
   clk_r_REG12963_S1 : DFF_X1 port map( D => n36838, CK => CLK, Q => n_2600, QN
                           => n41738);
   clk_r_REG12322_S1 : DFF_X1 port map( D => n36839, CK => CLK, Q => n_2601, QN
                           => n41737);
   clk_r_REG12452_S1 : DFF_X1 port map( D => n36840, CK => CLK, Q => n_2602, QN
                           => n41736);
   clk_r_REG12388_S1 : DFF_X1 port map( D => n36841, CK => CLK, Q => n_2603, QN
                           => n41735);
   clk_r_REG12492_S1 : DFF_X1 port map( D => n36842, CK => CLK, Q => n_2604, QN
                           => n41734);
   clk_r_REG13065_S1 : DFF_X1 port map( D => n36843, CK => CLK, Q => n_2605, QN
                           => n41733);
   clk_r_REG12450_S1 : DFF_X1 port map( D => n36844, CK => CLK, Q => n_2606, QN
                           => n41732);
   clk_r_REG12522_S1 : DFF_X1 port map( D => n36845, CK => CLK, Q => n_2607, QN
                           => n41731);
   clk_r_REG12520_S1 : DFF_X1 port map( D => n36846, CK => CLK, Q => n_2608, QN
                           => n41730);
   clk_r_REG12624_S1 : DFF_X1 port map( D => n36847, CK => CLK, Q => n_2609, QN
                           => n41729);
   clk_r_REG12961_S1 : DFF_X1 port map( D => n36848, CK => CLK, Q => n_2610, QN
                           => n41728);
   clk_r_REG12959_S1 : DFF_X1 port map( D => n36849, CK => CLK, Q => n_2611, QN
                           => n41727);
   clk_r_REG12518_S1 : DFF_X1 port map( D => n36850, CK => CLK, Q => n_2612, QN
                           => n41726);
   clk_r_REG10358_S1 : DFF_X1 port map( D => n36852, CK => CLK, Q => n_2613, QN
                           => n41725);
   clk_r_REG12580_S1 : DFF_X1 port map( D => n36853, CK => CLK, Q => n_2614, QN
                           => n41724);
   clk_r_REG12957_S1 : DFF_X1 port map( D => n36854, CK => CLK, Q => n_2615, QN
                           => n41723);
   clk_r_REG13001_S1 : DFF_X1 port map( D => n36856, CK => CLK, Q => n_2616, QN
                           => n41722);
   clk_r_REG12490_S1 : DFF_X1 port map( D => n36858, CK => CLK, Q => n_2617, QN
                           => n41721);
   clk_r_REG12999_S1 : DFF_X1 port map( D => n36859, CK => CLK, Q => n_2618, QN
                           => n41720);
   clk_r_REG12516_S1 : DFF_X1 port map( D => n36860, CK => CLK, Q => n_2619, QN
                           => n41719);
   clk_r_REG12386_S1 : DFF_X1 port map( D => n36861, CK => CLK, Q => n_2620, QN
                           => n41718);
   clk_r_REG12622_S1 : DFF_X1 port map( D => n36862, CK => CLK, Q => n_2621, QN
                           => n41717);
   clk_r_REG10456_S1 : DFF_X1 port map( D => n36864, CK => CLK, Q => n_2622, QN
                           => n41716);
   clk_r_REG12895_S1 : DFF_X1 port map( D => n36865, CK => CLK, Q => n_2623, QN
                           => n41715);
   clk_r_REG12937_S1 : DFF_X1 port map( D => n36867, CK => CLK, Q => n_2624, QN
                           => n41714);
   clk_r_REG12620_S1 : DFF_X1 port map( D => n36868, CK => CLK, Q => n_2625, QN
                           => n41713);
   clk_r_REG12366_S1 : DFF_X1 port map( D => n36869, CK => CLK, Q => n_2626, QN
                           => n41712);
   clk_r_REG12618_S1 : DFF_X1 port map( D => n36871, CK => CLK, Q => n_2627, QN
                           => n41711);
   clk_r_REG10463_S1 : DFF_X1 port map( D => n36873, CK => CLK, Q => n_2628, QN
                           => n41710);
   clk_r_REG12514_S1 : DFF_X1 port map( D => n36874, CK => CLK, Q => n_2629, QN
                           => n41709);
   clk_r_REG10449_S1 : DFF_X1 port map( D => n36876, CK => CLK, Q => n_2630, QN
                           => n41708);
   clk_r_REG12558_S1 : DFF_X1 port map( D => n36877, CK => CLK, Q => n_2631, QN
                           => n41707);
   clk_r_REG12364_S1 : DFF_X1 port map( D => n36879, CK => CLK, Q => n_2632, QN
                           => n41706);
   clk_r_REG10377_S1 : DFF_X1 port map( D => n36881, CK => CLK, Q => n_2633, QN
                           => n41705);
   clk_r_REG12997_S1 : DFF_X1 port map( D => n36883, CK => CLK, Q => n_2634, QN
                           => n41704);
   clk_r_REG10367_S1 : DFF_X1 port map( D => n36885, CK => CLK, Q => n_2635, QN
                           => n41703);
   clk_r_REG12578_S1 : DFF_X1 port map( D => n36886, CK => CLK, Q => n_2636, QN
                           => n41702);
   clk_r_REG10470_S1 : DFF_X1 port map( D => n36888, CK => CLK, Q => n_2637, QN
                           => n41701);
   clk_r_REG10440_S1 : DFF_X1 port map( D => n36890, CK => CLK, Q => n_2638, QN
                           => n41700);
   clk_r_REG13063_S1 : DFF_X1 port map( D => n36893, CK => CLK, Q => n_2639, QN
                           => n41699);
   clk_r_REG12424_S1 : DFF_X1 port map( D => n36895, CK => CLK, Q => n_2640, QN
                           => n41698);
   clk_r_REG12556_S1 : DFF_X1 port map( D => n36897, CK => CLK, Q => n_2641, QN
                           => n41697);
   clk_r_REG13469_S2 : DFFS_X1 port map( D => n1526, CK => CLK, SN => RESET_BAR
                           , Q => n_2642, QN => n47504);
   clk_r_REG13465_S2 : DFFS_X1 port map( D => n1525, CK => CLK, SN => RESET_BAR
                           , Q => n_2643, QN => n47505);
   clk_r_REG13472_S4 : DFFS_X1 port map( D => n47494, CK => CLK, SN => 
                           RESET_BAR, Q => n41694, QN => n_2644);
   clk_r_REG11825_S1 : DFF_X1 port map( D => n35853, CK => CLK, Q => n41693, QN
                           => n_2645);
   clk_r_REG13613_S7 : DFFR_X1 port map( D => n31164, CK => CLK, RN => 
                           RESET_BAR, Q => n41692, QN => n_2646);
   clk_r_REG13579_S7 : DFFR_X1 port map( D => n31168, CK => CLK, RN => 
                           RESET_BAR, Q => n41691, QN => n_2647);
   clk_r_REG13218_S1 : DFF_X1 port map( D => n36501, CK => CLK, Q => n41685, QN
                           => n_2648);
   clk_r_REG11486_S1 : DFF_X1 port map( D => n36033, CK => CLK, Q => n41684, QN
                           => n_2649);
   clk_r_REG11480_S1 : DFF_X1 port map( D => n36266, CK => CLK, Q => n41683, QN
                           => n_2650);
   clk_r_REG11472_S1 : DFF_X1 port map( D => n36297, CK => CLK, Q => n41682, QN
                           => n_2651);
   clk_r_REG11478_S1 : DFF_X1 port map( D => n36267, CK => CLK, Q => n41681, QN
                           => n_2652);
   clk_r_REG12651_S1 : DFF_X1 port map( D => n36268, CK => CLK, Q => n41680, QN
                           => n_2653);
   clk_r_REG11476_S1 : DFF_X1 port map( D => n36269, CK => CLK, Q => n41679, QN
                           => n_2654);
   clk_r_REG11474_S1 : DFF_X1 port map( D => n36270, CK => CLK, Q => n41678, QN
                           => n_2655);
   clk_r_REG11292_S1 : DFF_X1 port map( D => n36271, CK => CLK, Q => n41677, QN
                           => n_2656);
   clk_r_REG12683_S1 : DFF_X1 port map( D => n36034, CK => CLK, Q => n41676, QN
                           => n_2657);
   clk_r_REG11589_S1 : DFF_X1 port map( D => n36272, CK => CLK, Q => n41675, QN
                           => n_2658);
   clk_r_REG11484_S1 : DFF_X1 port map( D => n36039, CK => CLK, Q => n41674, QN
                           => n_2659);
   clk_r_REG12669_S1 : DFF_X1 port map( D => n36273, CK => CLK, Q => n41673, QN
                           => n_2660);
   clk_r_REG11735_S1 : DFF_X1 port map( D => n36274, CK => CLK, Q => n41672, QN
                           => n_2661);
   clk_r_REG11785_S1 : DFF_X1 port map( D => n36040, CK => CLK, Q => n41671, QN
                           => n_2662);
   clk_r_REG11890_S1 : DFF_X1 port map( D => n36060, CK => CLK, Q => n41670, QN
                           => n_2663);
   clk_r_REG11482_S1 : DFF_X1 port map( D => n36065, CK => CLK, Q => n41669, QN
                           => n_2664);
   clk_r_REG11775_S1 : DFF_X1 port map( D => n36275, CK => CLK, Q => n41668, QN
                           => n_2665);
   clk_r_REG11452_S1 : DFF_X1 port map( D => n36276, CK => CLK, Q => n41667, QN
                           => n_2666);
   clk_r_REG11773_S1 : DFF_X1 port map( D => n36277, CK => CLK, Q => n41666, QN
                           => n_2667);
   clk_r_REG11771_S1 : DFF_X1 port map( D => n36278, CK => CLK, Q => n41665, QN
                           => n_2668);
   clk_r_REG11470_S1 : DFF_X1 port map( D => n36073, CK => CLK, Q => n41664, QN
                           => n_2669);
   clk_r_REG12667_S1 : DFF_X1 port map( D => n36279, CK => CLK, Q => n41663, QN
                           => n_2670);
   clk_r_REG12679_S1 : DFF_X1 port map( D => n36078, CK => CLK, Q => n41662, QN
                           => n_2671);
   clk_r_REG12665_S1 : DFF_X1 port map( D => n36281, CK => CLK, Q => n41661, QN
                           => n_2672);
   clk_r_REG11783_S1 : DFF_X1 port map( D => n36074, CK => CLK, Q => n41660, QN
                           => n_2673);
   clk_r_REG11781_S1 : DFF_X1 port map( D => n36081, CK => CLK, Q => n41659, QN
                           => n_2674);
   clk_r_REG12677_S1 : DFF_X1 port map( D => n36082, CK => CLK, Q => n41658, QN
                           => n_2675);
   clk_r_REG11769_S1 : DFF_X1 port map( D => n36283, CK => CLK, Q => n41657, QN
                           => n_2676);
   clk_r_REG11513_S1 : DFF_X1 port map( D => n36284, CK => CLK, Q => n41656, QN
                           => n_2677);
   clk_r_REG11450_S1 : DFF_X1 port map( D => n36285, CK => CLK, Q => n41655, QN
                           => n_2678);
   clk_r_REG12681_S1 : DFF_X1 port map( D => n36072, CK => CLK, Q => n41654, QN
                           => n_2679);
   clk_r_REG12663_S1 : DFF_X1 port map( D => n36069, CK => CLK, Q => n41653, QN
                           => n_2680);
   clk_r_REG12649_S1 : DFF_X1 port map( D => n36286, CK => CLK, Q => n41652, QN
                           => n_2681);
   clk_r_REG12647_S1 : DFF_X1 port map( D => n36287, CK => CLK, Q => n41651, QN
                           => n_2682);
   clk_r_REG11559_S1 : DFF_X1 port map( D => n36289, CK => CLK, Q => n41650, QN
                           => n_2683);
   clk_r_REG11340_S1 : DFF_X1 port map( D => n36290, CK => CLK, Q => n41649, QN
                           => n_2684);
   clk_r_REG12645_S1 : DFF_X1 port map( D => n36291, CK => CLK, Q => n41648, QN
                           => n_2685);
   clk_r_REG11641_S1 : DFF_X1 port map( D => n36077, CK => CLK, Q => n41647, QN
                           => n_2686);
   clk_r_REG11346_S1 : DFF_X1 port map( D => n36075, CK => CLK, Q => n41646, QN
                           => n_2687);
   clk_r_REG11567_S1 : DFF_X1 port map( D => n36051, CK => CLK, Q => n41645, QN
                           => n_2688);
   clk_r_REG11557_S1 : DFF_X1 port map( D => n36294, CK => CLK, Q => n41644, QN
                           => n_2689);
   clk_r_REG11639_S1 : DFF_X1 port map( D => n36298, CK => CLK, Q => n41643, QN
                           => n_2690);
   clk_r_REG11555_S1 : DFF_X1 port map( D => n36299, CK => CLK, Q => n41642, QN
                           => n_2691);
   clk_r_REG11553_S1 : DFF_X1 port map( D => n36300, CK => CLK, Q => n41641, QN
                           => n_2692);
   clk_r_REG11926_S1 : DFF_X1 port map( D => n36301, CK => CLK, Q => n41640, QN
                           => n_2693);
   clk_r_REG11565_S1 : DFF_X1 port map( D => n36070, CK => CLK, Q => n41639, QN
                           => n_2694);
   clk_r_REG11924_S1 : DFF_X1 port map( D => n36302, CK => CLK, Q => n41638, QN
                           => n_2695);
   clk_r_REG11551_S1 : DFF_X1 port map( D => n36304, CK => CLK, Q => n41637, QN
                           => n_2696);
   clk_r_REG11338_S1 : DFF_X1 port map( D => n36305, CK => CLK, Q => n41636, QN
                           => n_2697);
   clk_r_REG11637_S1 : DFF_X1 port map( D => n36306, CK => CLK, Q => n41635, QN
                           => n_2698);
   clk_r_REG11531_S1 : DFF_X1 port map( D => n36046, CK => CLK, Q => n41634, QN
                           => n_2699);
   clk_r_REG11527_S1 : DFF_X1 port map( D => n36067, CK => CLK, Q => n41633, QN
                           => n_2700);
   clk_r_REG11733_S1 : DFF_X1 port map( D => n36307, CK => CLK, Q => n41632, QN
                           => n_2701);
   clk_r_REG11529_S1 : DFF_X1 port map( D => n36063, CK => CLK, Q => n41631, QN
                           => n_2702);
   clk_r_REG11922_S1 : DFF_X1 port map( D => n36308, CK => CLK, Q => n41630, QN
                           => n_2703);
   clk_r_REG11511_S1 : DFF_X1 port map( D => n36311, CK => CLK, Q => n41629, QN
                           => n_2704);
   clk_r_REG11932_S1 : DFF_X1 port map( D => n36062, CK => CLK, Q => n41628, QN
                           => n_2705);
   clk_r_REG11749_S1 : DFF_X1 port map( D => n36057, CK => CLK, Q => n41627, QN
                           => n_2706);
   clk_r_REG11643_S1 : DFF_X1 port map( D => n36056, CK => CLK, Q => n41626, QN
                           => n_2707);
   clk_r_REG11336_S1 : DFF_X1 port map( D => n36312, CK => CLK, Q => n41625, QN
                           => n_2708);
   clk_r_REG11334_S1 : DFF_X1 port map( D => n36313, CK => CLK, Q => n41624, QN
                           => n_2709);
   clk_r_REG11332_S1 : DFF_X1 port map( D => n36314, CK => CLK, Q => n41623, QN
                           => n_2710);
   clk_r_REG11330_S1 : DFF_X1 port map( D => n36316, CK => CLK, Q => n41622, QN
                           => n_2711);
   clk_r_REG11635_S1 : DFF_X1 port map( D => n36317, CK => CLK, Q => n41621, QN
                           => n_2712);
   clk_r_REG11633_S1 : DFF_X1 port map( D => n36318, CK => CLK, Q => n41620, QN
                           => n_2713);
   clk_r_REG11920_S1 : DFF_X1 port map( D => n36319, CK => CLK, Q => n41619, QN
                           => n_2714);
   clk_r_REG11918_S1 : DFF_X1 port map( D => n36320, CK => CLK, Q => n41618, QN
                           => n_2715);
   clk_r_REG11308_S1 : DFF_X1 port map( D => n36054, CK => CLK, Q => n41617, QN
                           => n_2716);
   clk_r_REG10826_S1 : DFF_X1 port map( D => n36516, CK => CLK, Q => n41616, QN
                           => n_2717);
   clk_r_REG11916_S1 : DFF_X1 port map( D => n36322, CK => CLK, Q => n41615, QN
                           => n_2718);
   clk_r_REG11631_S1 : DFF_X1 port map( D => n36323, CK => CLK, Q => n41614, QN
                           => n_2719);
   clk_r_REG11587_S1 : DFF_X1 port map( D => n36324, CK => CLK, Q => n41613, QN
                           => n_2720);
   clk_r_REG11751_S1 : DFF_X1 port map( D => n36053, CK => CLK, Q => n41612, QN
                           => n_2721);
   clk_r_REG11607_S1 : DFF_X1 port map( D => n36050, CK => CLK, Q => n41611, QN
                           => n_2722);
   clk_r_REG11609_S1 : DFF_X1 port map( D => n36049, CK => CLK, Q => n41610, QN
                           => n_2723);
   clk_r_REG11731_S1 : DFF_X1 port map( D => n36325, CK => CLK, Q => n41609, QN
                           => n_2724);
   clk_r_REG11611_S1 : DFF_X1 port map( D => n36048, CK => CLK, Q => n41608, QN
                           => n_2725);
   clk_r_REG11892_S1 : DFF_X1 port map( D => n36043, CK => CLK, Q => n41607, QN
                           => n_2726);
   clk_r_REG11310_S1 : DFF_X1 port map( D => n36042, CK => CLK, Q => n41606, QN
                           => n_2727);
   clk_r_REG11894_S1 : DFF_X1 port map( D => n36041, CK => CLK, Q => n41605, QN
                           => n_2728);
   clk_r_REG11896_S1 : DFF_X1 port map( D => n36038, CK => CLK, Q => n41604, QN
                           => n_2729);
   clk_r_REG11876_S1 : DFF_X1 port map( D => n36326, CK => CLK, Q => n41603, QN
                           => n_2730);
   clk_r_REG11312_S1 : DFF_X1 port map( D => n36037, CK => CLK, Q => n41602, QN
                           => n_2731);
   clk_r_REG11306_S1 : DFF_X1 port map( D => n36079, CK => CLK, Q => n41601, QN
                           => n_2732);
   clk_r_REG11314_S1 : DFF_X1 port map( D => n35954, CK => CLK, Q => n41600, QN
                           => n_2733);
   clk_r_REG11898_S1 : DFF_X1 port map( D => n35953, CK => CLK, Q => n41599, QN
                           => n_2734);
   clk_r_REG10793_S1 : DFF_X1 port map( D => n36328, CK => CLK, Q => n41598, QN
                           => n_2735);
   clk_r_REG12685_S1 : DFF_X1 port map( D => n35952, CK => CLK, Q => n41597, QN
                           => n_2736);
   clk_r_REG11613_S1 : DFF_X1 port map( D => n35951, CK => CLK, Q => n41596, QN
                           => n_2737);
   clk_r_REG11729_S1 : DFF_X1 port map( D => n36329, CK => CLK, Q => n41595, QN
                           => n_2738);
   clk_r_REG11874_S1 : DFF_X1 port map( D => n36330, CK => CLK, Q => n41594, QN
                           => n_2739);
   clk_r_REG11533_S1 : DFF_X1 port map( D => n35949, CK => CLK, Q => n41593, QN
                           => n_2740);
   clk_r_REG11509_S1 : DFF_X1 port map( D => n36332, CK => CLK, Q => n41592, QN
                           => n_2741);
   clk_r_REG11498_S1 : DFF_X1 port map( D => n35948, CK => CLK, Q => n41591, QN
                           => n_2742);
   clk_r_REG11290_S1 : DFF_X1 port map( D => n36333, CK => CLK, Q => n41590, QN
                           => n_2743);
   clk_r_REG11757_S1 : DFF_X1 port map( D => n35946, CK => CLK, Q => n41589, QN
                           => n_2744);
   clk_r_REG11446_S1 : DFF_X1 port map( D => n36334, CK => CLK, Q => n41588, QN
                           => n_2745);
   clk_r_REG12643_S1 : DFF_X1 port map( D => n36336, CK => CLK, Q => n41587, QN
                           => n_2746);
   clk_r_REG11900_S1 : DFF_X1 port map( D => n35945, CK => CLK, Q => n41586, QN
                           => n_2747);
   clk_r_REG11316_S1 : DFF_X1 port map( D => n35944, CK => CLK, Q => n41585, QN
                           => n_2748);
   clk_r_REG13108_S1 : DFF_X1 port map( D => n35943, CK => CLK, Q => n41584, QN
                           => n_2749);
   clk_r_REG12253_S1 : DFF_X1 port map( D => n35942, CK => CLK, Q => n41583, QN
                           => n_2750);
   clk_r_REG12687_S1 : DFF_X1 port map( D => n35941, CK => CLK, Q => n41582, QN
                           => n_2751);
   clk_r_REG11535_S1 : DFF_X1 port map( D => n35940, CK => CLK, Q => n41581, QN
                           => n_2752);
   clk_r_REG12036_S1 : DFF_X1 port map( D => n35939, CK => CLK, Q => n41580, QN
                           => n_2753);
   clk_r_REG11759_S1 : DFF_X1 port map( D => n35938, CK => CLK, Q => n41579, QN
                           => n_2754);
   clk_r_REG11500_S1 : DFF_X1 port map( D => n35937, CK => CLK, Q => n41578, QN
                           => n_2755);
   clk_r_REG11615_S1 : DFF_X1 port map( D => n35936, CK => CLK, Q => n41577, QN
                           => n_2756);
   clk_r_REG13234_S1 : DFF_X1 port map( D => n36337, CK => CLK, Q => n41576, QN
                           => n_2757);
   clk_r_REG13216_S1 : DFF_X1 port map( D => n36502, CK => CLK, Q => n41575, QN
                           => n_2758);
   clk_r_REG13224_S1 : DFF_X1 port map( D => n36498, CK => CLK, Q => n41574, QN
                           => n_2759);
   clk_r_REG13226_S1 : DFF_X1 port map( D => n36497, CK => CLK, Q => n41573, QN
                           => n_2760);
   clk_r_REG13228_S1 : DFF_X1 port map( D => n36496, CK => CLK, Q => n41572, QN
                           => n_2761);
   clk_r_REG13220_S1 : DFF_X1 port map( D => n36500, CK => CLK, Q => n41571, QN
                           => n_2762);
   clk_r_REG13230_S1 : DFF_X1 port map( D => n36495, CK => CLK, Q => n41570, QN
                           => n_2763);
   clk_r_REG13232_S1 : DFF_X1 port map( D => n36494, CK => CLK, Q => n41569, QN
                           => n_2764);
   clk_r_REG13264_S1 : DFF_X1 port map( D => n35930, CK => CLK, Q => n41568, QN
                           => n_2765);
   clk_r_REG13266_S1 : DFF_X1 port map( D => n35929, CK => CLK, Q => n41567, QN
                           => n_2766);
   clk_r_REG13268_S1 : DFF_X1 port map( D => n35927, CK => CLK, Q => n41566, QN
                           => n_2767);
   clk_r_REG11537_S1 : DFF_X1 port map( D => n35926, CK => CLK, Q => n41565, QN
                           => n_2768);
   clk_r_REG11539_S1 : DFF_X1 port map( D => n35923, CK => CLK, Q => n41564, QN
                           => n_2769);
   clk_r_REG11902_S1 : DFF_X1 port map( D => n35922, CK => CLK, Q => n41563, QN
                           => n_2770);
   clk_r_REG12691_S1 : DFF_X1 port map( D => n35921, CK => CLK, Q => n41562, QN
                           => n_2771);
   clk_r_REG12693_S1 : DFF_X1 port map( D => n35920, CK => CLK, Q => n41561, QN
                           => n_2772);
   clk_r_REG11318_S1 : DFF_X1 port map( D => n35919, CK => CLK, Q => n41560, QN
                           => n_2773);
   clk_r_REG11904_S1 : DFF_X1 port map( D => n35918, CK => CLK, Q => n41559, QN
                           => n_2774);
   clk_r_REG11320_S1 : DFF_X1 port map( D => n35917, CK => CLK, Q => n41558, QN
                           => n_2775);
   clk_r_REG13134_S1 : DFF_X1 port map( D => n35916, CK => CLK, Q => n41557, QN
                           => n_2776);
   clk_r_REG12052_S1 : DFF_X1 port map( D => n35915, CK => CLK, Q => n41556, QN
                           => n_2777);
   clk_r_REG11619_S1 : DFF_X1 port map( D => n35914, CK => CLK, Q => n41555, QN
                           => n_2778);
   clk_r_REG12054_S1 : DFF_X1 port map( D => n35913, CK => CLK, Q => n41554, QN
                           => n_2779);
   clk_r_REG11906_S1 : DFF_X1 port map( D => n35912, CK => CLK, Q => n41553, QN
                           => n_2780);
   clk_r_REG11502_S1 : DFF_X1 port map( D => n35911, CK => CLK, Q => n41552, QN
                           => n_2781);
   clk_r_REG11541_S1 : DFF_X1 port map( D => n35910, CK => CLK, Q => n41551, QN
                           => n_2782);
   clk_r_REG11506_S1 : DFF_X1 port map( D => n35907, CK => CLK, Q => n41550, QN
                           => n_2783);
   clk_r_REG11322_S1 : DFF_X1 port map( D => n35906, CK => CLK, Q => n41549, QN
                           => n_2784);
   clk_r_REG11621_S1 : DFF_X1 port map( D => n35908, CK => CLK, Q => n41548, QN
                           => n_2785);
   clk_r_REG11504_S1 : DFF_X1 port map( D => n35909, CK => CLK, Q => n41547, QN
                           => n_2786);
   clk_r_REG12689_S1 : DFF_X1 port map( D => n35924, CK => CLK, Q => n41546, QN
                           => n_2787);
   clk_r_REG12237_S1 : DFF_X1 port map( D => n36539, CK => CLK, Q => n41545, QN
                           => n_2788);
   clk_r_REG11617_S1 : DFF_X1 port map( D => n35925, CK => CLK, Q => n41544, QN
                           => n_2789);
   clk_r_REG11761_S1 : DFF_X1 port map( D => n35928, CK => CLK, Q => n41543, QN
                           => n_2790);
   clk_r_REG13132_S1 : DFF_X1 port map( D => n35947, CK => CLK, Q => n41542, QN
                           => n_2791);
   clk_r_REG12251_S1 : DFF_X1 port map( D => n35950, CK => CLK, Q => n41541, QN
                           => n_2792);
   clk_r_REG12050_S1 : DFF_X1 port map( D => n35955, CK => CLK, Q => n41540, QN
                           => n_2793);
   clk_r_REG13130_S1 : DFF_X1 port map( D => n35956, CK => CLK, Q => n41539, QN
                           => n_2794);
   clk_r_REG12239_S1 : DFF_X1 port map( D => n36526, CK => CLK, Q => n41538, QN
                           => n_2795);
   clk_r_REG11755_S1 : DFF_X1 port map( D => n35957, CK => CLK, Q => n41537, QN
                           => n_2796);
   clk_r_REG11753_S1 : DFF_X1 port map( D => n35958, CK => CLK, Q => n41536, QN
                           => n_2797);
   clk_r_REG12433_S1 : DFF_X1 port map( D => n36763, CK => CLK, Q => n41535, QN
                           => n_2798);
   clk_r_REG12555_S1 : DFF_X1 port map( D => n36527, CK => CLK, Q => n41534, QN
                           => n_2799);
   clk_r_REG12573_S1 : DFF_X1 port map( D => n36528, CK => CLK, Q => n41533, QN
                           => n_2800);
   clk_r_REG12559_S1 : DFF_X1 port map( D => n36877, CK => CLK, Q => n41532, QN
                           => n_2801);
   clk_r_REG12571_S1 : DFF_X1 port map( D => n36529, CK => CLK, Q => n41531, QN
                           => n_2802);
   clk_r_REG12241_S1 : DFF_X1 port map( D => n36364, CK => CLK, Q => n41530, QN
                           => n_2803);
   clk_r_REG12567_S1 : DFF_X1 port map( D => n36761, CK => CLK, Q => n41529, QN
                           => n_2804);
   clk_r_REG12557_S1 : DFF_X1 port map( D => n36897, CK => CLK, Q => n41528, QN
                           => n_2805);
   clk_r_REG12435_S1 : DFF_X1 port map( D => n36758, CK => CLK, Q => n41527, QN
                           => n_2806);
   clk_r_REG12569_S1 : DFF_X1 port map( D => n36755, CK => CLK, Q => n41526, QN
                           => n_2807);
   clk_r_REG12437_S1 : DFF_X1 port map( D => n36753, CK => CLK, Q => n41525, QN
                           => n_2808);
   clk_r_REG12425_S1 : DFF_X1 port map( D => n36895, CK => CLK, Q => n41524, QN
                           => n_2809);
   clk_r_REG12946_S1 : DFF_X1 port map( D => n36769, CK => CLK, Q => n41523, QN
                           => n_2810);
   clk_r_REG12443_S1 : DFF_X1 port map( D => n36530, CK => CLK, Q => n41522, QN
                           => n_2811);
   clk_r_REG12441_S1 : DFF_X1 port map( D => n36532, CK => CLK, Q => n41521, QN
                           => n_2812);
   clk_r_REG12439_S1 : DFF_X1 port map( D => n36735, CK => CLK, Q => n41520, QN
                           => n_2813);
   clk_r_REG12365_S1 : DFF_X1 port map( D => n36879, CK => CLK, Q => n41519, QN
                           => n_2814);
   clk_r_REG12379_S1 : DFF_X1 port map( D => n36518, CK => CLK, Q => n41518, QN
                           => n_2815);
   clk_r_REG12381_S1 : DFF_X1 port map( D => n36517, CK => CLK, Q => n41517, QN
                           => n_2816);
   clk_r_REG12383_S1 : DFF_X1 port map( D => n36513, CK => CLK, Q => n41516, QN
                           => n_2817);
   clk_r_REG12445_S1 : DFF_X1 port map( D => n36512, CK => CLK, Q => n41515, QN
                           => n_2818);
   clk_r_REG12387_S1 : DFF_X1 port map( D => n36861, CK => CLK, Q => n41514, QN
                           => n_2819);
   clk_r_REG12954_S1 : DFF_X1 port map( D => n36510, CK => CLK, Q => n41513, QN
                           => n_2820);
   clk_r_REG12373_S1 : DFF_X1 port map( D => n36722, CK => CLK, Q => n41512, QN
                           => n_2821);
   clk_r_REG12375_S1 : DFF_X1 port map( D => n36721, CK => CLK, Q => n41511, QN
                           => n_2822);
   clk_r_REG12575_S1 : DFF_X1 port map( D => n36509, CK => CLK, Q => n41510, QN
                           => n_2823);
   clk_r_REG12447_S1 : DFF_X1 port map( D => n36507, CK => CLK, Q => n41509, QN
                           => n_2824);
   clk_r_REG12956_S1 : DFF_X1 port map( D => n36506, CK => CLK, Q => n41508, QN
                           => n_2825);
   clk_r_REG12736_S1 : DFF_X1 port map( D => n36257, CK => CLK, Q => n41507, QN
                           => n_2826);
   clk_r_REG12371_S1 : DFF_X1 port map( D => n36724, CK => CLK, Q => n41506, QN
                           => n_2827);
   clk_r_REG12367_S1 : DFF_X1 port map( D => n36869, CK => CLK, Q => n41505, QN
                           => n_2828);
   clk_r_REG12363_S1 : DFF_X1 port map( D => n36520, CK => CLK, Q => n41504, QN
                           => n_2829);
   clk_r_REG12948_S1 : DFF_X1 port map( D => n36733, CK => CLK, Q => n41503, QN
                           => n_2830);
   clk_r_REG12337_S1 : DFF_X1 port map( D => n36786, CK => CLK, Q => n41502, QN
                           => n_2831);
   clk_r_REG13252_S1 : DFF_X1 port map( D => n36055, CK => CLK, Q => n41501, QN
                           => n_2832);
   clk_r_REG12950_S1 : DFF_X1 port map( D => n36667, CK => CLK, Q => n41500, QN
                           => n_2833);
   clk_r_REG12938_S1 : DFF_X1 port map( D => n36867, CK => CLK, Q => n41499, QN
                           => n_2834);
   clk_r_REG12942_S1 : DFF_X1 port map( D => n36793, CK => CLK, Q => n41498, QN
                           => n_2835);
   clk_r_REG12944_S1 : DFF_X1 port map( D => n36790, CK => CLK, Q => n41497, QN
                           => n_2836);
   clk_r_REG12896_S1 : DFF_X1 port map( D => n36865, CK => CLK, Q => n41496, QN
                           => n_2837);
   clk_r_REG12740_S1 : DFF_X1 port map( D => n36217, CK => CLK, Q => n41495, QN
                           => n_2838);
   clk_r_REG12726_S1 : DFF_X1 port map( D => n36752, CK => CLK, Q => n41494, QN
                           => n_2839);
   clk_r_REG12922_S1 : DFF_X1 port map( D => n36669, CK => CLK, Q => n41493, QN
                           => n_2840);
   clk_r_REG13250_S1 : DFF_X1 port map( D => n36059, CK => CLK, Q => n41492, QN
                           => n_2841);
   clk_r_REG12247_S1 : DFF_X1 port map( D => n36052, CK => CLK, Q => n41491, QN
                           => n_2842);
   clk_r_REG12728_S1 : DFF_X1 port map( D => n36750, CK => CLK, Q => n41490, QN
                           => n_2843);
   clk_r_REG12529_S1 : DFF_X1 port map( D => n36743, CK => CLK, Q => n41489, QN
                           => n_2844);
   clk_r_REG12814_S1 : DFF_X1 port map( D => n36032, CK => CLK, Q => n41488, QN
                           => n_2845);
   clk_r_REG13254_S1 : DFF_X1 port map( D => n36036, CK => CLK, Q => n41487, QN
                           => n_2846);
   clk_r_REG12806_S1 : DFF_X1 port map( D => n36288, CK => CLK, Q => n41486, QN
                           => n_2847);
   clk_r_REG12808_S1 : DFF_X1 port map( D => n36199, CK => CLK, Q => n41485, QN
                           => n_2848);
   clk_r_REG12810_S1 : DFF_X1 port map( D => n36154, CK => CLK, Q => n41484, QN
                           => n_2849);
   clk_r_REG12800_S1 : DFF_X1 port map( D => n36734, CK => CLK, Q => n41483, QN
                           => n_2850);
   clk_r_REG12812_S1 : DFF_X1 port map( D => n36149, CK => CLK, Q => n41482, QN
                           => n_2851);
   clk_r_REG12734_S1 : DFF_X1 port map( D => n36292, CK => CLK, Q => n41481, QN
                           => n_2852);
   clk_r_REG12802_S1 : DFF_X1 port map( D => n36728, CK => CLK, Q => n41480, QN
                           => n_2853);
   clk_r_REG12531_S1 : DFF_X1 port map( D => n36725, CK => CLK, Q => n41479, QN
                           => n_2854);
   clk_r_REG12804_S1 : DFF_X1 port map( D => n36293, CK => CLK, Q => n41478, QN
                           => n_2855);
   clk_r_REG12742_S1 : DFF_X1 port map( D => n36145, CK => CLK, Q => n41477, QN
                           => n_2856);
   clk_r_REG12732_S1 : DFF_X1 port map( D => n36295, CK => CLK, Q => n41476, QN
                           => n_2857);
   clk_r_REG12790_S1 : DFF_X1 port map( D => n36019, CK => CLK, Q => n41475, QN
                           => n_2858);
   clk_r_REG12744_S1 : DFF_X1 port map( D => n36018, CK => CLK, Q => n41474, QN
                           => n_2859);
   clk_r_REG12784_S1 : DFF_X1 port map( D => n36146, CK => CLK, Q => n41473, QN
                           => n_2860);
   clk_r_REG12746_S1 : DFF_X1 port map( D => n36016, CK => CLK, Q => n41472, QN
                           => n_2861);
   clk_r_REG10405_S1 : DFF_X1 port map( D => n36731, CK => CLK, Q => n41471, QN
                           => n_2862);
   clk_r_REG12245_S1 : DFF_X1 port map( D => n36147, CK => CLK, Q => n41470, QN
                           => n_2863);
   clk_r_REG11468_S1 : DFF_X1 port map( D => n36148, CK => CLK, Q => n41469, QN
                           => n_2864);
   clk_r_REG12243_S1 : DFF_X1 port map( D => n36150, CK => CLK, Q => n41468, QN
                           => n_2865);
   clk_r_REG12221_S1 : DFF_X1 port map( D => n36151, CK => CLK, Q => n41467, QN
                           => n_2866);
   clk_r_REG11466_S1 : DFF_X1 port map( D => n36152, CK => CLK, Q => n41466, QN
                           => n_2867);
   clk_r_REG11464_S1 : DFF_X1 port map( D => n36153, CK => CLK, Q => n41465, QN
                           => n_2868);
   clk_r_REG12207_S1 : DFF_X1 port map( D => n36309, CK => CLK, Q => n41464, QN
                           => n_2869);
   clk_r_REG11448_S1 : DFF_X1 port map( D => n36310, CK => CLK, Q => n41463, QN
                           => n_2870);
   clk_r_REG12219_S1 : DFF_X1 port map( D => n36155, CK => CLK, Q => n41462, QN
                           => n_2871);
   clk_r_REG12217_S1 : DFF_X1 port map( D => n36156, CK => CLK, Q => n41461, QN
                           => n_2872);
   clk_r_REG12227_S1 : DFF_X1 port map( D => n36004, CK => CLK, Q => n41460, QN
                           => n_2873);
   clk_r_REG12215_S1 : DFF_X1 port map( D => n36157, CK => CLK, Q => n41459, QN
                           => n_2874);
   clk_r_REG11462_S1 : DFF_X1 port map( D => n36160, CK => CLK, Q => n41458, QN
                           => n_2875);
   clk_r_REG11460_S1 : DFF_X1 port map( D => n36162, CK => CLK, Q => n41457, QN
                           => n_2876);
   clk_r_REG11488_S1 : DFF_X1 port map( D => n36000, CK => CLK, Q => n41456, QN
                           => n_2877);
   clk_r_REG11458_S1 : DFF_X1 port map( D => n36173, CK => CLK, Q => n41455, QN
                           => n_2878);
   clk_r_REG13256_S1 : DFF_X1 port map( D => n35998, CK => CLK, Q => n41454, QN
                           => n_2879);
   clk_r_REG11691_S1 : DFF_X1 port map( D => n36175, CK => CLK, Q => n41453, QN
                           => n_2880);
   clk_r_REG11703_S1 : DFF_X1 port map( D => n36178, CK => CLK, Q => n41452, QN
                           => n_2881);
   clk_r_REG11707_S1 : DFF_X1 port map( D => n35996, CK => CLK, Q => n41451, QN
                           => n_2882);
   clk_r_REG11701_S1 : DFF_X1 port map( D => n36180, CK => CLK, Q => n41450, QN
                           => n_2883);
   clk_r_REG11699_S1 : DFF_X1 port map( D => n36182, CK => CLK, Q => n41449, QN
                           => n_2884);
   clk_r_REG11709_S1 : DFF_X1 port map( D => n35994, CK => CLK, Q => n41448, QN
                           => n_2885);
   clk_r_REG11711_S1 : DFF_X1 port map( D => n35993, CK => CLK, Q => n41447, QN
                           => n_2886);
   clk_r_REG11697_S1 : DFF_X1 port map( D => n36185, CK => CLK, Q => n41446, QN
                           => n_2887);
   clk_r_REG11689_S1 : DFF_X1 port map( D => n36188, CK => CLK, Q => n41445, QN
                           => n_2888);
   clk_r_REG11669_S1 : DFF_X1 port map( D => n36571, CK => CLK, Q => n41444, QN
                           => n_2889);
   clk_r_REG11687_S1 : DFF_X1 port map( D => n36331, CK => CLK, Q => n41443, QN
                           => n_2890);
   clk_r_REG13258_S1 : DFF_X1 port map( D => n35991, CK => CLK, Q => n41442, QN
                           => n_2891);
   clk_r_REG13260_S1 : DFF_X1 port map( D => n35990, CK => CLK, Q => n41441, QN
                           => n_2892);
   clk_r_REG13262_S1 : DFF_X1 port map( D => n35989, CK => CLK, Q => n41440, QN
                           => n_2893);
   clk_r_REG12180_S1 : DFF_X1 port map( D => n36335, CK => CLK, Q => n41439, QN
                           => n_2894);
   clk_r_REG13178_S1 : DFF_X1 port map( D => n35987, CK => CLK, Q => n41438, QN
                           => n_2895);
   clk_r_REG13180_S1 : DFF_X1 port map( D => n35986, CK => CLK, Q => n41437, QN
                           => n_2896);
   clk_r_REG11951_S1 : DFF_X1 port map( D => n36338, CK => CLK, Q => n41436, QN
                           => n_2897);
   clk_r_REG12078_S1 : DFF_X1 port map( D => n36339, CK => CLK, Q => n41435, QN
                           => n_2898);
   clk_r_REG13200_S1 : DFF_X1 port map( D => n36340, CK => CLK, Q => n41434, QN
                           => n_2899);
   clk_r_REG12044_S1 : DFF_X1 port map( D => n36341, CK => CLK, Q => n41433, QN
                           => n_2900);
   clk_r_REG12269_S1 : DFF_X1 port map( D => n36342, CK => CLK, Q => n41432, QN
                           => n_2901);
   clk_r_REG13329_S1 : DFF_X1 port map( D => n36343, CK => CLK, Q => n41431, QN
                           => n_2902);
   clk_r_REG12205_S1 : DFF_X1 port map( D => n36344, CK => CLK, Q => n41430, QN
                           => n_2903);
   clk_r_REG12854_S1 : DFF_X1 port map( D => n36345, CK => CLK, Q => n41429, QN
                           => n_2904);
   clk_r_REG12778_S1 : DFF_X1 port map( D => n36346, CK => CLK, Q => n41428, QN
                           => n_2905);
   clk_r_REG12722_S1 : DFF_X1 port map( D => n36347, CK => CLK, Q => n41427, QN
                           => n_2906);
   clk_r_REG12583_S1 : DFF_X1 port map( D => n36834, CK => CLK, Q => n41426, QN
                           => n_2907);
   clk_r_REG13198_S1 : DFF_X1 port map( D => n36348, CK => CLK, Q => n41425, QN
                           => n_2908);
   clk_r_REG12517_S1 : DFF_X1 port map( D => n36860, CK => CLK, Q => n41424, QN
                           => n_2909);
   clk_r_REG13196_S1 : DFF_X1 port map( D => n36349, CK => CLK, Q => n41423, QN
                           => n_2910);
   clk_r_REG13204_S1 : DFF_X1 port map( D => n35971, CK => CLK, Q => n41422, QN
                           => n_2911);
   clk_r_REG13066_S1 : DFF_X1 port map( D => n36843, CK => CLK, Q => n41421, QN
                           => n_2912);
   clk_r_REG13122_S1 : DFF_X1 port map( D => n36350, CK => CLK, Q => n41420, QN
                           => n_2913);
   clk_r_REG12635_S1 : DFF_X1 port map( D => n36573, CK => CLK, Q => n41419, QN
                           => n_2914);
   clk_r_REG12625_S1 : DFF_X1 port map( D => n36847, CK => CLK, Q => n41418, QN
                           => n_2915);
   clk_r_REG13194_S1 : DFF_X1 port map( D => n36351, CK => CLK, Q => n41417, QN
                           => n_2916);
   clk_r_REG12633_S1 : DFF_X1 port map( D => n36576, CK => CLK, Q => n41416, QN
                           => n_2917);
   clk_r_REG12623_S1 : DFF_X1 port map( D => n36862, CK => CLK, Q => n41415, QN
                           => n_2918);
   clk_r_REG12631_S1 : DFF_X1 port map( D => n36578, CK => CLK, Q => n41414, QN
                           => n_2919);
   clk_r_REG13190_S1 : DFF_X1 port map( D => n36580, CK => CLK, Q => n41413, QN
                           => n_2920);
   clk_r_REG13158_S1 : DFF_X1 port map( D => n36352, CK => CLK, Q => n41412, QN
                           => n_2921);
   clk_r_REG13156_S1 : DFF_X1 port map( D => n36353, CK => CLK, Q => n41411, QN
                           => n_2922);
   clk_r_REG13182_S1 : DFF_X1 port map( D => n35961, CK => CLK, Q => n41410, QN
                           => n_2923);
   clk_r_REG13154_S1 : DFF_X1 port map( D => n36354, CK => CLK, Q => n41409, QN
                           => n_2924);
   clk_r_REG13184_S1 : DFF_X1 port map( D => n35959, CK => CLK, Q => n41408, QN
                           => n_2925);
   clk_r_REG13192_S1 : DFF_X1 port map( D => n36355, CK => CLK, Q => n41407, QN
                           => n_2926);
   clk_r_REG12621_S1 : DFF_X1 port map( D => n36868, CK => CLK, Q => n41406, QN
                           => n_2927);
   clk_r_REG12515_S1 : DFF_X1 port map( D => n36874, CK => CLK, Q => n41405, QN
                           => n_2928);
   clk_r_REG12451_S1 : DFF_X1 port map( D => n36844, CK => CLK, Q => n41404, QN
                           => n_2929);
   clk_r_REG10464_S1 : DFF_X1 port map( D => n36873, CK => CLK, Q => n41403, QN
                           => n_2930);
   clk_r_REG10471_S1 : DFF_X1 port map( D => n36888, CK => CLK, Q => n41402, QN
                           => n_2931);
   clk_r_REG12619_S1 : DFF_X1 port map( D => n36871, CK => CLK, Q => n41401, QN
                           => n_2932);
   clk_r_REG10441_S1 : DFF_X1 port map( D => n36890, CK => CLK, Q => n41400, QN
                           => n_2933);
   clk_r_REG12611_S1 : DFF_X1 port map( D => n36607, CK => CLK, Q => n41399, QN
                           => n_2934);
   clk_r_REG12581_S1 : DFF_X1 port map( D => n36853, CK => CLK, Q => n41398, QN
                           => n_2935);
   clk_r_REG12579_S1 : DFF_X1 port map( D => n36886, CK => CLK, Q => n41397, QN
                           => n_2936);
   clk_r_REG12609_S1 : DFF_X1 port map( D => n36610, CK => CLK, Q => n41396, QN
                           => n_2937);
   clk_r_REG13064_S1 : DFF_X1 port map( D => n36893, CK => CLK, Q => n41395, QN
                           => n_2938);
   clk_r_REG10378_S1 : DFF_X1 port map( D => n36881, CK => CLK, Q => n41394, QN
                           => n_2939);
   clk_r_REG10368_S1 : DFF_X1 port map( D => n36885, CK => CLK, Q => n41393, QN
                           => n_2940);
   clk_r_REG13118_S1 : DFF_X1 port map( D => n36613, CK => CLK, Q => n41392, QN
                           => n_2941);
   clk_r_REG13120_S1 : DFF_X1 port map( D => n36356, CK => CLK, Q => n41391, QN
                           => n_2942);
   clk_r_REG13116_S1 : DFF_X1 port map( D => n36619, CK => CLK, Q => n41390, QN
                           => n_2943);
   clk_r_REG13096_S1 : DFF_X1 port map( D => n36357, CK => CLK, Q => n41389, QN
                           => n_2944);
   clk_r_REG13110_S1 : DFF_X1 port map( D => n35935, CK => CLK, Q => n41388, QN
                           => n_2945);
   clk_r_REG13094_S1 : DFF_X1 port map( D => n36358, CK => CLK, Q => n41387, QN
                           => n_2946);
   clk_r_REG10920_S1 : DFF_X1 port map( D => n35934, CK => CLK, Q => n41386, QN
                           => n_2947);
   clk_r_REG11426_S1 : DFF_X1 port map( D => n35933, CK => CLK, Q => n41385, QN
                           => n_2948);
   clk_r_REG13092_S1 : DFF_X1 port map( D => n36359, CK => CLK, Q => n41384, QN
                           => n_2949);
   clk_r_REG13090_S1 : DFF_X1 port map( D => n36360, CK => CLK, Q => n41383, QN
                           => n_2950);
   clk_r_REG13112_S1 : DFF_X1 port map( D => n35932, CK => CLK, Q => n41382, QN
                           => n_2951);
   clk_r_REG13088_S1 : DFF_X1 port map( D => n36361, CK => CLK, Q => n41381, QN
                           => n_2952);
   clk_r_REG13086_S1 : DFF_X1 port map( D => n36362, CK => CLK, Q => n41380, QN
                           => n_2953);
   clk_r_REG13114_S1 : DFF_X1 port map( D => n35931, CK => CLK, Q => n41379, QN
                           => n_2954);
   clk_r_REG11835_S1 : DFF_X1 port map( D => n36363, CK => CLK, Q => n41378, QN
                           => n_2955);
   clk_r_REG13136_S1 : DFF_X1 port map( D => n35905, CK => CLK, Q => n41377, QN
                           => n_2956);
   clk_r_REG11655_S1 : DFF_X1 port map( D => n36626, CK => CLK, Q => n41376, QN
                           => n_2957);
   clk_r_REG11841_S1 : DFF_X1 port map( D => n35904, CK => CLK, Q => n41375, QN
                           => n_2958);
   clk_r_REG12184_S1 : DFF_X1 port map( D => n35903, CK => CLK, Q => n41374, QN
                           => n_2959);
   clk_r_REG12100_S1 : DFF_X1 port map( D => n35902, CK => CLK, Q => n41373, QN
                           => n_2960);
   clk_r_REG12539_S1 : DFF_X1 port map( D => n36628, CK => CLK, Q => n41372, QN
                           => n_2961);
   clk_r_REG11991_S1 : DFF_X1 port map( D => n35901, CK => CLK, Q => n41371, QN
                           => n_2962);
   clk_r_REG12056_S1 : DFF_X1 port map( D => n35900, CK => CLK, Q => n41370, QN
                           => n_2963);
   clk_r_REG12311_S1 : DFF_X1 port map( D => n35899, CK => CLK, Q => n41369, QN
                           => n_2964);
   clk_r_REG12882_S1 : DFF_X1 port map( D => n35898, CK => CLK, Q => n41368, QN
                           => n_2965);
   clk_r_REG12884_S1 : DFF_X1 port map( D => n35897, CK => CLK, Q => n41367, QN
                           => n_2966);
   clk_r_REG12878_S1 : DFF_X1 port map( D => n36365, CK => CLK, Q => n41366, QN
                           => n_2967);
   clk_r_REG12886_S1 : DFF_X1 port map( D => n35896, CK => CLK, Q => n41365, QN
                           => n_2968);
   clk_r_REG12876_S1 : DFF_X1 port map( D => n36366, CK => CLK, Q => n41364, QN
                           => n_2969);
   clk_r_REG12888_S1 : DFF_X1 port map( D => n35895, CK => CLK, Q => n41363, QN
                           => n_2970);
   clk_r_REG12874_S1 : DFF_X1 port map( D => n36367, CK => CLK, Q => n41362, QN
                           => n_2971);
   clk_r_REG13351_S1 : DFF_X1 port map( D => n35894, CK => CLK, Q => n41361, QN
                           => n_2972);
   clk_r_REG12255_S1 : DFF_X1 port map( D => n35893, CK => CLK, Q => n41360, QN
                           => n_2973);
   clk_r_REG12828_S1 : DFF_X1 port map( D => n35892, CK => CLK, Q => n41359, QN
                           => n_2974);
   clk_r_REG12764_S1 : DFF_X1 port map( D => n35891, CK => CLK, Q => n41358, QN
                           => n_2975);
   clk_r_REG12852_S1 : DFF_X1 port map( D => n36368, CK => CLK, Q => n41357, QN
                           => n_2976);
   clk_r_REG12850_S1 : DFF_X1 port map( D => n36369, CK => CLK, Q => n41356, QN
                           => n_2977);
   clk_r_REG12868_S1 : DFF_X1 port map( D => n35890, CK => CLK, Q => n41355, QN
                           => n_2978);
   clk_r_REG12848_S1 : DFF_X1 port map( D => n36370, CK => CLK, Q => n41354, QN
                           => n_2979);
   clk_r_REG12846_S1 : DFF_X1 port map( D => n36371, CK => CLK, Q => n41353, QN
                           => n_2980);
   clk_r_REG12836_S1 : DFF_X1 port map( D => n36629, CK => CLK, Q => n41352, QN
                           => n_2981);
   clk_r_REG12537_S1 : DFF_X1 port map( D => n36630, CK => CLK, Q => n41351, QN
                           => n_2982);
   clk_r_REG10450_S1 : DFF_X1 port map( D => n36876, CK => CLK, Q => n41350, QN
                           => n_2983);
   clk_r_REG12535_S1 : DFF_X1 port map( D => n36631, CK => CLK, Q => n41349, QN
                           => n_2984);
   clk_r_REG11685_S1 : DFF_X1 port map( D => n36372, CK => CLK, Q => n41348, QN
                           => n_2985);
   clk_r_REG11420_S1 : DFF_X1 port map( D => n36373, CK => CLK, Q => n41347, QN
                           => n_2986);
   clk_r_REG10934_S1 : DFF_X1 port map( D => n36374, CK => CLK, Q => n41346, QN
                           => n_2987);
   clk_r_REG11833_S1 : DFF_X1 port map( D => n36375, CK => CLK, Q => n41345, QN
                           => n_2988);
   clk_r_REG12178_S1 : DFF_X1 port map( D => n36376, CK => CLK, Q => n41344, QN
                           => n_2989);
   clk_r_REG12110_S1 : DFF_X1 port map( D => n36377, CK => CLK, Q => n41343, QN
                           => n_2990);
   clk_r_REG11983_S1 : DFF_X1 port map( D => n36378, CK => CLK, Q => n41342, QN
                           => n_2991);
   clk_r_REG12042_S1 : DFF_X1 port map( D => n36379, CK => CLK, Q => n41341, QN
                           => n_2992);
   clk_r_REG12305_S1 : DFF_X1 port map( D => n36380, CK => CLK, Q => n41340, QN
                           => n_2993);
   clk_r_REG13343_S1 : DFF_X1 port map( D => n36381, CK => CLK, Q => n41339, QN
                           => n_2994);
   clk_r_REG13014_S1 : DFF_X1 port map( D => n36640, CK => CLK, Q => n41338, QN
                           => n_2995);
   clk_r_REG12924_S1 : DFF_X1 port map( D => n36641, CK => CLK, Q => n41337, QN
                           => n_2996);
   clk_r_REG13078_S1 : DFF_X1 port map( D => n36642, CK => CLK, Q => n41336, QN
                           => n_2997);
   clk_r_REG12347_S1 : DFF_X1 port map( D => n36645, CK => CLK, Q => n41335, QN
                           => n_2998);
   clk_r_REG12411_S1 : DFF_X1 port map( D => n36647, CK => CLK, Q => n41334, QN
                           => n_2999);
   clk_r_REG12998_S1 : DFF_X1 port map( D => n36883, CK => CLK, Q => n41333, QN
                           => n_3000);
   clk_r_REG13012_S1 : DFF_X1 port map( D => n36649, CK => CLK, Q => n41332, QN
                           => n_3001);
   clk_r_REG13010_S1 : DFF_X1 port map( D => n36650, CK => CLK, Q => n41331, QN
                           => n_3002);
   clk_r_REG13008_S1 : DFF_X1 port map( D => n36651, CK => CLK, Q => n41330, QN
                           => n_3003);
   clk_r_REG13000_S1 : DFF_X1 port map( D => n36859, CK => CLK, Q => n41329, QN
                           => n_3004);
   clk_r_REG13002_S1 : DFF_X1 port map( D => n36856, CK => CLK, Q => n41328, QN
                           => n_3005);
   clk_r_REG12980_S1 : DFF_X1 port map( D => n36658, CK => CLK, Q => n41327, QN
                           => n_3006);
   clk_r_REG12958_S1 : DFF_X1 port map( D => n36854, CK => CLK, Q => n41326, QN
                           => n_3007);
   clk_r_REG12966_S1 : DFF_X1 port map( D => n36832, CK => CLK, Q => n41325, QN
                           => n_3008);
   clk_r_REG12499_S1 : DFF_X1 port map( D => n36660, CK => CLK, Q => n41324, QN
                           => n_3009);
   clk_r_REG12766_S1 : DFF_X1 port map( D => n35889, CK => CLK, Q => n41323, QN
                           => n_3010);
   clk_r_REG12960_S1 : DFF_X1 port map( D => n36849, CK => CLK, Q => n41322, QN
                           => n_3011);
   clk_r_REG12984_S1 : DFF_X1 port map( D => n36634, CK => CLK, Q => n41321, QN
                           => n_3012);
   clk_r_REG12962_S1 : DFF_X1 port map( D => n36848, CK => CLK, Q => n41320, QN
                           => n_3013);
   clk_r_REG12830_S1 : DFF_X1 port map( D => n35888, CK => CLK, Q => n41319, QN
                           => n_3014);
   clk_r_REG12257_S1 : DFF_X1 port map( D => n35887, CK => CLK, Q => n41318, QN
                           => n_3015);
   clk_r_REG13353_S1 : DFF_X1 port map( D => n35886, CK => CLK, Q => n41317, QN
                           => n_3016);
   clk_r_REG12313_S1 : DFF_X1 port map( D => n35885, CK => CLK, Q => n41316, QN
                           => n_3017);
   clk_r_REG12038_S1 : DFF_X1 port map( D => n36678, CK => CLK, Q => n41315, QN
                           => n_3018);
   clk_r_REG11993_S1 : DFF_X1 port map( D => n35884, CK => CLK, Q => n41314, QN
                           => n_3019);
   clk_r_REG12493_S1 : DFF_X1 port map( D => n36842, CK => CLK, Q => n41313, QN
                           => n_3020);
   clk_r_REG12389_S1 : DFF_X1 port map( D => n36841, CK => CLK, Q => n41312, QN
                           => n_3021);
   clk_r_REG12323_S1 : DFF_X1 port map( D => n36839, CK => CLK, Q => n41311, QN
                           => n_3022);
   clk_r_REG13068_S1 : DFF_X1 port map( D => n36837, CK => CLK, Q => n41310, QN
                           => n_3023);
   clk_r_REG12898_S1 : DFF_X1 port map( D => n36836, CK => CLK, Q => n41309, QN
                           => n_3024);
   clk_r_REG12116_S1 : DFF_X1 port map( D => n35883, CK => CLK, Q => n41308, QN
                           => n_3025);
   clk_r_REG12186_S1 : DFF_X1 port map( D => n35882, CK => CLK, Q => n41307, QN
                           => n_3026);
   clk_r_REG11843_S1 : DFF_X1 port map( D => n35881, CK => CLK, Q => n41306, QN
                           => n_3027);
   clk_r_REG10942_S1 : DFF_X1 port map( D => n35880, CK => CLK, Q => n41305, QN
                           => n_3028);
   clk_r_REG11428_S1 : DFF_X1 port map( D => n35879, CK => CLK, Q => n41304, QN
                           => n_3029);
   clk_r_REG11845_S1 : DFF_X1 port map( D => n35878, CK => CLK, Q => n41303, QN
                           => n_3030);
   clk_r_REG13074_S1 : DFF_X1 port map( D => n36802, CK => CLK, Q => n41302, QN
                           => n_3031);
   clk_r_REG13072_S1 : DFF_X1 port map( D => n36804, CK => CLK, Q => n41301, QN
                           => n_3032);
   clk_r_REG11430_S1 : DFF_X1 port map( D => n35877, CK => CLK, Q => n41300, QN
                           => n_3033);
   clk_r_REG10944_S1 : DFF_X1 port map( D => n35876, CK => CLK, Q => n41299, QN
                           => n_3034);
   clk_r_REG12188_S1 : DFF_X1 port map( D => n35875, CK => CLK, Q => n41298, QN
                           => n_3035);
   clk_r_REG12118_S1 : DFF_X1 port map( D => n35874, CK => CLK, Q => n41297, QN
                           => n_3036);
   clk_r_REG13076_S1 : DFF_X1 port map( D => n36673, CK => CLK, Q => n41296, QN
                           => n_3037);
   clk_r_REG13070_S1 : DFF_X1 port map( D => n36806, CK => CLK, Q => n41295, QN
                           => n_3038);
   clk_r_REG11995_S1 : DFF_X1 port map( D => n35873, CK => CLK, Q => n41294, QN
                           => n_3039);
   clk_r_REG13048_S1 : DFF_X1 port map( D => n36688, CK => CLK, Q => n41293, QN
                           => n_3040);
   clk_r_REG13046_S1 : DFF_X1 port map( D => n36689, CK => CLK, Q => n41292, QN
                           => n_3041);
   clk_r_REG13042_S1 : DFF_X1 port map( D => n36699, CK => CLK, Q => n41291, QN
                           => n_3042);
   clk_r_REG13024_S1 : DFF_X1 port map( D => n36808, CK => CLK, Q => n41290, QN
                           => n_3043);
   clk_r_REG13022_S1 : DFF_X1 port map( D => n36817, CK => CLK, Q => n41289, QN
                           => n_3044);
   clk_r_REG13044_S1 : DFF_X1 port map( D => n36697, CK => CLK, Q => n41288, QN
                           => n_3045);
   clk_r_REG12058_S1 : DFF_X1 port map( D => n35872, CK => CLK, Q => n41287, QN
                           => n_3046);
   clk_r_REG12297_S1 : DFF_X1 port map( D => n36693, CK => CLK, Q => n41286, QN
                           => n_3047);
   clk_r_REG10302_S1 : DFF_X1 port map( D => n36702, CK => CLK, Q => n41285, QN
                           => n_3048);
   clk_r_REG12908_S1 : DFF_X1 port map( D => n36820, CK => CLK, Q => n41284, QN
                           => n_3049);
   clk_r_REG12906_S1 : DFF_X1 port map( D => n36821, CK => CLK, Q => n41283, QN
                           => n_3050);
   clk_r_REG12327_S1 : DFF_X1 port map( D => n36823, CK => CLK, Q => n41282, QN
                           => n_3051);
   clk_r_REG12920_S1 : DFF_X1 port map( D => n36672, CK => CLK, Q => n41281, QN
                           => n_3052);
   clk_r_REG12916_S1 : DFF_X1 port map( D => n36695, CK => CLK, Q => n41280, QN
                           => n_3053);
   clk_r_REG12904_S1 : DFF_X1 port map( D => n36827, CK => CLK, Q => n41279, QN
                           => n_3054);
   clk_r_REG12902_S1 : DFF_X1 port map( D => n36828, CK => CLK, Q => n41278, QN
                           => n_3055);
   clk_r_REG12525_S1 : DFF_X1 port map( D => n36829, CK => CLK, Q => n41277, QN
                           => n_3056);
   clk_r_REG12918_S1 : DFF_X1 port map( D => n36690, CK => CLK, Q => n41276, QN
                           => n_3057);
   clk_r_REG12900_S1 : DFF_X1 port map( D => n36830, CK => CLK, Q => n41275, QN
                           => n_3058);
   clk_r_REG12507_S1 : DFF_X1 port map( D => n36632, CK => CLK, Q => n41274, QN
                           => n_3059);
   clk_r_REG12391_S1 : DFF_X1 port map( D => n36831, CK => CLK, Q => n41273, QN
                           => n_3060);
   clk_r_REG12403_S1 : DFF_X1 port map( D => n36686, CK => CLK, Q => n41272, QN
                           => n_3061);
   clk_r_REG12393_S1 : DFF_X1 port map( D => n36825, CK => CLK, Q => n41271, QN
                           => n_3062);
   clk_r_REG12395_S1 : DFF_X1 port map( D => n36824, CK => CLK, Q => n41270, QN
                           => n_3063);
   clk_r_REG12397_S1 : DFF_X1 port map( D => n36819, CK => CLK, Q => n41269, QN
                           => n_3064);
   clk_r_REG12405_S1 : DFF_X1 port map( D => n36682, CK => CLK, Q => n41268, QN
                           => n_3065);
   clk_r_REG12409_S1 : DFF_X1 port map( D => n36671, CK => CLK, Q => n41267, QN
                           => n_3066);
   clk_r_REG12399_S1 : DFF_X1 port map( D => n36818, CK => CLK, Q => n41266, QN
                           => n_3067);
   clk_r_REG12349_S1 : DFF_X1 port map( D => n36633, CK => CLK, Q => n41265, QN
                           => n_3068);
   clk_r_REG10932_S1 : DFF_X1 port map( D => n36382, CK => CLK, Q => n41264, QN
                           => n_3069);
   clk_r_REG12331_S1 : DFF_X1 port map( D => n36815, CK => CLK, Q => n41263, QN
                           => n_3070);
   clk_r_REG11418_S1 : DFF_X1 port map( D => n36383, CK => CLK, Q => n41262, QN
                           => n_3071);
   clk_r_REG12333_S1 : DFF_X1 port map( D => n36812, CK => CLK, Q => n41261, QN
                           => n_3072);
   clk_r_REG11683_S1 : DFF_X1 port map( D => n36384, CK => CLK, Q => n41260, QN
                           => n_3073);
   clk_r_REG12343_S1 : DFF_X1 port map( D => n36657, CK => CLK, Q => n41259, QN
                           => n_3074);
   clk_r_REG12345_S1 : DFF_X1 port map( D => n36656, CK => CLK, Q => n41258, QN
                           => n_3075);
   clk_r_REG11831_S1 : DFF_X1 port map( D => n36385, CK => CLK, Q => n41257, QN
                           => n_3076);
   clk_r_REG12176_S1 : DFF_X1 port map( D => n36386, CK => CLK, Q => n41256, QN
                           => n_3077);
   clk_r_REG12112_S1 : DFF_X1 port map( D => n36259, CK => CLK, Q => n41255, QN
                           => n_3078);
   clk_r_REG11985_S1 : DFF_X1 port map( D => n36260, CK => CLK, Q => n41254, QN
                           => n_3079);
   clk_r_REG12329_S1 : DFF_X1 port map( D => n36822, CK => CLK, Q => n41253, QN
                           => n_3080);
   clk_r_REG12325_S1 : DFF_X1 port map( D => n36826, CK => CLK, Q => n41252, QN
                           => n_3081);
   clk_r_REG12016_S1 : DFF_X1 port map( D => n36261, CK => CLK, Q => n41251, QN
                           => n_3082);
   clk_r_REG12307_S1 : DFF_X1 port map( D => n36262, CK => CLK, Q => n41250, QN
                           => n_3083);
   clk_r_REG12491_S1 : DFF_X1 port map( D => n36858, CK => CLK, Q => n41249, QN
                           => n_3084);
   clk_r_REG13345_S1 : DFF_X1 port map( D => n36263, CK => CLK, Q => n41248, QN
                           => n_3085);
   clk_r_REG12209_S1 : DFF_X1 port map( D => n36264, CK => CLK, Q => n41247, QN
                           => n_3086);
   clk_r_REG12780_S1 : DFF_X1 port map( D => n36265, CK => CLK, Q => n41246, QN
                           => n_3087);
   clk_r_REG12720_S1 : DFF_X1 port map( D => n36387, CK => CLK, Q => n41245, QN
                           => n_3088);
   clk_r_REG10398_S1 : DFF_X1 port map( D => n36488, CK => CLK, Q => n41244, QN
                           => n_3089);
   clk_r_REG12201_S1 : DFF_X1 port map( D => n36461, CK => CLK, Q => n41243, QN
                           => n_3090);
   clk_r_REG13339_S1 : DFF_X1 port map( D => n36459, CK => CLK, Q => n41242, QN
                           => n_3091);
   clk_r_REG12505_S1 : DFF_X1 port map( D => n36637, CK => CLK, Q => n41241, QN
                           => n_3092);
   clk_r_REG12710_S1 : DFF_X1 port map( D => n36491, CK => CLK, Q => n41240, QN
                           => n_3093);
   clk_r_REG12503_S1 : DFF_X1 port map( D => n36655, CK => CLK, Q => n41239, QN
                           => n_3094);
   clk_r_REG12501_S1 : DFF_X1 port map( D => n36659, CK => CLK, Q => n41238, QN
                           => n_3095);
   clk_r_REG12455_S1 : DFF_X1 port map( D => n36816, CK => CLK, Q => n41237, QN
                           => n_3096);
   clk_r_REG12457_S1 : DFF_X1 port map( D => n36814, CK => CLK, Q => n41236, QN
                           => n_3097);
   clk_r_REG12477_S1 : DFF_X1 port map( D => n36665, CK => CLK, Q => n41235, QN
                           => n_3098);
   clk_r_REG12459_S1 : DFF_X1 port map( D => n36810, CK => CLK, Q => n41234, QN
                           => n_3099);
   clk_r_REG12461_S1 : DFF_X1 port map( D => n36809, CK => CLK, Q => n41233, QN
                           => n_3100);
   clk_r_REG12301_S1 : DFF_X1 port map( D => n36438, CK => CLK, Q => n41232, QN
                           => n_3101);
   clk_r_REG12008_S1 : DFF_X1 port map( D => n36437, CK => CLK, Q => n41231, QN
                           => n_3102);
   clk_r_REG12453_S1 : DFF_X1 port map( D => n36840, CK => CLK, Q => n41230, QN
                           => n_3103);
   clk_r_REG11979_S1 : DFF_X1 port map( D => n36434, CK => CLK, Q => n41229, QN
                           => n_3104);
   clk_r_REG12106_S1 : DFF_X1 port map( D => n36432, CK => CLK, Q => n41228, QN
                           => n_3105);
   clk_r_REG12172_S1 : DFF_X1 port map( D => n36430, CK => CLK, Q => n41227, QN
                           => n_3106);
   clk_r_REG11827_S1 : DFF_X1 port map( D => n36428, CK => CLK, Q => n41226, QN
                           => n_3107);
   clk_r_REG11675_S1 : DFF_X1 port map( D => n36424, CK => CLK, Q => n41225, QN
                           => n_3108);
   clk_r_REG11412_S1 : DFF_X1 port map( D => n36423, CK => CLK, Q => n41224, QN
                           => n_3109);
   clk_r_REG10926_S1 : DFF_X1 port map( D => n36421, CK => CLK, Q => n41223, QN
                           => n_3110);
   clk_r_REG12523_S1 : DFF_X1 port map( D => n36845, CK => CLK, Q => n41222, QN
                           => n_3111);
   clk_r_REG12521_S1 : DFF_X1 port map( D => n36846, CK => CLK, Q => n41221, QN
                           => n_3112);
   clk_r_REG12533_S1 : DFF_X1 port map( D => n36635, CK => CLK, Q => n41220, QN
                           => n_3113);
   clk_r_REG12519_S1 : DFF_X1 port map( D => n36850, CK => CLK, Q => n41219, QN
                           => n_3114);
   clk_r_REG11414_S1 : DFF_X1 port map( D => n36415, CK => CLK, Q => n41218, QN
                           => n_3115);
   clk_r_REG11677_S1 : DFF_X1 port map( D => n36414, CK => CLK, Q => n41217, QN
                           => n_3116);
   clk_r_REG11679_S1 : DFF_X1 port map( D => n36412, CK => CLK, Q => n41216, QN
                           => n_3117);
   clk_r_REG10777_S1 : DFF_X1 port map( D => n36644, CK => CLK, Q => n41215, QN
                           => n_3118);
   clk_r_REG11681_S1 : DFF_X1 port map( D => n36405, CK => CLK, Q => n41214, QN
                           => n_3119);
   clk_r_REG11671_S1 : DFF_X1 port map( D => n36448, CK => CLK, Q => n41213, QN
                           => n_3120);
   clk_r_REG11705_S1 : DFF_X1 port map( D => n36044, CK => CLK, Q => n41212, QN
                           => n_3121);
   clk_r_REG10930_S1 : DFF_X1 port map( D => n36388, CK => CLK, Q => n41211, QN
                           => n_3122);
   clk_r_REG11416_S1 : DFF_X1 port map( D => n36389, CK => CLK, Q => n41210, QN
                           => n_3123);
   clk_r_REG11829_S1 : DFF_X1 port map( D => n36390, CK => CLK, Q => n41209, QN
                           => n_3124);
   clk_r_REG11801_S1 : DFF_X1 port map( D => n36391, CK => CLK, Q => n41208, QN
                           => n_3125);
   clk_r_REG11819_S1 : DFF_X1 port map( D => n36047, CK => CLK, Q => n41207, QN
                           => n_3126);
   clk_r_REG11799_S1 : DFF_X1 port map( D => n36392, CK => CLK, Q => n41206, QN
                           => n_3127);
   clk_r_REG11797_S1 : DFF_X1 port map( D => n36393, CK => CLK, Q => n41205, QN
                           => n_3128);
   clk_r_REG11817_S1 : DFF_X1 port map( D => n36058, CK => CLK, Q => n41204, QN
                           => n_3129);
   clk_r_REG11815_S1 : DFF_X1 port map( D => n36061, CK => CLK, Q => n41203, QN
                           => n_3130);
   clk_r_REG12174_S1 : DFF_X1 port map( D => n36394, CK => CLK, Q => n41202, QN
                           => n_3131);
   clk_r_REG12108_S1 : DFF_X1 port map( D => n36395, CK => CLK, Q => n41201, QN
                           => n_3132);
   clk_r_REG11981_S1 : DFF_X1 port map( D => n36396, CK => CLK, Q => n41200, QN
                           => n_3133);
   clk_r_REG12014_S1 : DFF_X1 port map( D => n36397, CK => CLK, Q => n41199, QN
                           => n_3134);
   clk_r_REG12303_S1 : DFF_X1 port map( D => n36400, CK => CLK, Q => n41198, QN
                           => n_3135);
   clk_r_REG13341_S1 : DFF_X1 port map( D => n36401, CK => CLK, Q => n41197, QN
                           => n_3136);
   clk_r_REG12203_S1 : DFF_X1 port map( D => n36402, CK => CLK, Q => n41196, QN
                           => n_3137);
   clk_r_REG12776_S1 : DFF_X1 port map( D => n36406, CK => CLK, Q => n41195, QN
                           => n_3138);
   clk_r_REG12148_S1 : DFF_X1 port map( D => n36407, CK => CLK, Q => n41194, QN
                           => n_3139);
   clk_r_REG12146_S1 : DFF_X1 port map( D => n36408, CK => CLK, Q => n41193, QN
                           => n_3140);
   clk_r_REG12162_S1 : DFF_X1 port map( D => n36064, CK => CLK, Q => n41192, QN
                           => n_3141);
   clk_r_REG12144_S1 : DFF_X1 port map( D => n36409, CK => CLK, Q => n41191, QN
                           => n_3142);
   clk_r_REG12160_S1 : DFF_X1 port map( D => n36066, CK => CLK, Q => n41190, QN
                           => n_3143);
   clk_r_REG12158_S1 : DFF_X1 port map( D => n36071, CK => CLK, Q => n41189, QN
                           => n_3144);
   clk_r_REG12718_S1 : DFF_X1 port map( D => n36410, CK => CLK, Q => n41188, QN
                           => n_3145);
   clk_r_REG12076_S1 : DFF_X1 port map( D => n36411, CK => CLK, Q => n41187, QN
                           => n_3146);
   clk_r_REG12074_S1 : DFF_X1 port map( D => n36413, CK => CLK, Q => n41186, QN
                           => n_3147);
   clk_r_REG12096_S1 : DFF_X1 port map( D => n36068, CK => CLK, Q => n41185, QN
                           => n_3148);
   clk_r_REG12072_S1 : DFF_X1 port map( D => n36416, CK => CLK, Q => n41184, QN
                           => n_3149);
   clk_r_REG12094_S1 : DFF_X1 port map( D => n36080, CK => CLK, Q => n41183, QN
                           => n_3150);
   clk_r_REG12114_S1 : DFF_X1 port map( D => n36076, CK => CLK, Q => n41182, QN
                           => n_3151);
   clk_r_REG10928_S1 : DFF_X1 port map( D => n36417, CK => CLK, Q => n41181, QN
                           => n_3152);
   clk_r_REG11392_S1 : DFF_X1 port map( D => n36418, CK => CLK, Q => n41180, QN
                           => n_3153);
   clk_r_REG11949_S1 : DFF_X1 port map( D => n36419, CK => CLK, Q => n41179, QN
                           => n_3154);
   clk_r_REG12012_S1 : DFF_X1 port map( D => n36435, CK => CLK, Q => n41178, QN
                           => n_3155);
   clk_r_REG12010_S1 : DFF_X1 port map( D => n36436, CK => CLK, Q => n41177, QN
                           => n_3156);
   clk_r_REG12006_S1 : DFF_X1 port map( D => n36439, CK => CLK, Q => n41176, QN
                           => n_3157);
   clk_r_REG12030_S1 : DFF_X1 port map( D => n36045, CK => CLK, Q => n41175, QN
                           => n_3158);
   clk_r_REG12032_S1 : DFF_X1 port map( D => n36035, CK => CLK, Q => n41174, QN
                           => n_3159);
   clk_r_REG12034_S1 : DFF_X1 port map( D => n36031, CK => CLK, Q => n41173, QN
                           => n_3160);
   clk_r_REG11673_S1 : DFF_X1 port map( D => n36440, CK => CLK, Q => n41172, QN
                           => n_3161);
   clk_r_REG10840_S1 : DFF_X1 port map( D => n36675, CK => CLK, Q => n41171, QN
                           => n_3162);
   clk_r_REG11406_S1 : DFF_X1 port map( D => n36030, CK => CLK, Q => n41170, QN
                           => n_3163);
   clk_r_REG11388_S1 : DFF_X1 port map( D => n36444, CK => CLK, Q => n41169, QN
                           => n_3164);
   clk_r_REG11386_S1 : DFF_X1 port map( D => n36445, CK => CLK, Q => n41168, QN
                           => n_3165);
   clk_r_REG11378_S1 : DFF_X1 port map( D => n36668, CK => CLK, Q => n41167, QN
                           => n_3166);
   clk_r_REG12706_S1 : DFF_X1 port map( D => n36691, CK => CLK, Q => n41166, QN
                           => n_3167);
   clk_r_REG12786_S1 : DFF_X1 port map( D => n36029, CK => CLK, Q => n41165, QN
                           => n_3168);
   clk_r_REG12223_S1 : DFF_X1 port map( D => n36028, CK => CLK, Q => n41164, QN
                           => n_3169);
   clk_r_REG13311_S1 : DFF_X1 port map( D => n36670, CK => CLK, Q => n41163, QN
                           => n_3170);
   clk_r_REG12285_S1 : DFF_X1 port map( D => n36027, CK => CLK, Q => n41162, QN
                           => n_3171);
   clk_r_REG10908_S1 : DFF_X1 port map( D => n36026, CK => CLK, Q => n41161, QN
                           => n_3172);
   clk_r_REG10896_S1 : DFF_X1 port map( D => n36446, CK => CLK, Q => n41160, QN
                           => n_3173);
   clk_r_REG10894_S1 : DFF_X1 port map( D => n36447, CK => CLK, Q => n41159, QN
                           => n_3174);
   clk_r_REG11961_S1 : DFF_X1 port map( D => n36025, CK => CLK, Q => n41158, QN
                           => n_3175);
   clk_r_REG10879_S1 : DFF_X1 port map( D => n36458, CK => CLK, Q => n41157, QN
                           => n_3176);
   clk_r_REG10910_S1 : DFF_X1 port map( D => n36024, CK => CLK, Q => n41156, QN
                           => n_3177);
   clk_r_REG10912_S1 : DFF_X1 port map( D => n36022, CK => CLK, Q => n41155, QN
                           => n_3178);
   clk_r_REG12716_S1 : DFF_X1 port map( D => n36452, CK => CLK, Q => n41154, QN
                           => n_3179);
   clk_r_REG12774_S1 : DFF_X1 port map( D => n36453, CK => CLK, Q => n41153, QN
                           => n_3180);
   clk_r_REG12197_S1 : DFF_X1 port map( D => n36463, CK => CLK, Q => n41152, QN
                           => n_3181);
   clk_r_REG13327_S1 : DFF_X1 port map( D => n36464, CK => CLK, Q => n41151, QN
                           => n_3182);
   clk_r_REG12267_S1 : DFF_X1 port map( D => n36460, CK => CLK, Q => n41150, QN
                           => n_3183);
   clk_r_REG11945_S1 : DFF_X1 port map( D => n36467, CK => CLK, Q => n41149, QN
                           => n_3184);
   clk_r_REG12599_S1 : DFF_X1 port map( D => n36680, CK => CLK, Q => n41148, QN
                           => n_3185);
   clk_r_REG12714_S1 : DFF_X1 port map( D => n36468, CK => CLK, Q => n41147, QN
                           => n_3186);
   clk_r_REG12772_S1 : DFF_X1 port map( D => n36471, CK => CLK, Q => n41146, QN
                           => n_3187);
   clk_r_REG10489_S1 : DFF_X1 port map( D => n36473, CK => CLK, Q => n41145, QN
                           => n_3188);
   clk_r_REG13325_S1 : DFF_X1 port map( D => n36466, CK => CLK, Q => n41144, QN
                           => n_3189);
   clk_r_REG12263_S1 : DFF_X1 port map( D => n36482, CK => CLK, Q => n41143, QN
                           => n_3190);
   clk_r_REG11943_S1 : DFF_X1 port map( D => n36476, CK => CLK, Q => n41142, QN
                           => n_3191);
   clk_r_REG12265_S1 : DFF_X1 port map( D => n36479, CK => CLK, Q => n41141, QN
                           => n_3192);
   clk_r_REG10482_S1 : DFF_X1 port map( D => n36663, CK => CLK, Q => n41140, QN
                           => n_3193);
   clk_r_REG12287_S1 : DFF_X1 port map( D => n36021, CK => CLK, Q => n41139, QN
                           => n_3194);
   clk_r_REG12770_S1 : DFF_X1 port map( D => n36475, CK => CLK, Q => n41138, QN
                           => n_3195);
   clk_r_REG12788_S1 : DFF_X1 port map( D => n36020, CK => CLK, Q => n41137, QN
                           => n_3196);
   clk_r_REG12792_S1 : DFF_X1 port map( D => n36017, CK => CLK, Q => n41136, QN
                           => n_3197);
   clk_r_REG12748_S1 : DFF_X1 port map( D => n36015, CK => CLK, Q => n41135, QN
                           => n_3198);
   clk_r_REG12750_S1 : DFF_X1 port map( D => n36014, CK => CLK, Q => n41134, QN
                           => n_3199);
   clk_r_REG12712_S1 : DFF_X1 port map( D => n36481, CK => CLK, Q => n41133, QN
                           => n_3200);
   clk_r_REG12225_S1 : DFF_X1 port map( D => n36013, CK => CLK, Q => n41132, QN
                           => n_3201);
   clk_r_REG13313_S1 : DFF_X1 port map( D => n36653, CK => CLK, Q => n41131, QN
                           => n_3202);
   clk_r_REG13315_S1 : DFF_X1 port map( D => n36646, CK => CLK, Q => n41130, QN
                           => n_3203);
   clk_r_REG13321_S1 : DFF_X1 port map( D => n36492, CK => CLK, Q => n41129, QN
                           => n_3204);
   clk_r_REG11963_S1 : DFF_X1 port map( D => n36012, CK => CLK, Q => n41128, QN
                           => n_3205);
   clk_r_REG12249_S1 : DFF_X1 port map( D => n36011, CK => CLK, Q => n41127, QN
                           => n_3206);
   clk_r_REG12199_S1 : DFF_X1 port map( D => n36462, CK => CLK, Q => n41126, QN
                           => n_3207);
   clk_r_REG11965_S1 : DFF_X1 port map( D => n36010, CK => CLK, Q => n41125, QN
                           => n_3208);
   clk_r_REG11967_S1 : DFF_X1 port map( D => n36009, CK => CLK, Q => n41124, QN
                           => n_3209);
   clk_r_REG12982_S1 : DFF_X1 port map( D => n36639, CK => CLK, Q => n41123, QN
                           => n_3210);
   clk_r_REG11408_S1 : DFF_X1 port map( D => n36008, CK => CLK, Q => n41122, QN
                           => n_3211);
   clk_r_REG12752_S1 : DFF_X1 port map( D => n36007, CK => CLK, Q => n41121, QN
                           => n_3212);
   clk_r_REG10914_S1 : DFF_X1 port map( D => n36006, CK => CLK, Q => n41120, QN
                           => n_3213);
   clk_r_REG12351_S1 : DFF_X1 port map( D => n36604, CK => CLK, Q => n41119, QN
                           => n_3214);
   clk_r_REG12289_S1 : DFF_X1 port map( D => n36005, CK => CLK, Q => n41118, QN
                           => n_3215);
   clk_r_REG12098_S1 : DFF_X1 port map( D => n36003, CK => CLK, Q => n41117, QN
                           => n_3216);
   clk_r_REG13176_S1 : DFF_X1 port map( D => n36002, CK => CLK, Q => n41116, QN
                           => n_3217);
   clk_r_REG12483_S1 : DFF_X1 port map( D => n36603, CK => CLK, Q => n41115, QN
                           => n_3218);
   clk_r_REG12613_S1 : DFF_X1 port map( D => n36601, CK => CLK, Q => n41114, QN
                           => n_3219);
   clk_r_REG12794_S1 : DFF_X1 port map( D => n36001, CK => CLK, Q => n41113, QN
                           => n_3220);
   clk_r_REG11663_S1 : DFF_X1 port map( D => n36600, CK => CLK, Q => n41112, QN
                           => n_3221);
   clk_r_REG12838_S1 : DFF_X1 port map( D => n36599, CK => CLK, Q => n41111, QN
                           => n_3222);
   clk_r_REG11821_S1 : DFF_X1 port map( D => n35999, CK => CLK, Q => n41110, QN
                           => n_3223);
   clk_r_REG12164_S1 : DFF_X1 port map( D => n35997, CK => CLK, Q => n41109, QN
                           => n_3224);
   clk_r_REG12541_S1 : DFF_X1 port map( D => n36596, CK => CLK, Q => n41108, QN
                           => n_3225);
   clk_r_REG13058_S1 : DFF_X1 port map( D => n36595, CK => CLK, Q => n41107, QN
                           => n_3226);
   clk_r_REG13317_S1 : DFF_X1 port map( D => n36590, CK => CLK, Q => n41106, QN
                           => n_3227);
   clk_r_REG12413_S1 : DFF_X1 port map( D => n36588, CK => CLK, Q => n41105, QN
                           => n_3228);
   clk_r_REG12926_S1 : DFF_X1 port map( D => n36587, CK => CLK, Q => n41104, QN
                           => n_3229);
   clk_r_REG12910_S1 : DFF_X1 port map( D => n36787, CK => CLK, Q => n41103, QN
                           => n_3230);
   clk_r_REG12565_S1 : DFF_X1 port map( D => n36764, CK => CLK, Q => n41102, QN
                           => n_3231);
   clk_r_REG12235_S1 : DFF_X1 port map( D => n36585, CK => CLK, Q => n41101, QN
                           => n_3232);
   clk_r_REG12211_S1 : DFF_X1 port map( D => n36237, CK => CLK, Q => n41100, QN
                           => n_3233);
   clk_r_REG12213_S1 : DFF_X1 port map( D => n36236, CK => CLK, Q => n41099, QN
                           => n_3234);
   clk_r_REG12914_S1 : DFF_X1 port map( D => n36770, CK => CLK, Q => n41098, QN
                           => n_3235);
   clk_r_REG12543_S1 : DFF_X1 port map( D => n36581, CK => CLK, Q => n41097, QN
                           => n_3236);
   clk_r_REG12423_S1 : DFF_X1 port map( D => n36542, CK => CLK, Q => n41096, QN
                           => n_3237);
   clk_r_REG12754_S1 : DFF_X1 port map( D => n35995, CK => CLK, Q => n41095, QN
                           => n_3238);
   clk_r_REG12341_S1 : DFF_X1 port map( D => n36778, CK => CLK, Q => n41094, QN
                           => n_3239);
   clk_r_REG12724_S1 : DFF_X1 port map( D => n36234, CK => CLK, Q => n41093, QN
                           => n_3240);
   clk_r_REG12730_S1 : DFF_X1 port map( D => n36575, CK => CLK, Q => n41092, QN
                           => n_3241);
   clk_r_REG12928_S1 : DFF_X1 port map( D => n36574, CK => CLK, Q => n41091, QN
                           => n_3242);
   clk_r_REG12527_S1 : DFF_X1 port map( D => n36794, CK => CLK, Q => n41090, QN
                           => n_3243);
   clk_r_REG12782_S1 : DFF_X1 port map( D => n36254, CK => CLK, Q => n41089, QN
                           => n_3244);
   clk_r_REG12339_S1 : DFF_X1 port map( D => n36782, CK => CLK, Q => n41088, QN
                           => n_3245);
   clk_r_REG12912_S1 : DFF_X1 port map( D => n36771, CK => CLK, Q => n41087, QN
                           => n_3246);
   clk_r_REG12229_S1 : DFF_X1 port map( D => n35992, CK => CLK, Q => n41086, QN
                           => n_3247);
   clk_r_REG12401_S1 : DFF_X1 port map( D => n36796, CK => CLK, Q => n41085, QN
                           => n_3248);
   clk_r_REG12353_S1 : DFF_X1 port map( D => n36569, CK => CLK, Q => n41084, QN
                           => n_3249);
   clk_r_REG12369_S1 : DFF_X1 port map( D => n36785, CK => CLK, Q => n41083, QN
                           => n_3250);
   clk_r_REG12798_S1 : DFF_X1 port map( D => n36789, CK => CLK, Q => n41082, QN
                           => n_3251);
   clk_r_REG12738_S1 : DFF_X1 port map( D => n36251, CK => CLK, Q => n41081, QN
                           => n_3252);
   clk_r_REG12561_S1 : DFF_X1 port map( D => n36797, CK => CLK, Q => n41080, QN
                           => n_3253);
   clk_r_REG12431_S1 : DFF_X1 port map( D => n36779, CK => CLK, Q => n41079, QN
                           => n_3254);
   clk_r_REG12549_S1 : DFF_X1 port map( D => n36560, CK => CLK, Q => n41078, QN
                           => n_3255);
   clk_r_REG12421_S1 : DFF_X1 port map( D => n36555, CK => CLK, Q => n41077, QN
                           => n_3256);
   clk_r_REG12377_S1 : DFF_X1 port map( D => n36554, CK => CLK, Q => n41076, QN
                           => n_3257);
   clk_r_REG12952_S1 : DFF_X1 port map( D => n36553, CK => CLK, Q => n41075, QN
                           => n_3258);
   clk_r_REG12231_S1 : DFF_X1 port map( D => n35988, CK => CLK, Q => n41074, QN
                           => n_3259);
   clk_r_REG12796_S1 : DFF_X1 port map( D => n35985, CK => CLK, Q => n41073, QN
                           => n_3260);
   clk_r_REG12816_S1 : DFF_X1 port map( D => n35984, CK => CLK, Q => n41072, QN
                           => n_3261);
   clk_r_REG12427_S1 : DFF_X1 port map( D => n36795, CK => CLK, Q => n41071, QN
                           => n_3262);
   clk_r_REG12359_S1 : DFF_X1 port map( D => n36549, CK => CLK, Q => n41070, QN
                           => n_3263);
   clk_r_REG12563_S1 : DFF_X1 port map( D => n36776, CK => CLK, Q => n41069, QN
                           => n_3264);
   clk_r_REG12429_S1 : DFF_X1 port map( D => n36781, CK => CLK, Q => n41068, QN
                           => n_3265);
   clk_r_REG12335_S1 : DFF_X1 port map( D => n36792, CK => CLK, Q => n41067, QN
                           => n_3266);
   clk_r_REG12940_S1 : DFF_X1 port map( D => n36798, CK => CLK, Q => n41066, QN
                           => n_3267);
   clk_r_REG12553_S1 : DFF_X1 port map( D => n36544, CK => CLK, Q => n41065, QN
                           => n_3268);
   clk_r_REG12407_S1 : DFF_X1 port map( D => n36681, CK => CLK, Q => n41064, QN
                           => n_3269);
   clk_r_REG12361_S1 : DFF_X1 port map( D => n36545, CK => CLK, Q => n41063, QN
                           => n_3270);
   clk_r_REG12936_S1 : DFF_X1 port map( D => n36546, CK => CLK, Q => n41062, QN
                           => n_3271);
   clk_r_REG12233_S1 : DFF_X1 port map( D => n35983, CK => CLK, Q => n41061, QN
                           => n_3272);
   clk_r_REG12818_S1 : DFF_X1 port map( D => n35982, CK => CLK, Q => n41060, QN
                           => n_3273);
   clk_r_REG12820_S1 : DFF_X1 port map( D => n35981, CK => CLK, Q => n41059, QN
                           => n_3274);
   clk_r_REG12756_S1 : DFF_X1 port map( D => n35980, CK => CLK, Q => n41058, QN
                           => n_3275);
   clk_r_REG12551_S1 : DFF_X1 port map( D => n36551, CK => CLK, Q => n41057, QN
                           => n_3276);
   clk_r_REG12419_S1 : DFF_X1 port map( D => n36556, CK => CLK, Q => n41056, QN
                           => n_3277);
   clk_r_REG12357_S1 : DFF_X1 port map( D => n36557, CK => CLK, Q => n41055, QN
                           => n_3278);
   clk_r_REG12934_S1 : DFF_X1 port map( D => n36558, CK => CLK, Q => n41054, QN
                           => n_3279);
   clk_r_REG12708_S1 : DFF_X1 port map( D => n36559, CK => CLK, Q => n41053, QN
                           => n_3280);
   clk_r_REG12822_S1 : DFF_X1 port map( D => n35979, CK => CLK, Q => n41052, QN
                           => n_3281);
   clk_r_REG12758_S1 : DFF_X1 port map( D => n35978, CK => CLK, Q => n41051, QN
                           => n_3282);
   clk_r_REG12547_S1 : DFF_X1 port map( D => n36561, CK => CLK, Q => n41050, QN
                           => n_3283);
   clk_r_REG12417_S1 : DFF_X1 port map( D => n36562, CK => CLK, Q => n41049, QN
                           => n_3284);
   clk_r_REG12355_S1 : DFF_X1 port map( D => n36563, CK => CLK, Q => n41048, QN
                           => n_3285);
   clk_r_REG12932_S1 : DFF_X1 port map( D => n36564, CK => CLK, Q => n41047, QN
                           => n_3286);
   clk_r_REG12824_S1 : DFF_X1 port map( D => n35977, CK => CLK, Q => n41046, QN
                           => n_3287);
   clk_r_REG12760_S1 : DFF_X1 port map( D => n35976, CK => CLK, Q => n41045, QN
                           => n_3288);
   clk_r_REG12826_S1 : DFF_X1 port map( D => n35975, CK => CLK, Q => n41044, QN
                           => n_3289);
   clk_r_REG12545_S1 : DFF_X1 port map( D => n36566, CK => CLK, Q => n41043, QN
                           => n_3290);
   clk_r_REG12762_S1 : DFF_X1 port map( D => n35974, CK => CLK, Q => n41042, QN
                           => n_3291);
   clk_r_REG12415_S1 : DFF_X1 port map( D => n36567, CK => CLK, Q => n41041, QN
                           => n_3292);
   clk_r_REG12930_S1 : DFF_X1 port map( D => n36568, CK => CLK, Q => n41040, QN
                           => n_3293);
   clk_r_REG11490_S1 : DFF_X1 port map( D => n35973, CK => CLK, Q => n41039, QN
                           => n_3294);
   clk_r_REG11492_S1 : DFF_X1 port map( D => n35972, CK => CLK, Q => n41038, QN
                           => n_3295);
   clk_r_REG11454_S1 : DFF_X1 port map( D => n36190, CK => CLK, Q => n41037, QN
                           => n_3296);
   clk_r_REG11456_S1 : DFF_X1 port map( D => n36189, CK => CLK, Q => n41036, QN
                           => n_3297);
   clk_r_REG11494_S1 : DFF_X1 port map( D => n35970, CK => CLK, Q => n41035, QN
                           => n_3298);
   clk_r_REG11496_S1 : DFF_X1 port map( D => n35969, CK => CLK, Q => n41034, QN
                           => n_3299);
   clk_r_REG12166_S1 : DFF_X1 port map( D => n35968, CK => CLK, Q => n41033, QN
                           => n_3300);
   clk_r_REG12168_S1 : DFF_X1 port map( D => n35967, CK => CLK, Q => n41032, QN
                           => n_3301);
   clk_r_REG12842_S1 : DFF_X1 port map( D => n36577, CK => CLK, Q => n41031, QN
                           => n_3302);
   clk_r_REG11969_S1 : DFF_X1 port map( D => n35966, CK => CLK, Q => n41030, QN
                           => n_3303);
   clk_r_REG10916_S1 : DFF_X1 port map( D => n35965, CK => CLK, Q => n41029, QN
                           => n_3304);
   clk_r_REG11971_S1 : DFF_X1 port map( D => n35964, CK => CLK, Q => n41028, QN
                           => n_3305);
   clk_r_REG12994_S1 : DFF_X1 port map( D => n36582, CK => CLK, Q => n41027, QN
                           => n_3306);
   clk_r_REG11667_S1 : DFF_X1 port map( D => n36583, CK => CLK, Q => n41026, QN
                           => n_3307);
   clk_r_REG11410_S1 : DFF_X1 port map( D => n35963, CK => CLK, Q => n41025, QN
                           => n_3308);
   clk_r_REG10918_S1 : DFF_X1 port map( D => n35962, CK => CLK, Q => n41024, QN
                           => n_3309);
   clk_r_REG12291_S1 : DFF_X1 port map( D => n35960, CK => CLK, Q => n41023, QN
                           => n_3310);
   clk_r_REG13208_S1 : DFF_X1 port map( D => n35819, CK => CLK, Q => n41022, QN
                           => n_3311);
   clk_r_REG12487_S1 : DFF_X1 port map( D => n36589, CK => CLK, Q => n41021, QN
                           => n_3312);
   clk_r_REG12485_S1 : DFF_X1 port map( D => n36591, CK => CLK, Q => n41020, QN
                           => n_3313);
   clk_r_REG11851_S1 : DFF_X1 port map( D => n35817, CK => CLK, Q => n41019, QN
                           => n_3314);
   clk_r_REG12617_S1 : DFF_X1 port map( D => n36592, CK => CLK, Q => n41018, QN
                           => n_3315);
   clk_r_REG13359_S1 : DFF_X1 port map( D => n35816, CK => CLK, Q => n41017, QN
                           => n_3316);
   clk_r_REG11665_S1 : DFF_X1 port map( D => n36593, CK => CLK, Q => n41016, QN
                           => n_3317);
   clk_r_REG12840_S1 : DFF_X1 port map( D => n36594, CK => CLK, Q => n41015, QN
                           => n_3318);
   clk_r_REG13361_S1 : DFF_X1 port map( D => n35813, CK => CLK, Q => n41014, QN
                           => n_3319);
   clk_r_REG12319_S1 : DFF_X1 port map( D => n35812, CK => CLK, Q => n41013, QN
                           => n_3320);
   clk_r_REG13363_S1 : DFF_X1 port map( D => n35811, CK => CLK, Q => n41012, QN
                           => n_3321);
   clk_r_REG12124_S1 : DFF_X1 port map( D => n35810, CK => CLK, Q => n41011, QN
                           => n_3322);
   clk_r_REG12615_S1 : DFF_X1 port map( D => n36598, CK => CLK, Q => n41010, QN
                           => n_3323);
   clk_r_REG13150_S1 : DFF_X1 port map( D => n36602, CK => CLK, Q => n41009, QN
                           => n_3324);
   clk_r_REG12990_S1 : DFF_X1 port map( D => n36605, CK => CLK, Q => n41008, QN
                           => n_3325);
   clk_r_REG11999_S1 : DFF_X1 port map( D => n35808, CK => CLK, Q => n41007, QN
                           => n_3326);
   clk_r_REG13056_S1 : DFF_X1 port map( D => n36608, CK => CLK, Q => n41006, QN
                           => n_3327);
   clk_r_REG13210_S1 : DFF_X1 port map( D => n35807, CK => CLK, Q => n41005, QN
                           => n_3328);
   clk_r_REG12894_S1 : DFF_X1 port map( D => n35806, CK => CLK, Q => n41004, QN
                           => n_3329);
   clk_r_REG12194_S1 : DFF_X1 port map( D => n35805, CK => CLK, Q => n41003, QN
                           => n_3330);
   clk_r_REG11853_S1 : DFF_X1 port map( D => n35804, CK => CLK, Q => n41002, QN
                           => n_3331);
   clk_r_REG12128_S1 : DFF_X1 port map( D => n35803, CK => CLK, Q => n41001, QN
                           => n_3332);
   clk_r_REG11384_S1 : DFF_X1 port map( D => n36611, CK => CLK, Q => n41000, QN
                           => n_3333);
   clk_r_REG11855_S1 : DFF_X1 port map( D => n35801, CK => CLK, Q => n40999, QN
                           => n_3334);
   clk_r_REG12481_S1 : DFF_X1 port map( D => n36612, CK => CLK, Q => n40998, QN
                           => n_3335);
   clk_r_REG10952_S1 : DFF_X1 port map( D => n35800, CK => CLK, Q => n40997, QN
                           => n_3336);
   clk_r_REG13054_S1 : DFF_X1 port map( D => n36615, CK => CLK, Q => n40996, QN
                           => n_3337);
   clk_r_REG13052_S1 : DFF_X1 port map( D => n36616, CK => CLK, Q => n40995, QN
                           => n_3338);
   clk_r_REG12130_S1 : DFF_X1 port map( D => n35799, CK => CLK, Q => n40994, QN
                           => n_3339);
   clk_r_REG12261_S1 : DFF_X1 port map( D => n36617, CK => CLK, Q => n40993, QN
                           => n_3340);
   clk_r_REG11713_S1 : DFF_X1 port map( D => n35798, CK => CLK, Q => n40992, QN
                           => n_3341);
   clk_r_REG11438_S1 : DFF_X1 port map( D => n35797, CK => CLK, Q => n40991, QN
                           => n_3342);
   clk_r_REG12607_S1 : DFF_X1 port map( D => n36620, CK => CLK, Q => n40990, QN
                           => n_3343);
   clk_r_REG12988_S1 : DFF_X1 port map( D => n36621, CK => CLK, Q => n40989, QN
                           => n_3344);
   clk_r_REG11661_S1 : DFF_X1 port map( D => n36622, CK => CLK, Q => n40988, QN
                           => n_3345);
   clk_r_REG11715_S1 : DFF_X1 port map( D => n35796, CK => CLK, Q => n40987, QN
                           => n_3346);
   clk_r_REG11659_S1 : DFF_X1 port map( D => n36623, CK => CLK, Q => n40986, QN
                           => n_3347);
   clk_r_REG11695_S1 : DFF_X1 port map( D => n36158, CK => CLK, Q => n40985, QN
                           => n_3348);
   clk_r_REG11693_S1 : DFF_X1 port map( D => n36159, CK => CLK, Q => n40984, QN
                           => n_3349);
   clk_r_REG11657_S1 : DFF_X1 port map( D => n36625, CK => CLK, Q => n40983, QN
                           => n_3350);
   clk_r_REG11765_S1 : DFF_X1 port map( D => n35793, CK => CLK, Q => n40982, QN
                           => n_3351);
   clk_r_REG11625_S1 : DFF_X1 port map( D => n35792, CK => CLK, Q => n40981, QN
                           => n_3352);
   clk_r_REG11910_S1 : DFF_X1 port map( D => n35791, CK => CLK, Q => n40980, QN
                           => n_3353);
   clk_r_REG11547_S1 : DFF_X1 port map( D => n35790, CK => CLK, Q => n40979, QN
                           => n_3354);
   clk_r_REG11627_S1 : DFF_X1 port map( D => n35788, CK => CLK, Q => n40978, QN
                           => n_3355);
   clk_r_REG11767_S1 : DFF_X1 port map( D => n35787, CK => CLK, Q => n40977, QN
                           => n_3356);
   clk_r_REG12699_S1 : DFF_X1 port map( D => n35786, CK => CLK, Q => n40976, QN
                           => n_3357);
   clk_r_REG11647_S1 : DFF_X1 port map( D => n35784, CK => CLK, Q => n40975, QN
                           => n_3358);
   clk_r_REG12701_S1 : DFF_X1 port map( D => n35783, CK => CLK, Q => n40974, QN
                           => n_3359);
   clk_r_REG11326_S1 : DFF_X1 port map( D => n35782, CK => CLK, Q => n40973, QN
                           => n_3360);
   clk_r_REG11328_S1 : DFF_X1 port map( D => n35781, CK => CLK, Q => n40972, QN
                           => n_3361);
   clk_r_REG11787_S1 : DFF_X1 port map( D => n35780, CK => CLK, Q => n40971, QN
                           => n_3362);
   clk_r_REG11549_S1 : DFF_X1 port map( D => n35779, CK => CLK, Q => n40970, QN
                           => n_3363);
   clk_r_REG11348_S1 : DFF_X1 port map( D => n35778, CK => CLK, Q => n40969, QN
                           => n_3364);
   clk_r_REG11569_S1 : DFF_X1 port map( D => n35777, CK => CLK, Q => n40968, QN
                           => n_3365);
   clk_r_REG11350_S1 : DFF_X1 port map( D => n35776, CK => CLK, Q => n40967, QN
                           => n_3366);
   clk_r_REG12675_S1 : DFF_X1 port map( D => n36161, CK => CLK, Q => n40966, QN
                           => n_3367);
   clk_r_REG11525_S1 : DFF_X1 port map( D => n36163, CK => CLK, Q => n40965, QN
                           => n_3368);
   clk_r_REG11304_S1 : DFF_X1 port map( D => n36164, CK => CLK, Q => n40964, QN
                           => n_3369);
   clk_r_REG11914_S1 : DFF_X1 port map( D => n35773, CK => CLK, Q => n40963, QN
                           => n_3370);
   clk_r_REG11605_S1 : DFF_X1 port map( D => n36165, CK => CLK, Q => n40962, QN
                           => n_3371);
   clk_r_REG11789_S1 : DFF_X1 port map( D => n35772, CK => CLK, Q => n40961, QN
                           => n_3372);
   clk_r_REG11934_S1 : DFF_X1 port map( D => n35770, CK => CLK, Q => n40960, QN
                           => n_3373);
   clk_r_REG11747_S1 : DFF_X1 port map( D => n36166, CK => CLK, Q => n40959, QN
                           => n_3374);
   clk_r_REG12695_S1 : DFF_X1 port map( D => n35820, CK => CLK, Q => n40958, QN
                           => n_3375);
   clk_r_REG12703_S1 : DFF_X1 port map( D => n35771, CK => CLK, Q => n40957, QN
                           => n_3376);
   clk_r_REG11888_S1 : DFF_X1 port map( D => n36167, CK => CLK, Q => n40956, QN
                           => n_3377);
   clk_r_REG11912_S1 : DFF_X1 port map( D => n35775, CK => CLK, Q => n40955, QN
                           => n_3378);
   clk_r_REG11745_S1 : DFF_X1 port map( D => n36168, CK => CLK, Q => n40954, QN
                           => n_3379);
   clk_r_REG11603_S1 : DFF_X1 port map( D => n36169, CK => CLK, Q => n40953, QN
                           => n_3380);
   clk_r_REG11302_S1 : DFF_X1 port map( D => n36170, CK => CLK, Q => n40952, QN
                           => n_3381);
   clk_r_REG11523_S1 : DFF_X1 port map( D => n36171, CK => CLK, Q => n40951, QN
                           => n_3382);
   clk_r_REG11543_S1 : DFF_X1 port map( D => n35815, CK => CLK, Q => n40950, QN
                           => n_3383);
   clk_r_REG11886_S1 : DFF_X1 port map( D => n36172, CK => CLK, Q => n40949, QN
                           => n_3384);
   clk_r_REG12661_S1 : DFF_X1 port map( D => n36174, CK => CLK, Q => n40948, QN
                           => n_3385);
   clk_r_REG11623_S1 : DFF_X1 port map( D => n35818, CK => CLK, Q => n40947, QN
                           => n_3386);
   clk_r_REG13248_S1 : DFF_X1 port map( D => n36176, CK => CLK, Q => n40946, QN
                           => n_3387);
   clk_r_REG13246_S1 : DFF_X1 port map( D => n36177, CK => CLK, Q => n40945, QN
                           => n_3388);
   clk_r_REG13238_S1 : DFF_X1 port map( D => n36225, CK => CLK, Q => n40944, QN
                           => n_3389);
   clk_r_REG13244_S1 : DFF_X1 port map( D => n36179, CK => CLK, Q => n40943, QN
                           => n_3390);
   clk_r_REG13242_S1 : DFF_X1 port map( D => n36181, CK => CLK, Q => n40942, QN
                           => n_3391);
   clk_r_REG13272_S1 : DFF_X1 port map( D => n35821, CK => CLK, Q => n40941, QN
                           => n_3392);
   clk_r_REG13240_S1 : DFF_X1 port map( D => n36183, CK => CLK, Q => n40940, QN
                           => n_3393);
   clk_r_REG10351_S1 : DFF_X1 port map( D => n36399, CK => CLK, Q => n40939, QN
                           => n_3394);
   clk_r_REG13104_S1 : DFF_X1 port map( D => n36186, CK => CLK, Q => n40938, QN
                           => n_3395);
   clk_r_REG13124_S1 : DFF_X1 port map( D => n36187, CK => CLK, Q => n40937, QN
                           => n_3396);
   clk_r_REG11884_S1 : DFF_X1 port map( D => n36191, CK => CLK, Q => n40936, QN
                           => n_3397);
   clk_r_REG13102_S1 : DFF_X1 port map( D => n36192, CK => CLK, Q => n40935, QN
                           => n_3398);
   clk_r_REG13160_S1 : DFF_X1 port map( D => n36193, CK => CLK, Q => n40934, QN
                           => n_3399);
   clk_r_REG13146_S1 : DFF_X1 port map( D => n35826, CK => CLK, Q => n40933, QN
                           => n_3400);
   clk_r_REG11300_S1 : DFF_X1 port map( D => n36194, CK => CLK, Q => n40932, QN
                           => n_3401);
   clk_r_REG13100_S1 : DFF_X1 port map( D => n36195, CK => CLK, Q => n40931, QN
                           => n_3402);
   clk_r_REG11882_S1 : DFF_X1 port map( D => n36196, CK => CLK, Q => n40930, QN
                           => n_3403);
   clk_r_REG13098_S1 : DFF_X1 port map( D => n36197, CK => CLK, Q => n40929, QN
                           => n_3404);
   clk_r_REG11298_S1 : DFF_X1 port map( D => n36198, CK => CLK, Q => n40928, QN
                           => n_3405);
   clk_r_REG10764_S1 : DFF_X1 port map( D => n36404, CK => CLK, Q => n40927, QN
                           => n_3406);
   clk_r_REG11743_S1 : DFF_X1 port map( D => n36200, CK => CLK, Q => n40926, QN
                           => n_3407);
   clk_r_REG11953_S1 : DFF_X1 port map( D => n36201, CK => CLK, Q => n40925, QN
                           => n_3408);
   clk_r_REG11779_S1 : DFF_X1 port map( D => n36202, CK => CLK, Q => n40924, QN
                           => n_3409);
   clk_r_REG11930_S1 : DFF_X1 port map( D => n36203, CK => CLK, Q => n40923, QN
                           => n_3410);
   clk_r_REG11928_S1 : DFF_X1 port map( D => n36204, CK => CLK, Q => n40922, QN
                           => n_3411);
   clk_r_REG11880_S1 : DFF_X1 port map( D => n36205, CK => CLK, Q => n40921, QN
                           => n_3412);
   clk_r_REG11878_S1 : DFF_X1 port map( D => n36206, CK => CLK, Q => n40920, QN
                           => n_3413);
   clk_r_REG12659_S1 : DFF_X1 port map( D => n36207, CK => CLK, Q => n40919, QN
                           => n_3414);
   clk_r_REG11344_S1 : DFF_X1 port map( D => n36208, CK => CLK, Q => n40918, QN
                           => n_3415);
   clk_r_REG10696_S1 : DFF_X1 port map( D => n36426, CK => CLK, Q => n40917, QN
                           => n_3416);
   clk_r_REG11601_S1 : DFF_X1 port map( D => n36209, CK => CLK, Q => n40916, QN
                           => n_3417);
   clk_r_REG11777_S1 : DFF_X1 port map( D => n36210, CK => CLK, Q => n40915, QN
                           => n_3418);
   clk_r_REG11741_S1 : DFF_X1 port map( D => n36211, CK => CLK, Q => n40914, QN
                           => n_3419);
   clk_r_REG11908_S1 : DFF_X1 port map( D => n35839, CK => CLK, Q => n40913, QN
                           => n_3420);
   clk_r_REG11342_S1 : DFF_X1 port map( D => n36212, CK => CLK, Q => n40912, QN
                           => n_3421);
   clk_r_REG11296_S1 : DFF_X1 port map( D => n36213, CK => CLK, Q => n40911, QN
                           => n_3422);
   clk_r_REG11599_S1 : DFF_X1 port map( D => n36214, CK => CLK, Q => n40910, QN
                           => n_3423);
   clk_r_REG11629_S1 : DFF_X1 port map( D => n36490, CK => CLK, Q => n40909, QN
                           => n_3424);
   clk_r_REG11645_S1 : DFF_X1 port map( D => n35841, CK => CLK, Q => n40908, QN
                           => n_3425);
   clk_r_REG11597_S1 : DFF_X1 port map( D => n36215, CK => CLK, Q => n40907, QN
                           => n_3426);
   clk_r_REG11739_S1 : DFF_X1 port map( D => n36216, CK => CLK, Q => n40906, QN
                           => n_3427);
   clk_r_REG11294_S1 : DFF_X1 port map( D => n36218, CK => CLK, Q => n40905, QN
                           => n_3428);
   clk_r_REG12024_S1 : DFF_X1 port map( D => n36219, CK => CLK, Q => n40904, QN
                           => n_3429);
   clk_r_REG11737_S1 : DFF_X1 port map( D => n36220, CK => CLK, Q => n40903, QN
                           => n_3430);
   clk_r_REG11763_S1 : DFF_X1 port map( D => n35846, CK => CLK, Q => n40902, QN
                           => n_3431);
   clk_r_REG10866_S1 : DFF_X1 port map( D => n36442, CK => CLK, Q => n40901, QN
                           => n_3432);
   clk_r_REG11324_S1 : DFF_X1 port map( D => n35848, CK => CLK, Q => n40900, QN
                           => n_3433);
   clk_r_REG11595_S1 : DFF_X1 port map( D => n36221, CK => CLK, Q => n40899, QN
                           => n_3434);
   clk_r_REG12657_S1 : DFF_X1 port map( D => n36222, CK => CLK, Q => n40898, QN
                           => n_3435);
   clk_r_REG11521_S1 : DFF_X1 port map( D => n36223, CK => CLK, Q => n40897, QN
                           => n_3436);
   clk_r_REG11593_S1 : DFF_X1 port map( D => n36224, CK => CLK, Q => n40896, QN
                           => n_3437);
   clk_r_REG11591_S1 : DFF_X1 port map( D => n36227, CK => CLK, Q => n40895, QN
                           => n_3438);
   clk_r_REG11517_S1 : DFF_X1 port map( D => n36240, CK => CLK, Q => n40894, QN
                           => n_3439);
   clk_r_REG12020_S1 : DFF_X1 port map( D => n36242, CK => CLK, Q => n40893, QN
                           => n_3440);
   clk_r_REG12046_S1 : DFF_X1 port map( D => n36243, CK => CLK, Q => n40892, QN
                           => n_3441);
   clk_r_REG10620_S1 : DFF_X1 port map( D => n36450, CK => CLK, Q => n40891, QN
                           => n_3442);
   clk_r_REG12673_S1 : DFF_X1 port map( D => n36247, CK => CLK, Q => n40890, QN
                           => n_3443);
   clk_r_REG11561_S1 : DFF_X1 port map( D => n36250, CK => CLK, Q => n40889, QN
                           => n_3444);
   clk_r_REG12064_S1 : DFF_X1 port map( D => n35850, CK => CLK, Q => n40888, QN
                           => n_3445);
   clk_r_REG12022_S1 : DFF_X1 port map( D => n36229, CK => CLK, Q => n40887, QN
                           => n_3446);
   clk_r_REG11563_S1 : DFF_X1 port map( D => n36249, CK => CLK, Q => n40886, QN
                           => n_3447);
   clk_r_REG12671_S1 : DFF_X1 port map( D => n36256, CK => CLK, Q => n40885, QN
                           => n_3448);
   clk_r_REG12697_S1 : DFF_X1 port map( D => n35814, CK => CLK, Q => n40884, QN
                           => n_3449);
   clk_r_REG10417_S1 : DFF_X1 port map( D => n36455, CK => CLK, Q => n40883, QN
                           => n_3450);
   clk_r_REG12018_S1 : DFF_X1 port map( D => n36258, CK => CLK, Q => n40882, QN
                           => n_3451);
   clk_r_REG12655_S1 : DFF_X1 port map( D => n36245, CK => CLK, Q => n40881, QN
                           => n_3452);
   clk_r_REG12653_S1 : DFF_X1 port map( D => n36246, CK => CLK, Q => n40880, QN
                           => n_3453);
   clk_r_REG11519_S1 : DFF_X1 port map( D => n36228, CK => CLK, Q => n40879, QN
                           => n_3454);
   clk_r_REG11545_S1 : DFF_X1 port map( D => n35802, CK => CLK, Q => n40878, QN
                           => n_3455);
   clk_r_REG11515_S1 : DFF_X1 port map( D => n36255, CK => CLK, Q => n40877, QN
                           => n_3456);
   clk_r_REG10807_S1 : DFF_X1 port map( D => n36470, CK => CLK, Q => n40876, QN
                           => n_3457);
   clk_r_REG10323_S1 : DFF_X1 port map( D => n36504, CK => CLK, Q => n40875, QN
                           => n_3458);
   clk_r_REG13222_S1 : DFF_X1 port map( D => n36499, CK => CLK, Q => n40874, QN
                           => n_3459);
   clk_r_REG13274_S1 : DFF_X1 port map( D => n35795, CK => CLK, Q => n40873, QN
                           => n_3460);
   clk_r_REG13270_S1 : DFF_X1 port map( D => n35871, CK => CLK, Q => n40872, QN
                           => n_3461);
   clk_r_REG13236_S1 : DFF_X1 port map( D => n36226, CK => CLK, Q => n40871, QN
                           => n_3462);
   clk_r_REG13276_S1 : DFF_X1 port map( D => n35789, CK => CLK, Q => n40870, QN
                           => n_3463);
   clk_r_REG13365_S1 : DFF_X1 port map( D => n35785, CK => CLK, Q => n40869, QN
                           => n_3464);
   clk_r_REG13323_S1 : DFF_X1 port map( D => n36480, CK => CLK, Q => n40868, QN
                           => n_3465);
   clk_r_REG13347_S1 : DFF_X1 port map( D => n36241, CK => CLK, Q => n40867, QN
                           => n_3466);
   clk_r_REG13307_S1 : DFF_X1 port map( D => n36709, CK => CLK, Q => n40866, QN
                           => n_3467);
   clk_r_REG13309_S1 : DFF_X1 port map( D => n36706, CK => CLK, Q => n40865, QN
                           => n_3468);
   clk_r_REG12271_S1 : DFF_X1 port map( D => n36253, CK => CLK, Q => n40864, QN
                           => n_3469);
   clk_r_REG12321_S1 : DFF_X1 port map( D => n35794, CK => CLK, Q => n40863, QN
                           => n_3470);
   clk_r_REG12299_S1 : DFF_X1 port map( D => n36483, CK => CLK, Q => n40862, QN
                           => n_3471);
   clk_r_REG12275_S1 : DFF_X1 port map( D => n36235, CK => CLK, Q => n40861, QN
                           => n_3472);
   clk_r_REG12277_S1 : DFF_X1 port map( D => n36233, CK => CLK, Q => n40860, QN
                           => n_3473);
   clk_r_REG12279_S1 : DFF_X1 port map( D => n36232, CK => CLK, Q => n40859, QN
                           => n_3474);
   clk_r_REG12273_S1 : DFF_X1 port map( D => n36252, CK => CLK, Q => n40858, QN
                           => n_3475);
   clk_r_REG12864_S1 : DFF_X1 port map( D => n36230, CK => CLK, Q => n40857, QN
                           => n_3476);
   clk_r_REG12834_S1 : DFF_X1 port map( D => n36685, CK => CLK, Q => n40856, QN
                           => n_3477);
   clk_r_REG12872_S1 : DFF_X1 port map( D => n36478, CK => CLK, Q => n40855, QN
                           => n_3478);
   clk_r_REG12856_S1 : DFF_X1 port map( D => n36248, CK => CLK, Q => n40854, QN
                           => n_3479);
   clk_r_REG12858_S1 : DFF_X1 port map( D => n36244, CK => CLK, Q => n40853, QN
                           => n_3480);
   clk_r_REG10309_S1 : DFF_X1 port map( D => n36719, CK => CLK, Q => n40852, QN
                           => n_3481);
   clk_r_REG12860_S1 : DFF_X1 port map( D => n36239, CK => CLK, Q => n40851, QN
                           => n_3482);
   clk_r_REG12862_S1 : DFF_X1 port map( D => n36238, CK => CLK, Q => n40850, QN
                           => n_3483);
   clk_r_REG13331_S1 : DFF_X1 port map( D => n36231, CK => CLK, Q => n40849, QN
                           => n_3484);
   clk_r_REG10391_S1 : DFF_X1 port map( D => n36716, CK => CLK, Q => n40848, QN
                           => n_3485);
   clk_r_REG13172_S1 : DFF_X1 port map( D => n36083, CK => CLK, Q => n40847, QN
                           => n_3486);
   clk_r_REG11857_S1 : DFF_X1 port map( D => n35774, CK => CLK, Q => n40846, QN
                           => n_3487);
   clk_r_REG13188_S1 : DFF_X1 port map( D => n35847, CK => CLK, Q => n40845, QN
                           => n_3488);
   clk_r_REG13152_S1 : DFF_X1 port map( D => n36484, CK => CLK, Q => n40844, QN
                           => n_3489);
   clk_r_REG13170_S1 : DFF_X1 port map( D => n36084, CK => CLK, Q => n40843, QN
                           => n_3490);
   clk_r_REG13168_S1 : DFF_X1 port map( D => n36085, CK => CLK, Q => n40842, QN
                           => n_3491);
   clk_r_REG13166_S1 : DFF_X1 port map( D => n36086, CK => CLK, Q => n40841, QN
                           => n_3492);
   clk_r_REG13164_S1 : DFF_X1 port map( D => n36087, CK => CLK, Q => n40840, QN
                           => n_3493);
   clk_r_REG10712_S1 : DFF_X1 port map( D => n36486, CK => CLK, Q => n40839, QN
                           => n_3494);
   clk_r_REG11813_S1 : DFF_X1 port map( D => n36088, CK => CLK, Q => n40838, QN
                           => n_3495);
   clk_r_REG13335_S1 : DFF_X1 port map( D => n36089, CK => CLK, Q => n40837, QN
                           => n_3496);
   clk_r_REG11811_S1 : DFF_X1 port map( D => n36090, CK => CLK, Q => n40836, QN
                           => n_3497);
   clk_r_REG11809_S1 : DFF_X1 port map( D => n36091, CK => CLK, Q => n40835, QN
                           => n_3498);
   clk_r_REG11839_S1 : DFF_X1 port map( D => n36092, CK => CLK, Q => n40834, QN
                           => n_3499);
   clk_r_REG11807_S1 : DFF_X1 port map( D => n36093, CK => CLK, Q => n40833, QN
                           => n_3500);
   clk_r_REG11837_S1 : DFF_X1 port map( D => n36094, CK => CLK, Q => n40832, QN
                           => n_3501);
   clk_r_REG12986_S1 : DFF_X1 port map( D => n36624, CK => CLK, Q => n40831, QN
                           => n_3502);
   clk_r_REG13128_S1 : DFF_X1 port map( D => n36095, CK => CLK, Q => n40830, QN
                           => n_3503);
   clk_r_REG12142_S1 : DFF_X1 port map( D => n36474, CK => CLK, Q => n40829, QN
                           => n_3504);
   clk_r_REG12156_S1 : DFF_X1 port map( D => n36096, CK => CLK, Q => n40828, QN
                           => n_3505);
   clk_r_REG12154_S1 : DFF_X1 port map( D => n36097, CK => CLK, Q => n40827, QN
                           => n_3506);
   clk_r_REG12152_S1 : DFF_X1 port map( D => n36098, CK => CLK, Q => n40826, QN
                           => n_3507);
   clk_r_REG12136_S1 : DFF_X1 port map( D => n36707, CK => CLK, Q => n40825, QN
                           => n_3508);
   clk_r_REG12150_S1 : DFF_X1 port map( D => n36099, CK => CLK, Q => n40824, QN
                           => n_3509);
   clk_r_REG12978_S1 : DFF_X1 port map( D => n36711, CK => CLK, Q => n40823, QN
                           => n_3510);
   clk_r_REG12283_S1 : DFF_X1 port map( D => n36100, CK => CLK, Q => n40822, QN
                           => n_3511);
   clk_r_REG12182_S1 : DFF_X1 port map( D => n36101, CK => CLK, Q => n40821, QN
                           => n_3512);
   clk_r_REG12138_S1 : DFF_X1 port map( D => n36565, CK => CLK, Q => n40820, QN
                           => n_3513);
   clk_r_REG12092_S1 : DFF_X1 port map( D => n36102, CK => CLK, Q => n40819, QN
                           => n_3514);
   clk_r_REG10542_S1 : DFF_X1 port map( D => n36713, CK => CLK, Q => n40818, QN
                           => n_3515);
   clk_r_REG12090_S1 : DFF_X1 port map( D => n36103, CK => CLK, Q => n40817, QN
                           => n_3516);
   clk_r_REG12088_S1 : DFF_X1 port map( D => n36104, CK => CLK, Q => n40816, QN
                           => n_3517);
   clk_r_REG12086_S1 : DFF_X1 port map( D => n36105, CK => CLK, Q => n40815, QN
                           => n_3518);
   clk_r_REG13060_S1 : DFF_X1 port map( D => n36548, CK => CLK, Q => n40814, QN
                           => n_3519);
   clk_r_REG12489_S1 : DFF_X1 port map( D => n36547, CK => CLK, Q => n40813, QN
                           => n_3520);
   clk_r_REG13016_S1 : DFF_X1 port map( D => n36552, CK => CLK, Q => n40812, QN
                           => n_3521);
   clk_r_REG12084_S1 : DFF_X1 port map( D => n36106, CK => CLK, Q => n40811, QN
                           => n_3522);
   clk_r_REG12126_S1 : DFF_X1 port map( D => n35809, CK => CLK, Q => n40810, QN
                           => n_3523);
   clk_r_REG12070_S1 : DFF_X1 port map( D => n36465, CK => CLK, Q => n40809, QN
                           => n_3524);
   clk_r_REG12996_S1 : DFF_X1 port map( D => n36570, CK => CLK, Q => n40808, QN
                           => n_3525);
   clk_r_REG10457_S1 : DFF_X1 port map( D => n36864, CK => CLK, Q => n40807, QN
                           => n_3526);
   clk_r_REG12495_S1 : DFF_X1 port map( D => n36775, CK => CLK, Q => n40806, QN
                           => n_3527);
   clk_r_REG12465_S1 : DFF_X1 port map( D => n36766, CK => CLK, Q => n40805, QN
                           => n_3528);
   clk_r_REG12467_S1 : DFF_X1 port map( D => n36765, CK => CLK, Q => n40804, QN
                           => n_3529);
   clk_r_REG12992_S1 : DFF_X1 port map( D => n36597, CK => CLK, Q => n40803, QN
                           => n_3530);
   clk_r_REG11959_S1 : DFF_X1 port map( D => n36107, CK => CLK, Q => n40802, QN
                           => n_3531);
   clk_r_REG11989_S1 : DFF_X1 port map( D => n36108, CK => CLK, Q => n40801, QN
                           => n_3532);
   clk_r_REG11947_S1 : DFF_X1 port map( D => n36456, CK => CLK, Q => n40800, QN
                           => n_3533);
   clk_r_REG12048_S1 : DFF_X1 port map( D => n36109, CK => CLK, Q => n40799, QN
                           => n_3534);
   clk_r_REG12001_S1 : DFF_X1 port map( D => n35769, CK => CLK, Q => n40798, QN
                           => n_3535);
   clk_r_REG11941_S1 : DFF_X1 port map( D => n36747, CK => CLK, Q => n40797, QN
                           => n_3536);
   clk_r_REG11957_S1 : DFF_X1 port map( D => n36110, CK => CLK, Q => n40796, QN
                           => n_3537);
   clk_r_REG11987_S1 : DFF_X1 port map( D => n36111, CK => CLK, Q => n40795, QN
                           => n_3538);
   clk_r_REG12473_S1 : DFF_X1 port map( D => n36742, CK => CLK, Q => n40794, QN
                           => n_3539);
   clk_r_REG12479_S1 : DFF_X1 port map( D => n36614, CK => CLK, Q => n40793, QN
                           => n_3540);
   clk_r_REG13034_S1 : DFF_X1 port map( D => n36741, CK => CLK, Q => n40792, QN
                           => n_3541);
   clk_r_REG13036_S1 : DFF_X1 port map( D => n36740, CK => CLK, Q => n40791, QN
                           => n_3542);
   clk_r_REG13038_S1 : DFF_X1 port map( D => n36738, CK => CLK, Q => n40790, QN
                           => n_3543);
   clk_r_REG12976_S1 : DFF_X1 port map( D => n36737, CK => CLK, Q => n40789, QN
                           => n_3544);
   clk_r_REG10359_S1 : DFF_X1 port map( D => n36852, CK => CLK, Q => n40788, QN
                           => n_3545);
   clk_r_REG13050_S1 : DFF_X1 port map( D => n36627, CK => CLK, Q => n40787, QN
                           => n_3546);
   clk_r_REG13040_S1 : DFF_X1 port map( D => n36732, CK => CLK, Q => n40786, QN
                           => n_3547);
   clk_r_REG10924_S1 : DFF_X1 port map( D => n35849, CK => CLK, Q => n40785, QN
                           => n_3548);
   clk_r_REG10892_S1 : DFF_X1 port map( D => n36451, CK => CLK, Q => n40784, QN
                           => n_3549);
   clk_r_REG10940_S1 : DFF_X1 port map( D => n36112, CK => CLK, Q => n40783, QN
                           => n_3550);
   clk_r_REG10906_S1 : DFF_X1 port map( D => n36113, CK => CLK, Q => n40782, QN
                           => n_3551);
   clk_r_REG10904_S1 : DFF_X1 port map( D => n36114, CK => CLK, Q => n40781, QN
                           => n_3552);
   clk_r_REG10902_S1 : DFF_X1 port map( D => n36115, CK => CLK, Q => n40780, QN
                           => n_3553);
   clk_r_REG10938_S1 : DFF_X1 port map( D => n36116, CK => CLK, Q => n40779, QN
                           => n_3554);
   clk_r_REG10900_S1 : DFF_X1 port map( D => n36117, CK => CLK, Q => n40778, QN
                           => n_3555);
   clk_r_REG12591_S1 : DFF_X1 port map( D => n36729, CK => CLK, Q => n40777, QN
                           => n_3556);
   clk_r_REG12593_S1 : DFF_X1 port map( D => n36727, CK => CLK, Q => n40776, QN
                           => n_3557);
   clk_r_REG12629_S1 : DFF_X1 port map( D => n36723, CK => CLK, Q => n40775, QN
                           => n_3558);
   clk_r_REG12595_S1 : DFF_X1 port map( D => n36720, CK => CLK, Q => n40774, QN
                           => n_3559);
   clk_r_REG12605_S1 : DFF_X1 port map( D => n36648, CK => CLK, Q => n40773, QN
                           => n_3560);
   clk_r_REG12585_S1 : DFF_X1 port map( D => n36800, CK => CLK, Q => n40772, QN
                           => n_3561);
   clk_r_REG12603_S1 : DFF_X1 port map( D => n36652, CK => CLK, Q => n40771, QN
                           => n_3562);
   clk_r_REG11382_S1 : DFF_X1 port map( D => n36654, CK => CLK, Q => n40770, QN
                           => n_3563);
   clk_r_REG11404_S1 : DFF_X1 port map( D => n36118, CK => CLK, Q => n40769, QN
                           => n_3564);
   clk_r_REG11390_S1 : DFF_X1 port map( D => n36443, CK => CLK, Q => n40768, QN
                           => n_3565);
   clk_r_REG11402_S1 : DFF_X1 port map( D => n36119, CK => CLK, Q => n40767, QN
                           => n_3566);
   clk_r_REG11400_S1 : DFF_X1 port map( D => n36120, CK => CLK, Q => n40766, QN
                           => n_3567);
   clk_r_REG11398_S1 : DFF_X1 port map( D => n36121, CK => CLK, Q => n40765, QN
                           => n_3568);
   clk_r_REG11424_S1 : DFF_X1 port map( D => n36122, CK => CLK, Q => n40764, QN
                           => n_3569);
   clk_r_REG11396_S1 : DFF_X1 port map( D => n36123, CK => CLK, Q => n40763, QN
                           => n_3570);
   clk_r_REG12120_S1 : DFF_X1 port map( D => n35845, CK => CLK, Q => n40762, QN
                           => n_3571);
   clk_r_REG11977_S1 : DFF_X1 port map( D => n35844, CK => CLK, Q => n40761, QN
                           => n_3572);
   clk_r_REG11847_S1 : DFF_X1 port map( D => n35843, CK => CLK, Q => n40760, QN
                           => n_3573);
   clk_r_REG13080_S1 : DFF_X1 port map( D => n36636, CK => CLK, Q => n40759, QN
                           => n_3574);
   clk_r_REG12475_S1 : DFF_X1 port map( D => n36739, CK => CLK, Q => n40758, QN
                           => n_3575);
   clk_r_REG12890_S1 : DFF_X1 port map( D => n35842, CK => CLK, Q => n40757, QN
                           => n_3576);
   clk_r_REG12190_S1 : DFF_X1 port map( D => n35840, CK => CLK, Q => n40756, QN
                           => n_3577);
   clk_r_REG10936_S1 : DFF_X1 port map( D => n36124, CK => CLK, Q => n40755, QN
                           => n_3578);
   clk_r_REG10344_S1 : DFF_X1 port map( D => n36684, CK => CLK, Q => n40754, QN
                           => n_3579);
   clk_r_REG11422_S1 : DFF_X1 port map( D => n36125, CK => CLK, Q => n40753, QN
                           => n_3580);
   clk_r_REG11805_S1 : DFF_X1 port map( D => n36126, CK => CLK, Q => n40752, QN
                           => n_3581);
   clk_r_REG12601_S1 : DFF_X1 port map( D => n36664, CK => CLK, Q => n40751, QN
                           => n_3582);
   clk_r_REG13355_S1 : DFF_X1 port map( D => n35838, CK => CLK, Q => n40750, QN
                           => n_3583);
   clk_r_REG12066_S1 : DFF_X1 port map( D => n35837, CK => CLK, Q => n40749, QN
                           => n_3584);
   clk_r_REG12134_S1 : DFF_X1 port map( D => n36756, CK => CLK, Q => n40748, QN
                           => n_3585);
   clk_r_REG12315_S1 : DFF_X1 port map( D => n35836, CK => CLK, Q => n40747, QN
                           => n_3586);
   clk_r_REG13030_S1 : DFF_X1 port map( D => n36760, CK => CLK, Q => n40746, QN
                           => n_3587);
   clk_r_REG12082_S1 : DFF_X1 port map( D => n36127, CK => CLK, Q => n40745, QN
                           => n_3588);
   clk_r_REG12192_S1 : DFF_X1 port map( D => n35835, CK => CLK, Q => n40744, QN
                           => n_3589);
   clk_r_REG12587_S1 : DFF_X1 port map( D => n36791, CK => CLK, Q => n40743, QN
                           => n_3590);
   clk_r_REG12122_S1 : DFF_X1 port map( D => n35834, CK => CLK, Q => n40742, QN
                           => n_3591);
   clk_r_REG11380_S1 : DFF_X1 port map( D => n36661, CK => CLK, Q => n40741, QN
                           => n_3592);
   clk_r_REG11997_S1 : DFF_X1 port map( D => n35833, CK => CLK, Q => n40740, QN
                           => n_3593);
   clk_r_REG12497_S1 : DFF_X1 port map( D => n36679, CK => CLK, Q => n40739, QN
                           => n_3594);
   clk_r_REG12040_S1 : DFF_X1 port map( D => n36666, CK => CLK, Q => n40738, QN
                           => n_3595);
   clk_r_REG12880_S1 : DFF_X1 port map( D => n36128, CK => CLK, Q => n40737, QN
                           => n_3596);
   clk_r_REG13206_S1 : DFF_X1 port map( D => n35832, CK => CLK, Q => n40736, QN
                           => n_3597);
   clk_r_REG10946_S1 : DFF_X1 port map( D => n35831, CK => CLK, Q => n40735, QN
                           => n_3598);
   clk_r_REG13144_S1 : DFF_X1 port map( D => n35830, CK => CLK, Q => n40734, QN
                           => n_3599);
   clk_r_REG11436_S1 : DFF_X1 port map( D => n35829, CK => CLK, Q => n40733, QN
                           => n_3600);
   clk_r_REG11849_S1 : DFF_X1 port map( D => n35828, CK => CLK, Q => n40732, QN
                           => n_3601);
   clk_r_REG13349_S1 : DFF_X1 port map( D => n36129, CK => CLK, Q => n40731, QN
                           => n_3602);
   clk_r_REG10948_S1 : DFF_X1 port map( D => n35827, CK => CLK, Q => n40730, QN
                           => n_3603);
   clk_r_REG12309_S1 : DFF_X1 port map( D => n36130, CK => CLK, Q => n40729, QN
                           => n_3604);
   clk_r_REG13202_S1 : DFF_X1 port map( D => n36131, CK => CLK, Q => n40728, QN
                           => n_3605);
   clk_r_REG13126_S1 : DFF_X1 port map( D => n36132, CK => CLK, Q => n40727, QN
                           => n_3606);
   clk_r_REG13162_S1 : DFF_X1 port map( D => n36133, CK => CLK, Q => n40726, QN
                           => n_3607);
   clk_r_REG12028_S1 : DFF_X1 port map( D => n36134, CK => CLK, Q => n40725, QN
                           => n_3608);
   clk_r_REG12317_S1 : DFF_X1 port map( D => n35825, CK => CLK, Q => n40724, QN
                           => n_3609);
   clk_r_REG13357_S1 : DFF_X1 port map( D => n35824, CK => CLK, Q => n40723, QN
                           => n_3610);
   clk_r_REG12892_S1 : DFF_X1 port map( D => n35823, CK => CLK, Q => n40722, QN
                           => n_3611);
   clk_r_REG12637_S1 : DFF_X1 port map( D => n36541, CK => CLK, Q => n40721, QN
                           => n_3612);
   clk_r_REG12509_S1 : DFF_X1 port map( D => n36540, CK => CLK, Q => n40720, QN
                           => n_3613);
   clk_r_REG13082_S1 : DFF_X1 port map( D => n36536, CK => CLK, Q => n40719, QN
                           => n_3614);
   clk_r_REG10950_S1 : DFF_X1 port map( D => n35822, CK => CLK, Q => n40718, QN
                           => n_3615);
   clk_r_REG11955_S1 : DFF_X1 port map( D => n36135, CK => CLK, Q => n40717, QN
                           => n_3616);
   clk_r_REG12080_S1 : DFF_X1 port map( D => n36136, CK => CLK, Q => n40716, QN
                           => n_3617);
   clk_r_REG12870_S1 : DFF_X1 port map( D => n35870, CK => CLK, Q => n40715, QN
                           => n_3618);
   clk_r_REG10523_S1 : DFF_X1 port map( D => n36784, CK => CLK, Q => n40714, QN
                           => n_3619);
   clk_r_REG11803_S1 : DFF_X1 port map( D => n36137, CK => CLK, Q => n40713, QN
                           => n_3620);
   clk_r_REG13319_S1 : DFF_X1 port map( D => n36534, CK => CLK, Q => n40712, QN
                           => n_3621);
   clk_r_REG11394_S1 : DFF_X1 port map( D => n36138, CK => CLK, Q => n40711, QN
                           => n_3622);
   clk_r_REG10898_S1 : DFF_X1 port map( D => n36139, CK => CLK, Q => n40710, QN
                           => n_3623);
   clk_r_REG11432_S1 : DFF_X1 port map( D => n35869, CK => CLK, Q => n40709, QN
                           => n_3624);
   clk_r_REG12293_S1 : DFF_X1 port map( D => n35868, CK => CLK, Q => n40708, QN
                           => n_3625);
   clk_r_REG11823_S1 : DFF_X1 port map( D => n35867, CK => CLK, Q => n40707, QN
                           => n_3626);
   clk_r_REG12140_S1 : DFF_X1 port map( D => n36523, CK => CLK, Q => n40706, QN
                           => n_3627);
   clk_r_REG12102_S1 : DFF_X1 port map( D => n35866, CK => CLK, Q => n40705, QN
                           => n_3628);
   clk_r_REG12844_S1 : DFF_X1 port map( D => n36521, CK => CLK, Q => n40704, QN
                           => n_3629);
   clk_r_REG11973_S1 : DFF_X1 port map( D => n35865, CK => CLK, Q => n40703, QN
                           => n_3630);
   clk_r_REG13138_S1 : DFF_X1 port map( D => n35864, CK => CLK, Q => n40702, QN
                           => n_3631);
   clk_r_REG12060_S1 : DFF_X1 port map( D => n35863, CK => CLK, Q => n40701, QN
                           => n_3632);
   clk_r_REG13337_S1 : DFF_X1 port map( D => n35862, CK => CLK, Q => n40700, QN
                           => n_3633);
   clk_r_REG12295_S1 : DFF_X1 port map( D => n35861, CK => CLK, Q => n40699, QN
                           => n_3634);
   clk_r_REG13140_S1 : DFF_X1 port map( D => n35860, CK => CLK, Q => n40698, QN
                           => n_3635);
   clk_r_REG13186_S1 : DFF_X1 port map( D => n35859, CK => CLK, Q => n40697, QN
                           => n_3636);
   clk_r_REG12062_S1 : DFF_X1 port map( D => n35858, CK => CLK, Q => n40696, QN
                           => n_3637);
   clk_r_REG13142_S1 : DFF_X1 port map( D => n35857, CK => CLK, Q => n40695, QN
                           => n_3638);
   clk_r_REG13174_S1 : DFF_X1 port map( D => n36023, CK => CLK, Q => n40694, QN
                           => n_3639);
   clk_r_REG13032_S1 : DFF_X1 port map( D => n36744, CK => CLK, Q => n40693, QN
                           => n_3640);
   clk_r_REG11975_S1 : DFF_X1 port map( D => n35856, CK => CLK, Q => n40692, QN
                           => n_3641);
   clk_r_REG12104_S1 : DFF_X1 port map( D => n35855, CK => CLK, Q => n40691, QN
                           => n_3642);
   clk_r_REG12170_S1 : DFF_X1 port map( D => n35854, CK => CLK, Q => n40690, QN
                           => n_3643);
   clk_r_REG11434_S1 : DFF_X1 port map( D => n35852, CK => CLK, Q => n40689, QN
                           => n_3644);
   clk_r_REG10922_S1 : DFF_X1 port map( D => n35851, CK => CLK, Q => n40688, QN
                           => n_3645);
   clk_r_REG12471_S1 : DFF_X1 port map( D => n36745, CK => CLK, Q => n40687, QN
                           => n_3646);
   clk_r_REG12627_S1 : DFF_X1 port map( D => n36746, CK => CLK, Q => n40686, QN
                           => n_3647);
   clk_r_REG12866_S1 : DFF_X1 port map( D => n36140, CK => CLK, Q => n40685, QN
                           => n_3648);
   clk_r_REG10636_S1 : DFF_X1 port map( D => n36749, CK => CLK, Q => n40684, QN
                           => n_3649);
   clk_r_REG13333_S1 : DFF_X1 port map( D => n36141, CK => CLK, Q => n40683, QN
                           => n_3650);
   clk_r_REG13062_S1 : DFF_X1 port map( D => n36537, CK => CLK, Q => n40682, QN
                           => n_3651);
   clk_r_REG12511_S1 : DFF_X1 port map( D => n36533, CK => CLK, Q => n40681, QN
                           => n_3652);
   clk_r_REG12281_S1 : DFF_X1 port map( D => n36142, CK => CLK, Q => n40680, QN
                           => n_3653);
   clk_r_REG12639_S1 : DFF_X1 port map( D => n36531, CK => CLK, Q => n40679, QN
                           => n_3654);
   clk_r_REG13106_S1 : DFF_X1 port map( D => n36143, CK => CLK, Q => n40678, QN
                           => n_3655);
   clk_r_REG12026_S1 : DFF_X1 port map( D => n36144, CK => CLK, Q => n40677, QN
                           => n_3656);
   clk_r_REG12974_S1 : DFF_X1 port map( D => n36754, CK => CLK, Q => n40676, QN
                           => n_3657);
   clk_r_REG12469_S1 : DFF_X1 port map( D => n36757, CK => CLK, Q => n40675, QN
                           => n_3658);
   clk_r_REG12589_S1 : DFF_X1 port map( D => n36759, CK => CLK, Q => n40674, QN
                           => n_3659);
   clk_r_REG13006_S1 : DFF_X1 port map( D => n36762, CK => CLK, Q => n40673, QN
                           => n_3660);
   clk_r_REG13018_S1 : DFF_X1 port map( D => n36524, CK => CLK, Q => n40672, QN
                           => n_3661);
   clk_r_REG13004_S1 : DFF_X1 port map( D => n36767, CK => CLK, Q => n40671, QN
                           => n_3662);
   clk_r_REG12972_S1 : DFF_X1 port map( D => n36768, CK => CLK, Q => n40670, QN
                           => n_3663);
   clk_r_REG13028_S1 : DFF_X1 port map( D => n36772, CK => CLK, Q => n40669, QN
                           => n_3664);
   clk_r_REG13026_S1 : DFF_X1 port map( D => n36773, CK => CLK, Q => n40668, QN
                           => n_3665);
   clk_r_REG12463_S1 : DFF_X1 port map( D => n36774, CK => CLK, Q => n40667, QN
                           => n_3666);
   clk_r_REG12597_S1 : DFF_X1 port map( D => n36704, CK => CLK, Q => n40666, QN
                           => n_3667);
   clk_r_REG12970_S1 : DFF_X1 port map( D => n36777, CK => CLK, Q => n40665, QN
                           => n_3668);
   clk_r_REG12968_S1 : DFF_X1 port map( D => n36780, CK => CLK, Q => n40664, QN
                           => n_3669);
   clk_r_REG12964_S1 : DFF_X1 port map( D => n36838, CK => CLK, Q => n40663, QN
                           => n_3670);
   clk_r_REG13468_S4 : DFFS_X1 port map( D => n47493, CK => CLK, SN => 
                           RESET_BAR, Q => n40662, QN => n_3671);
   clk_r_REG13466_S3 : DFFR_X1 port map( D => n47505, CK => CLK, RN => 
                           RESET_BAR, Q => n_3672, QN => n47493);
   clk_r_REG13467_S4 : DFFS_X1 port map( D => n47493, CK => CLK, SN => 
                           RESET_BAR, Q => n_3673, QN => n40660);
   clk_r_REG13470_S3 : DFFR_X1 port map( D => n47504, CK => CLK, RN => 
                           RESET_BAR, Q => n_3674, QN => n47494);
   clk_r_REG13471_S4 : DFFS_X1 port map( D => n47494, CK => CLK, SN => 
                           RESET_BAR, Q => n_3675, QN => n40658);
   clk_r_REG13621_S7 : DFFR_X1 port map( D => ADD_RD2(3), CK => CLK, RN => 
                           RESET_BAR, Q => n40657, QN => n_3676);
   clk_r_REG13519_S7 : DFFR_X1 port map( D => ADD_RD1(3), CK => CLK, RN => 
                           RESET_BAR, Q => n40656, QN => n_3677);
   clk_r_REG13595_S7 : DFFS_X1 port map( D => n47498, CK => CLK, SN => 
                           RESET_BAR, Q => n47432, QN => n49081);
   clk_r_REG13583_S7 : DFFS_X1 port map( D => n47503, CK => CLK, SN => 
                           RESET_BAR, Q => n_3678, QN => n49077);
   clk_r_REG13580_S7 : DFFS_X1 port map( D => n47497, CK => CLK, SN => n47506, 
                           Q => n_3679, QN => n49079);
   clk_r_REG13592_S7 : DFFS_X1 port map( D => n47502, CK => CLK, SN => n47506, 
                           Q => n47449, QN => n49080);
   clk_r_REG13456_S2 : DFFR_X1 port map( D => n30121, CK => CLK, RN => 
                           RESET_BAR, Q => n40645, QN => n_3680);
   clk_r_REG13457_S3 : DFFR_X1 port map( D => n40645, CK => CLK, RN => 
                           RESET_BAR, Q => n40644, QN => n_3681);
   clk_r_REG13458_S4 : DFFR_X1 port map( D => n40644, CK => CLK, RN => 
                           RESET_BAR, Q => n40643, QN => n_3682);
   clk_r_REG13453_S2 : DFFR_X1 port map( D => n30118, CK => CLK, RN => 
                           RESET_BAR, Q => n40641, QN => n_3683);
   clk_r_REG13454_S3 : DFFR_X1 port map( D => n40641, CK => CLK, RN => 
                           RESET_BAR, Q => n40640, QN => n_3684);
   clk_r_REG13455_S4 : DFFR_X1 port map( D => n40640, CK => CLK, RN => 
                           RESET_BAR, Q => n40639, QN => n_3685);
   clk_r_REG13444_S2 : DFFR_X1 port map( D => n30113, CK => CLK, RN => 
                           RESET_BAR, Q => n40635, QN => n_3686);
   clk_r_REG13445_S3 : DFFR_X1 port map( D => n40635, CK => CLK, RN => n47506, 
                           Q => n40634, QN => n_3687);
   clk_r_REG13446_S4 : DFFR_X1 port map( D => n40634, CK => CLK, RN => 
                           RESET_BAR, Q => n40633, QN => n_3688);
   clk_r_REG13441_S2 : DFFR_X1 port map( D => n30110, CK => CLK, RN => 
                           RESET_BAR, Q => n40631, QN => n_3689);
   clk_r_REG13442_S3 : DFFR_X1 port map( D => n40631, CK => CLK, RN => 
                           RESET_BAR, Q => n40630, QN => n_3690);
   clk_r_REG13443_S4 : DFFR_X1 port map( D => n40630, CK => CLK, RN => 
                           RESET_BAR, Q => n40629, QN => n_3691);
   clk_r_REG13588_S7 : DFFR_X1 port map( D => n30083, CK => CLK, RN => 
                           RESET_BAR, Q => n49092, QN => n_3692);
   clk_r_REG13578_S7 : DFFR_X1 port map( D => n30082, CK => CLK, RN => 
                           RESET_BAR, Q => n49093, QN => n_3693);
   clk_r_REG13585_S7 : DFFR_X1 port map( D => n30081, CK => CLK, RN => 
                           RESET_BAR, Q => n49094, QN => n_3694);
   clk_r_REG13577_S7 : DFFR_X1 port map( D => n30080, CK => CLK, RN => 
                           RESET_BAR, Q => n49087, QN => n_3695);
   clk_r_REG13594_S7 : DFFR_X1 port map( D => n30079, CK => CLK, RN => 
                           RESET_BAR, Q => n49089, QN => n_3696);
   clk_r_REG13597_S7 : DFFR_X1 port map( D => n30078, CK => CLK, RN => 
                           RESET_BAR, Q => n49091, QN => n_3697);
   clk_r_REG13584_S7 : DFFR_X1 port map( D => n30077, CK => CLK, RN => 
                           RESET_BAR, Q => n49090, QN => n_3698);
   clk_r_REG13600_S7 : DFFR_X1 port map( D => n30076, CK => CLK, RN => 
                           RESET_BAR, Q => n49086, QN => n_3699);
   clk_r_REG13590_S7 : DFFR_X1 port map( D => n30075, CK => CLK, RN => 
                           RESET_BAR, Q => n49088, QN => n_3700);
   clk_r_REG13593_S7 : DFFR_X1 port map( D => n30071, CK => CLK, RN => 
                           RESET_BAR, Q => n49085, QN => n_3701);
   clk_r_REG13513_S7 : DFFR_X1 port map( D => n30060, CK => CLK, RN => 
                           RESET_BAR, Q => n49095, QN => n_3702);
   clk_r_REG13500_S7 : DFFR_X1 port map( D => n30056, CK => CLK, RN => 
                           RESET_BAR, Q => n49096, QN => n_3703);
   clk_r_REG13509_S7 : DFFR_X1 port map( D => n30054, CK => CLK, RN => 
                           RESET_BAR, Q => n49097, QN => n_3704);
   clk_r_REG13598_S7 : DFFR_X1 port map( D => n47500, CK => CLK, RN => 
                           RESET_BAR, Q => n_3705, QN => n49076);
   clk_r_REG13604_S7 : DFFS_X1 port map( D => n47499, CK => CLK, SN => 
                           RESET_BAR, Q => n47447, QN => n49083);
   clk_r_REG13607_S7 : DFFS_X1 port map( D => n47501, CK => CLK, SN => 
                           RESET_BAR, Q => n47446, QN => n49084);
   clk_r_REG13589_S7 : DFFS_X1 port map( D => n47495, CK => CLK, SN => 
                           RESET_BAR, Q => n47453, QN => n49082);
   clk_r_REG13586_S7 : DFFS_X1 port map( D => n47496, CK => CLK, SN => 
                           RESET_BAR, Q => n_3706, QN => n49078);
   clk_r_REG13462_S2 : DFFS_X1 port map( D => n30048, CK => CLK, SN => 
                           RESET_BAR, Q => n40563, QN => n_3707);
   clk_r_REG13463_S3 : DFFS_X1 port map( D => n40563, CK => CLK, SN => 
                           RESET_BAR, Q => n40562, QN => n_3708);
   clk_r_REG13464_S4 : DFFS_X1 port map( D => n40562, CK => CLK, SN => 
                           RESET_BAR, Q => n40561, QN => n_3709);
   clk_r_REG13459_S2 : DFFR_X1 port map( D => n30046, CK => CLK, RN => 
                           RESET_BAR, Q => n40560, QN => n_3710);
   clk_r_REG13460_S3 : DFFR_X1 port map( D => n40560, CK => CLK, RN => 
                           RESET_BAR, Q => n40559, QN => n_3711);
   clk_r_REG13461_S4 : DFFR_X1 port map( D => n40559, CK => CLK, RN => 
                           RESET_BAR, Q => n40558, QN => n_3712);
   clk_r_REG13450_S2 : DFFR_X1 port map( D => n30044, CK => CLK, RN => 
                           RESET_BAR, Q => n40557, QN => n_3713);
   clk_r_REG13451_S3 : DFFR_X1 port map( D => n40557, CK => CLK, RN => 
                           RESET_BAR, Q => n40556, QN => n_3714);
   clk_r_REG13452_S4 : DFFR_X1 port map( D => n40556, CK => CLK, RN => 
                           RESET_BAR, Q => n40555, QN => n_3715);
   clk_r_REG13447_S2 : DFFR_X1 port map( D => n30042, CK => CLK, RN => 
                           RESET_BAR, Q => n40554, QN => n_3716);
   clk_r_REG13448_S3 : DFFR_X1 port map( D => n40554, CK => CLK, RN => 
                           RESET_BAR, Q => n40553, QN => n_3717);
   clk_r_REG13449_S4 : DFFR_X1 port map( D => n40553, CK => CLK, RN => 
                           RESET_BAR, Q => n40552, QN => n_3718);
   clk_r_REG13501_S7 : DFFR_X1 port map( D => n30058, CK => CLK, RN => 
                           RESET_BAR, Q => n40577, QN => n_3719);
   clk_r_REG13502_S7 : DFFR_X1 port map( D => n30061, CK => CLK, RN => 
                           RESET_BAR, Q => n40580, QN => n_3720);
   clk_r_REG13512_S7 : DFFR_X1 port map( D => n30059, CK => CLK, RN => 
                           RESET_BAR, Q => n47430, QN => n_3721);
   clk_r_REG13505_S7 : DFFR_X1 port map( D => n30064, CK => CLK, RN => 
                           RESET_BAR, Q => n40583, QN => n_3722);
   clk_r_REG13515_S7 : DFFR_X1 port map( D => n30068, CK => CLK, RN => 
                           RESET_BAR, Q => n40587, QN => n_3723);
   clk_r_REG13582_S7 : DFFR_X1 port map( D => n30073, CK => CLK, RN => 
                           RESET_BAR, Q => n40592, QN => n_3724);
   clk_r_REG13581_S7 : DFFR_X1 port map( D => n30072, CK => CLK, RN => 
                           RESET_BAR, Q => n40591, QN => n_3725);
   clk_r_REG13596_S7 : DFFR_X1 port map( D => n30069, CK => CLK, RN => 
                           RESET_BAR, Q => n40588, QN => n_3726);
   clk_r_REG13599_S7 : DFFR_X1 port map( D => n30074, CK => CLK, RN => 
                           RESET_BAR, Q => n47428, QN => n_3727);
   clk_r_REG13612_S7 : DFFS_X1 port map( D => n1530, CK => CLK, SN => RESET_BAR
                           , Q => n_3728, QN => n40655);
   clk_r_REG13576_S7 : DFFS_X1 port map( D => n1533, CK => CLK, SN => n47506, Q
                           => n_3729, QN => n40565);
   clk_r_REG13605_S7 : DFFS_X1 port map( D => n1528, CK => CLK, SN => n47506, Q
                           => n_3730, QN => n40648);
   clk_r_REG13504_S7 : DFFR_X1 port map( D => n30063, CK => CLK, RN => 
                           RESET_BAR, Q => n40582, QN => n_3731);
   clk_r_REG13514_S7 : DFFR_X1 port map( D => n30065, CK => CLK, RN => 
                           RESET_BAR, Q => n40584, QN => n_3732);
   clk_r_REG13510_S7 : DFFR_X1 port map( D => n30055, CK => CLK, RN => 
                           RESET_BAR, Q => n40574, QN => n_3733);
   clk_r_REG13508_S7 : DFFR_X1 port map( D => n30053, CK => CLK, RN => 
                           RESET_BAR, Q => n47431, QN => n_3734);
   clk_r_REG13503_S7 : DFFR_X1 port map( D => n30062, CK => CLK, RN => 
                           RESET_BAR, Q => n40581, QN => n_3735);
   clk_r_REG13587_S7 : DFFR_X1 port map( D => n30070, CK => CLK, RN => 
                           RESET_BAR, Q => n40589, QN => n_3736);
   clk_r_REG13591_S7 : DFFR_X1 port map( D => n30084, CK => CLK, RN => 
                           RESET_BAR, Q => n47429, QN => n_3737);
   clk_r_REG13614_S7 : DFFR_X1 port map( D => n1529, CK => CLK, RN => RESET_BAR
                           , Q => n_3738, QN => n40571);
   clk_r_REG13610_S7 : DFFS_X1 port map( D => n1531, CK => CLK, SN => RESET_BAR
                           , Q => n_3739, QN => n40654);
   clk_r_REG13602_S7 : DFFS_X1 port map( D => n1527, CK => CLK, SN => n47506, Q
                           => n_3740, QN => n40649);
   clk_r_REG13507_S7 : DFFR_X1 port map( D => n30067, CK => CLK, RN => 
                           RESET_BAR, Q => n40586, QN => n_3741);
   clk_r_REG13511_S7 : DFFR_X1 port map( D => n30057, CK => CLK, RN => 
                           RESET_BAR, Q => n40576, QN => n_3742);
   clk_r_REG13506_S7 : DFFR_X1 port map( D => n30066, CK => CLK, RN => 
                           RESET_BAR, Q => n40585, QN => n_3743);
   clk_r_REG13608_S7 : DFFS_X1 port map( D => n1532, CK => CLK, SN => n47506, Q
                           => n_3744, QN => n40568);
   clk_r_REG13615_S7 : DFFS_X1 port map( D => n31166, CK => CLK, SN => n47506, 
                           Q => n41690, QN => n_3745);
   clk_r_REG13611_S7 : DFFR_X1 port map( D => n31169, CK => CLK, RN => 
                           RESET_BAR, Q => n41688, QN => n_3746);
   clk_r_REG13603_S7 : DFFR_X1 port map( D => n31167, CK => CLK, RN => 
                           RESET_BAR, Q => n41687, QN => n_3747);
   clk_r_REG13606_S7 : DFFR_X1 port map( D => n31171, CK => CLK, RN => 
                           RESET_BAR, Q => n41689, QN => n_3748);
   clk_r_REG13609_S7 : DFFR_X1 port map( D => n31170, CK => CLK, RN => 
                           RESET_BAR, Q => n41686, QN => n_3749);
   clk_r_REG13397_S2 : DFFS_X2 port map( D => n30094, CK => CLK, SN => 
                           RESET_BAR, Q => n40613, QN => n_3750);
   clk_r_REG13399_S2 : DFFS_X2 port map( D => n30096, CK => CLK, SN => n47506, 
                           Q => n40615, QN => n_3751);
   clk_r_REG13400_S2 : DFFS_X2 port map( D => n30097, CK => CLK, SN => 
                           RESET_BAR, Q => n40616, QN => n_3752);
   clk_r_REG13401_S2 : DFFS_X2 port map( D => n30098, CK => CLK, SN => 
                           RESET_BAR, Q => n40617, QN => n_3753);
   clk_r_REG13402_S2 : DFFS_X2 port map( D => n30099, CK => CLK, SN => 
                           RESET_BAR, Q => n40618, QN => n_3754);
   clk_r_REG13388_S2 : DFFS_X2 port map( D => n30101, CK => CLK, SN => n47506, 
                           Q => n40620, QN => n_3755);
   clk_r_REG13390_S2 : DFFS_X2 port map( D => n30103, CK => CLK, SN => 
                           RESET_BAR, Q => n40622, QN => n_3756);
   clk_r_REG13392_S2 : DFFS_X2 port map( D => n30105, CK => CLK, SN => 
                           RESET_BAR, Q => n40624, QN => n_3757);
   clk_r_REG13411_S2 : DFFS_X2 port map( D => n30124, CK => CLK, SN => n47506, 
                           Q => n40647, QN => n_3758);
   clk_r_REG13396_S2 : DFFS_X2 port map( D => n30093, CK => CLK, SN => n47506, 
                           Q => n40612, QN => n_3759);
   clk_r_REG13409_S2 : DFFS_X2 port map( D => n30120, CK => CLK, SN => 
                           RESET_BAR, Q => n40642, QN => n_3760);
   clk_r_REG13407_S2 : DFFS_X2 port map( D => n30116, CK => CLK, SN => 
                           RESET_BAR, Q => n40637, QN => n_3761);
   clk_r_REG13408_S2 : DFFS_X2 port map( D => n30117, CK => CLK, SN => 
                           RESET_BAR, Q => n40638, QN => n_3762);
   clk_r_REG13405_S2 : DFFS_X2 port map( D => n30112, CK => CLK, SN => 
                           RESET_BAR, Q => n40632, QN => n_3763);
   clk_r_REG13406_S2 : DFFS_X2 port map( D => n30115, CK => CLK, SN => 
                           RESET_BAR, Q => n40636, QN => n_3764);
   clk_r_REG13395_S2 : DFFS_X2 port map( D => n30108, CK => CLK, SN => n47506, 
                           Q => n40627, QN => n_3765);
   clk_r_REG13404_S2 : DFFS_X2 port map( D => n30109, CK => CLK, SN => 
                           RESET_BAR, Q => n40628, QN => n_3766);
   clk_r_REG13393_S2 : DFFS_X2 port map( D => n30106, CK => CLK, SN => n47506, 
                           Q => n40625, QN => n_3767);
   clk_r_REG13394_S2 : DFFS_X2 port map( D => n30107, CK => CLK, SN => n47506, 
                           Q => n40626, QN => n_3768);
   clk_r_REG13389_S2 : DFFS_X2 port map( D => n30102, CK => CLK, SN => n47506, 
                           Q => n40621, QN => n_3769);
   clk_r_REG13391_S2 : DFFS_X2 port map( D => n30104, CK => CLK, SN => 
                           RESET_BAR, Q => n40623, QN => n_3770);
   clk_r_REG13398_S2 : DFFS_X2 port map( D => n30095, CK => CLK, SN => n47506, 
                           Q => n40614, QN => n_3771);
   clk_r_REG13403_S2 : DFFS_X2 port map( D => n30100, CK => CLK, SN => n47506, 
                           Q => n40619, QN => n_3772);
   clk_r_REG13386_S2 : DFFS_X2 port map( D => n30091, CK => CLK, SN => n47506, 
                           Q => n40610, QN => n_3773);
   clk_r_REG13387_S2 : DFFS_X2 port map( D => n30092, CK => CLK, SN => n47506, 
                           Q => n40611, QN => n_3774);
   clk_r_REG13384_S2 : DFFS_X2 port map( D => n30089, CK => CLK, SN => n47506, 
                           Q => n40608, QN => n_3775);
   clk_r_REG13385_S2 : DFFS_X2 port map( D => n30090, CK => CLK, SN => 
                           RESET_BAR, Q => n40609, QN => n_3776);
   clk_r_REG13382_S2 : DFFS_X2 port map( D => n30087, CK => CLK, SN => n47506, 
                           Q => n40606, QN => n_3777);
   clk_r_REG13383_S2 : DFFS_X2 port map( D => n30088, CK => CLK, SN => 
                           RESET_BAR, Q => n40607, QN => n_3778);
   clk_r_REG13380_S2 : DFFS_X2 port map( D => n30085, CK => CLK, SN => 
                           RESET_BAR, Q => n40604, QN => n_3779);
   clk_r_REG13381_S2 : DFFS_X2 port map( D => n30086, CK => CLK, SN => 
                           RESET_BAR, Q => n40605, QN => n_3780);
   clk_r_REG13410_S2 : DFFS_X2 port map( D => n30123, CK => CLK, SN => 
                           RESET_BAR, Q => n40646, QN => n_3781);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n47506);
   U4 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40646, ZN => n47562);
   U5 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40604, ZN => n47566);
   U6 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40605, ZN => n47565);
   U7 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40606, ZN => n47551);
   U8 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40607, ZN => n47550);
   U9 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40608, ZN => n47548);
   U10 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40609, ZN => n47544);
   U11 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40610, ZN => n47540);
   U12 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40611, ZN => n47543);
   U13 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40620, ZN => n47558);
   U14 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40621, ZN => n47539);
   U15 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40622, ZN => n47546);
   U16 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40623, ZN => n47535);
   U17 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40624, ZN => n47556);
   U18 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40625, ZN => n47552);
   U19 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40626, ZN => n47553);
   U20 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40627, ZN => n47554);
   U21 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40612, ZN => n47559);
   U22 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40613, ZN => n47532);
   U23 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40614, ZN => n47536);
   U24 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40615, ZN => n47545);
   U25 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40616, ZN => n47560);
   U26 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40617, ZN => n47538);
   U27 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40618, ZN => n47557);
   U28 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40619, ZN => n47541);
   U29 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40628, ZN => n47512);
   U30 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40632, ZN => n47547);
   U31 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40636, ZN => n47542);
   U32 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40637, ZN => n47511);
   U33 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40638, ZN => n47563);
   U34 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40642, ZN => n47561);
   U35 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n40647, ZN => n47567);
   U36 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n42749, ZN => n47570);
   U37 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n42742, ZN => n47549);
   U38 : NAND3_X1 port map( A1 => n47506, A2 => n42760, A3 => n42757, ZN => 
                           n48334);
   U39 : CLKBUF_X1 port map( A => n48334, Z => n48133);
   U40 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n42760, A3 => n42758, ZN => 
                           n49075);
   U41 : CLKBUF_X1 port map( A => n49075, Z => n49012);
   U42 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), A3 => ADD_RD1(0)
                           , ZN => n31166);
   U43 : INV_X1 port map( A => n31166, ZN => n1529);
   U44 : NAND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n47507);
   U45 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n47507, ZN => n31171);
   U46 : INV_X1 port map( A => n31171, ZN => n1528);
   U47 : INV_X1 port map( A => ADD_RD1(2), ZN => n47509);
   U48 : NOR2_X1 port map( A1 => n47509, A2 => n47507, ZN => n31169);
   U49 : INV_X1 port map( A => n31169, ZN => n1531);
   U50 : INV_X1 port map( A => ADD_RD1(1), ZN => n47508);
   U51 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => n47508, ZN
                           => n31170);
   U52 : INV_X1 port map( A => n31170, ZN => n1532);
   U53 : OR3_X1 port map( A1 => n47508, A2 => n47509, A3 => ADD_RD1(0), ZN => 
                           n47501);
   U54 : INV_X1 port map( A => ADD_RD2(2), ZN => n47588);
   U55 : INV_X1 port map( A => ADD_RD2(1), ZN => n47590);
   U56 : OR3_X1 port map( A1 => n47588, A2 => n47590, A3 => ADD_RD2(0), ZN => 
                           n47496);
   U57 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n47508, ZN => n47510);
   U58 : NOR2_X1 port map( A1 => n47509, A2 => n47510, ZN => n31164);
   U59 : INV_X1 port map( A => n31164, ZN => n1530);
   U60 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n47510, ZN => n31167);
   U61 : INV_X1 port map( A => n31167, ZN => n1527);
   U62 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => n47590, ZN
                           => n31168);
   U63 : INV_X1 port map( A => n31168, ZN => n1533);
   U64 : INV_X1 port map( A => ADD_WR(3), ZN => n1526);
   U65 : INV_X1 port map( A => ADD_WR(4), ZN => n1525);
   U66 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42737, ZN => n47528);
   U67 : OAI22_X1 port map( A1 => n40632, A2 => n47528, B1 => n42720, B2 => 
                           n47547, ZN => n35769);
   U68 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42724, ZN => n47519);
   U69 : OAI22_X1 port map( A1 => n40606, A2 => n47519, B1 => n42719, B2 => 
                           n47551, ZN => n35770);
   U70 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42729, ZN => n47514);
   U71 : OAI22_X1 port map( A1 => n40606, A2 => n47514, B1 => n42718, B2 => 
                           n47551, ZN => n35771);
   U72 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42725, ZN => n47517);
   U73 : OAI22_X1 port map( A1 => n40606, A2 => n47517, B1 => n42717, B2 => 
                           n47551, ZN => n35772);
   U74 : OAI22_X1 port map( A1 => n40607, A2 => n47519, B1 => n42716, B2 => 
                           n47550, ZN => n35773);
   U75 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42734, ZN => n47524);
   U76 : OAI22_X1 port map( A1 => n40632, A2 => n47524, B1 => n42715, B2 => 
                           n47547, ZN => n35774);
   U77 : OAI22_X1 port map( A1 => n40609, A2 => n47519, B1 => n42714, B2 => 
                           n47544, ZN => n35775);
   U78 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42727, ZN => n47515);
   U79 : OAI22_X1 port map( A1 => n40607, A2 => n47515, B1 => n42713, B2 => 
                           n47550, ZN => n35776);
   U80 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42728, ZN => n47518);
   U81 : OAI22_X1 port map( A1 => n40607, A2 => n47518, B1 => n42712, B2 => 
                           n47550, ZN => n35777);
   U82 : OAI22_X1 port map( A1 => n40608, A2 => n47515, B1 => n42711, B2 => 
                           n47548, ZN => n35778);
   U83 : OAI22_X1 port map( A1 => n40606, A2 => n47518, B1 => n42710, B2 => 
                           n47551, ZN => n35779);
   U84 : OAI22_X1 port map( A1 => n40608, A2 => n47517, B1 => n42709, B2 => 
                           n47548, ZN => n35780);
   U85 : OAI22_X1 port map( A1 => n40609, A2 => n47515, B1 => n42708, B2 => 
                           n47544, ZN => n35781);
   U86 : OAI22_X1 port map( A1 => n40606, A2 => n47515, B1 => n42707, B2 => 
                           n47551, ZN => n35782);
   U87 : OAI22_X1 port map( A1 => n40609, A2 => n47514, B1 => n42706, B2 => 
                           n47544, ZN => n35783);
   U88 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42726, ZN => n47516);
   U89 : OAI22_X1 port map( A1 => n40608, A2 => n47516, B1 => n42705, B2 => 
                           n47548, ZN => n35784);
   U90 : OAI22_X1 port map( A1 => n40632, A2 => n47549, B1 => n42704, B2 => 
                           n47547, ZN => n35785);
   U91 : OAI22_X1 port map( A1 => n40608, A2 => n47514, B1 => n42703, B2 => 
                           n47548, ZN => n35786);
   U92 : OAI22_X1 port map( A1 => n40609, A2 => n47517, B1 => n42702, B2 => 
                           n47544, ZN => n35787);
   U93 : OAI22_X1 port map( A1 => n40609, A2 => n47516, B1 => n42701, B2 => 
                           n47544, ZN => n35788);
   U94 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42723, ZN => n47537);
   U95 : OAI22_X1 port map( A1 => n40609, A2 => n47537, B1 => n42700, B2 => 
                           n47544, ZN => n35789);
   U96 : OAI22_X1 port map( A1 => n40608, A2 => n47518, B1 => n42699, B2 => 
                           n47548, ZN => n35790);
   U97 : OAI22_X1 port map( A1 => n40608, A2 => n47519, B1 => n42698, B2 => 
                           n47548, ZN => n35791);
   U98 : OAI22_X1 port map( A1 => n40607, A2 => n47516, B1 => n42697, B2 => 
                           n47550, ZN => n35792);
   U99 : OAI22_X1 port map( A1 => n40607, A2 => n47517, B1 => n42696, B2 => 
                           n47550, ZN => n35793);
   U100 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42741, ZN => n47530);
   U101 : OAI22_X1 port map( A1 => n40632, A2 => n47530, B1 => n42695, B2 => 
                           n47547, ZN => n35794);
   U102 : OAI22_X1 port map( A1 => n40608, A2 => n47537, B1 => n42694, B2 => 
                           n47548, ZN => n35795);
   U103 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42733, ZN => n47555);
   U104 : OAI22_X1 port map( A1 => n40606, A2 => n47555, B1 => n42693, B2 => 
                           n47551, ZN => n35796);
   U105 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42732, ZN => n47533);
   U106 : OAI22_X1 port map( A1 => n40627, A2 => n47533, B1 => n42692, B2 => 
                           n47554, ZN => n35797);
   U107 : OAI22_X1 port map( A1 => n40625, A2 => n47555, B1 => n42691, B2 => 
                           n47552, ZN => n35798);
   U108 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42736, ZN => n47520);
   U109 : OAI22_X1 port map( A1 => n40625, A2 => n47520, B1 => n42690, B2 => 
                           n47552, ZN => n35799);
   U110 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42731, ZN => n47527);
   U111 : OAI22_X1 port map( A1 => n40625, A2 => n47527, B1 => n42689, B2 => 
                           n47552, ZN => n35800);
   U112 : OAI22_X1 port map( A1 => n40626, A2 => n47524, B1 => n42688, B2 => 
                           n47553, ZN => n35801);
   U113 : OAI22_X1 port map( A1 => n40632, A2 => n47518, B1 => n42687, B2 => 
                           n47547, ZN => n35802);
   U114 : OAI22_X1 port map( A1 => n40626, A2 => n47520, B1 => n42686, B2 => 
                           n47553, ZN => n35803);
   U115 : OAI22_X1 port map( A1 => n40625, A2 => n47524, B1 => n42685, B2 => 
                           n47552, ZN => n35804);
   U116 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42735, ZN => n47531);
   U117 : OAI22_X1 port map( A1 => n40625, A2 => n47531, B1 => n42684, B2 => 
                           n47552, ZN => n35805);
   U118 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42744, ZN => n47526);
   U119 : OAI22_X1 port map( A1 => n40627, A2 => n47526, B1 => n42683, B2 => 
                           n47554, ZN => n35806);
   U120 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42739, ZN => n47522);
   U121 : OAI22_X1 port map( A1 => n40627, A2 => n47522, B1 => n42682, B2 => 
                           n47554, ZN => n35807);
   U122 : OAI22_X1 port map( A1 => n40625, A2 => n47528, B1 => n42681, B2 => 
                           n47552, ZN => n35808);
   U123 : OAI22_X1 port map( A1 => n40632, A2 => n47520, B1 => n42680, B2 => 
                           n47547, ZN => n35809);
   U124 : OAI22_X1 port map( A1 => n40627, A2 => n47520, B1 => n42679, B2 => 
                           n47554, ZN => n35810);
   U125 : OAI22_X1 port map( A1 => n40627, A2 => n47549, B1 => n42678, B2 => 
                           n47554, ZN => n35811);
   U126 : OAI22_X1 port map( A1 => n40625, A2 => n47530, B1 => n42677, B2 => 
                           n47552, ZN => n35812);
   U127 : OAI22_X1 port map( A1 => n40625, A2 => n47549, B1 => n42676, B2 => 
                           n47552, ZN => n35813);
   U128 : OAI22_X1 port map( A1 => n40632, A2 => n47514, B1 => n42675, B2 => 
                           n47547, ZN => n35814);
   U129 : OAI22_X1 port map( A1 => n40609, A2 => n47518, B1 => n42674, B2 => 
                           n47544, ZN => n35815);
   U130 : OAI22_X1 port map( A1 => n40626, A2 => n47549, B1 => n42673, B2 => 
                           n47553, ZN => n35816);
   U131 : OAI22_X1 port map( A1 => n40627, A2 => n47524, B1 => n42672, B2 => 
                           n47554, ZN => n35817);
   U132 : OAI22_X1 port map( A1 => n40606, A2 => n47516, B1 => n42671, B2 => 
                           n47551, ZN => n35818);
   U133 : OAI22_X1 port map( A1 => n40626, A2 => n47522, B1 => n42670, B2 => 
                           n47553, ZN => n35819);
   U134 : OAI22_X1 port map( A1 => n40607, A2 => n47514, B1 => n42669, B2 => 
                           n47550, ZN => n35820);
   U135 : OAI22_X1 port map( A1 => n40632, A2 => n47537, B1 => n42668, B2 => 
                           n47547, ZN => n35821);
   U136 : OAI22_X1 port map( A1 => n40608, A2 => n47527, B1 => n42667, B2 => 
                           n47548, ZN => n35822);
   U137 : OAI22_X1 port map( A1 => n40607, A2 => n47526, B1 => n42666, B2 => 
                           n47550, ZN => n35823);
   U138 : OAI22_X1 port map( A1 => n40607, A2 => n47549, B1 => n42665, B2 => 
                           n47550, ZN => n35824);
   U139 : OAI22_X1 port map( A1 => n40607, A2 => n47530, B1 => n42664, B2 => 
                           n47550, ZN => n35825);
   U140 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42740, ZN => n47523);
   U141 : OAI22_X1 port map( A1 => n40632, A2 => n47523, B1 => n42663, B2 => 
                           n47547, ZN => n35826);
   U142 : OAI22_X1 port map( A1 => n40606, A2 => n47527, B1 => n42662, B2 => 
                           n47551, ZN => n35827);
   U143 : OAI22_X1 port map( A1 => n40607, A2 => n47524, B1 => n42661, B2 => 
                           n47550, ZN => n35828);
   U144 : OAI22_X1 port map( A1 => n40607, A2 => n47533, B1 => n42660, B2 => 
                           n47550, ZN => n35829);
   U145 : OAI22_X1 port map( A1 => n40607, A2 => n47523, B1 => n42659, B2 => 
                           n47550, ZN => n35830);
   U146 : OAI22_X1 port map( A1 => n40607, A2 => n47527, B1 => n42658, B2 => 
                           n47550, ZN => n35831);
   U147 : OAI22_X1 port map( A1 => n40607, A2 => n47522, B1 => n42657, B2 => 
                           n47550, ZN => n35832);
   U148 : OAI22_X1 port map( A1 => n40607, A2 => n47528, B1 => n42656, B2 => 
                           n47550, ZN => n35833);
   U149 : OAI22_X1 port map( A1 => n40607, A2 => n47520, B1 => n42655, B2 => 
                           n47550, ZN => n35834);
   U150 : OAI22_X1 port map( A1 => n40606, A2 => n47531, B1 => n42654, B2 => 
                           n47551, ZN => n35835);
   U151 : OAI22_X1 port map( A1 => n40606, A2 => n47530, B1 => n42653, B2 => 
                           n47551, ZN => n35836);
   U152 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42738, ZN => n47529);
   U153 : OAI22_X1 port map( A1 => n40606, A2 => n47529, B1 => n42652, B2 => 
                           n47551, ZN => n35837);
   U154 : OAI22_X1 port map( A1 => n40606, A2 => n47549, B1 => n42651, B2 => 
                           n47551, ZN => n35838);
   U155 : OAI22_X1 port map( A1 => n40632, A2 => n47519, B1 => n42650, B2 => 
                           n47547, ZN => n35839);
   U156 : OAI22_X1 port map( A1 => n40607, A2 => n47531, B1 => n42649, B2 => 
                           n47550, ZN => n35840);
   U157 : OAI22_X1 port map( A1 => n40632, A2 => n47516, B1 => n42648, B2 => 
                           n47547, ZN => n35841);
   U158 : OAI22_X1 port map( A1 => n40606, A2 => n47526, B1 => n42647, B2 => 
                           n47551, ZN => n35842);
   U159 : OAI22_X1 port map( A1 => n40606, A2 => n47524, B1 => n42646, B2 => 
                           n47551, ZN => n35843);
   U160 : OAI22_X1 port map( A1 => n40606, A2 => n47528, B1 => n42645, B2 => 
                           n47551, ZN => n35844);
   U161 : OAI22_X1 port map( A1 => n40606, A2 => n47520, B1 => n42644, B2 => 
                           n47551, ZN => n35845);
   U162 : OAI22_X1 port map( A1 => n40632, A2 => n47517, B1 => n42643, B2 => 
                           n47547, ZN => n35846);
   U163 : OAI22_X1 port map( A1 => n40632, A2 => n47522, B1 => n42642, B2 => 
                           n47547, ZN => n35847);
   U164 : OAI22_X1 port map( A1 => n40632, A2 => n47515, B1 => n42641, B2 => 
                           n47547, ZN => n35848);
   U165 : OAI22_X1 port map( A1 => n40632, A2 => n47527, B1 => n42640, B2 => 
                           n47547, ZN => n35849);
   U166 : OAI22_X1 port map( A1 => n40632, A2 => n47529, B1 => n42639, B2 => 
                           n47547, ZN => n35850);
   U167 : OAI22_X1 port map( A1 => n40609, A2 => n47527, B1 => n42638, B2 => 
                           n47544, ZN => n35851);
   U168 : OAI22_X1 port map( A1 => n40609, A2 => n47533, B1 => n42637, B2 => 
                           n47544, ZN => n35852);
   U169 : OAI22_X1 port map( A1 => n40609, A2 => n47524, B1 => n42636, B2 => 
                           n47544, ZN => n35853);
   U170 : OAI22_X1 port map( A1 => n40609, A2 => n47531, B1 => n42635, B2 => 
                           n47544, ZN => n35854);
   U171 : OAI22_X1 port map( A1 => n40609, A2 => n47520, B1 => n42634, B2 => 
                           n47544, ZN => n35855);
   U172 : OAI22_X1 port map( A1 => n40609, A2 => n47528, B1 => n42633, B2 => 
                           n47544, ZN => n35856);
   U173 : OAI22_X1 port map( A1 => n40606, A2 => n47523, B1 => n42632, B2 => 
                           n47551, ZN => n35857);
   U174 : OAI22_X1 port map( A1 => n40609, A2 => n47529, B1 => n42631, B2 => 
                           n47544, ZN => n35858);
   U175 : OAI22_X1 port map( A1 => n40609, A2 => n47522, B1 => n42630, B2 => 
                           n47544, ZN => n35859);
   U176 : OAI22_X1 port map( A1 => n40609, A2 => n47523, B1 => n42629, B2 => 
                           n47544, ZN => n35860);
   U177 : OAI22_X1 port map( A1 => n40609, A2 => n47530, B1 => n42628, B2 => 
                           n47544, ZN => n35861);
   U178 : OAI22_X1 port map( A1 => n40609, A2 => n47549, B1 => n42627, B2 => 
                           n47544, ZN => n35862);
   U179 : OAI22_X1 port map( A1 => n40608, A2 => n47529, B1 => n42626, B2 => 
                           n47548, ZN => n35863);
   U180 : OAI22_X1 port map( A1 => n40608, A2 => n47523, B1 => n42625, B2 => 
                           n47548, ZN => n35864);
   U181 : OAI22_X1 port map( A1 => n40608, A2 => n47528, B1 => n42624, B2 => 
                           n47548, ZN => n35865);
   U182 : OAI22_X1 port map( A1 => n40608, A2 => n47520, B1 => n42623, B2 => 
                           n47548, ZN => n35866);
   U183 : OAI22_X1 port map( A1 => n40608, A2 => n47524, B1 => n42622, B2 => 
                           n47548, ZN => n35867);
   U184 : OAI22_X1 port map( A1 => n40608, A2 => n47530, B1 => n42621, B2 => 
                           n47548, ZN => n35868);
   U185 : OAI22_X1 port map( A1 => n40608, A2 => n47533, B1 => n42620, B2 => 
                           n47548, ZN => n35869);
   U186 : OAI22_X1 port map( A1 => n40608, A2 => n47526, B1 => n42619, B2 => 
                           n47548, ZN => n35870);
   U187 : OAI22_X1 port map( A1 => n40606, A2 => n47537, B1 => n42618, B2 => 
                           n47551, ZN => n35871);
   U188 : OAI22_X1 port map( A1 => n40622, A2 => n47529, B1 => n42617, B2 => 
                           n47546, ZN => n35872);
   U189 : OAI22_X1 port map( A1 => n40622, A2 => n47528, B1 => n42616, B2 => 
                           n47546, ZN => n35873);
   U190 : OAI22_X1 port map( A1 => n40622, A2 => n47520, B1 => n42615, B2 => 
                           n47546, ZN => n35874);
   U191 : OAI22_X1 port map( A1 => n40622, A2 => n47531, B1 => n42614, B2 => 
                           n47546, ZN => n35875);
   U192 : OAI22_X1 port map( A1 => n40620, A2 => n47527, B1 => n42613, B2 => 
                           n47558, ZN => n35876);
   U193 : OAI22_X1 port map( A1 => n40620, A2 => n47533, B1 => n42612, B2 => 
                           n47558, ZN => n35877);
   U194 : OAI22_X1 port map( A1 => n40622, A2 => n47524, B1 => n42611, B2 => 
                           n47546, ZN => n35878);
   U195 : OAI22_X1 port map( A1 => n40622, A2 => n47533, B1 => n42610, B2 => 
                           n47546, ZN => n35879);
   U196 : OAI22_X1 port map( A1 => n40622, A2 => n47527, B1 => n42609, B2 => 
                           n47546, ZN => n35880);
   U197 : OAI22_X1 port map( A1 => n40620, A2 => n47524, B1 => n42608, B2 => 
                           n47558, ZN => n35881);
   U198 : OAI22_X1 port map( A1 => n40620, A2 => n47531, B1 => n42607, B2 => 
                           n47558, ZN => n35882);
   U199 : OAI22_X1 port map( A1 => n40620, A2 => n47520, B1 => n42606, B2 => 
                           n47558, ZN => n35883);
   U200 : OAI22_X1 port map( A1 => n40620, A2 => n47528, B1 => n42605, B2 => 
                           n47558, ZN => n35884);
   U201 : OAI22_X1 port map( A1 => n40620, A2 => n47530, B1 => n42604, B2 => 
                           n47558, ZN => n35885);
   U202 : OAI22_X1 port map( A1 => n40620, A2 => n47549, B1 => n42603, B2 => 
                           n47558, ZN => n35886);
   U203 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42743, ZN => n47525);
   U204 : OAI22_X1 port map( A1 => n40620, A2 => n47525, B1 => n42602, B2 => 
                           n47558, ZN => n35887);
   U205 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42745, ZN => n47521);
   U206 : OAI22_X1 port map( A1 => n40620, A2 => n47521, B1 => n42601, B2 => 
                           n47558, ZN => n35888);
   U207 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42746, ZN => n47534);
   U208 : OAI22_X1 port map( A1 => n40620, A2 => n47534, B1 => n42600, B2 => 
                           n47558, ZN => n35889);
   U209 : OAI22_X1 port map( A1 => n40612, A2 => n47526, B1 => n42599, B2 => 
                           n47559, ZN => n35890);
   U210 : OAI22_X1 port map( A1 => n40618, A2 => n47534, B1 => n42598, B2 => 
                           n47557, ZN => n35891);
   U211 : OAI22_X1 port map( A1 => n40618, A2 => n47521, B1 => n42597, B2 => 
                           n47557, ZN => n35892);
   U212 : OAI22_X1 port map( A1 => n40618, A2 => n47525, B1 => n42596, B2 => 
                           n47557, ZN => n35893);
   U213 : OAI22_X1 port map( A1 => n40618, A2 => n47549, B1 => n42595, B2 => 
                           n47557, ZN => n35894);
   U214 : OAI22_X1 port map( A1 => n40622, A2 => n47526, B1 => n42594, B2 => 
                           n47546, ZN => n35895);
   U215 : OAI22_X1 port map( A1 => n40620, A2 => n47526, B1 => n42593, B2 => 
                           n47558, ZN => n35896);
   U216 : OAI22_X1 port map( A1 => n40618, A2 => n47526, B1 => n42592, B2 => 
                           n47557, ZN => n35897);
   U217 : OAI22_X1 port map( A1 => n40616, A2 => n47526, B1 => n42591, B2 => 
                           n47560, ZN => n35898);
   U218 : OAI22_X1 port map( A1 => n40618, A2 => n47530, B1 => n42590, B2 => 
                           n47557, ZN => n35899);
   U219 : OAI22_X1 port map( A1 => n40618, A2 => n47529, B1 => n42589, B2 => 
                           n47557, ZN => n35900);
   U220 : OAI22_X1 port map( A1 => n40618, A2 => n47528, B1 => n42588, B2 => 
                           n47557, ZN => n35901);
   U221 : OAI22_X1 port map( A1 => n40618, A2 => n47520, B1 => n42587, B2 => 
                           n47557, ZN => n35902);
   U222 : OAI22_X1 port map( A1 => n40618, A2 => n47531, B1 => n42586, B2 => 
                           n47557, ZN => n35903);
   U223 : OAI22_X1 port map( A1 => n40618, A2 => n47524, B1 => n42585, B2 => 
                           n47557, ZN => n35904);
   U224 : OAI22_X1 port map( A1 => n40616, A2 => n47523, B1 => n42584, B2 => 
                           n47560, ZN => n35905);
   U225 : OAI22_X1 port map( A1 => n40626, A2 => n47515, B1 => n42583, B2 => 
                           n47553, ZN => n35906);
   U226 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42730, ZN => n47513);
   U227 : OAI22_X1 port map( A1 => n40626, A2 => n47513, B1 => n42582, B2 => 
                           n47553, ZN => n35907);
   U228 : OAI22_X1 port map( A1 => n40627, A2 => n47516, B1 => n42581, B2 => 
                           n47554, ZN => n35908);
   U229 : OAI22_X1 port map( A1 => n40627, A2 => n47513, B1 => n42580, B2 => 
                           n47554, ZN => n35909);
   U230 : OAI22_X1 port map( A1 => n40626, A2 => n47518, B1 => n42579, B2 => 
                           n47553, ZN => n35910);
   U231 : OAI22_X1 port map( A1 => n40625, A2 => n47513, B1 => n42578, B2 => 
                           n47552, ZN => n35911);
   U232 : OAI22_X1 port map( A1 => n40627, A2 => n47519, B1 => n42577, B2 => 
                           n47554, ZN => n35912);
   U233 : OAI22_X1 port map( A1 => n40627, A2 => n47529, B1 => n42576, B2 => 
                           n47554, ZN => n35913);
   U234 : OAI22_X1 port map( A1 => n40625, A2 => n47516, B1 => n42575, B2 => 
                           n47552, ZN => n35914);
   U235 : OAI22_X1 port map( A1 => n40625, A2 => n47529, B1 => n42574, B2 => 
                           n47552, ZN => n35915);
   U236 : OAI22_X1 port map( A1 => n40627, A2 => n47523, B1 => n42573, B2 => 
                           n47554, ZN => n35916);
   U237 : OAI22_X1 port map( A1 => n40625, A2 => n47515, B1 => n42572, B2 => 
                           n47552, ZN => n35917);
   U238 : OAI22_X1 port map( A1 => n40626, A2 => n47519, B1 => n42571, B2 => 
                           n47553, ZN => n35918);
   U239 : OAI22_X1 port map( A1 => n40627, A2 => n47515, B1 => n42570, B2 => 
                           n47554, ZN => n35919);
   U240 : OAI22_X1 port map( A1 => n40626, A2 => n47514, B1 => n42569, B2 => 
                           n47553, ZN => n35920);
   U241 : OAI22_X1 port map( A1 => n40625, A2 => n47514, B1 => n42568, B2 => 
                           n47552, ZN => n35921);
   U242 : OAI22_X1 port map( A1 => n40625, A2 => n47519, B1 => n42567, B2 => 
                           n47552, ZN => n35922);
   U243 : OAI22_X1 port map( A1 => n40627, A2 => n47518, B1 => n42566, B2 => 
                           n47554, ZN => n35923);
   U244 : OAI22_X1 port map( A1 => n40627, A2 => n47514, B1 => n42565, B2 => 
                           n47554, ZN => n35924);
   U245 : OAI22_X1 port map( A1 => n40626, A2 => n47516, B1 => n42564, B2 => 
                           n47553, ZN => n35925);
   U246 : OAI22_X1 port map( A1 => n40625, A2 => n47518, B1 => n42563, B2 => 
                           n47552, ZN => n35926);
   U247 : OAI22_X1 port map( A1 => n40616, A2 => n47537, B1 => n42562, B2 => 
                           n47560, ZN => n35927);
   U248 : OAI22_X1 port map( A1 => n40627, A2 => n47517, B1 => n42561, B2 => 
                           n47554, ZN => n35928);
   U249 : OAI22_X1 port map( A1 => n40612, A2 => n47537, B1 => n42560, B2 => 
                           n47559, ZN => n35929);
   U250 : OAI22_X1 port map( A1 => n40622, A2 => n47537, B1 => n42559, B2 => 
                           n47546, ZN => n35930);
   U251 : OAI22_X1 port map( A1 => n40615, A2 => n47523, B1 => n42558, B2 => 
                           n47545, ZN => n35931);
   U252 : OAI22_X1 port map( A1 => n40612, A2 => n47523, B1 => n42557, B2 => 
                           n47559, ZN => n35932);
   U253 : OAI22_X1 port map( A1 => n40618, A2 => n47533, B1 => n42556, B2 => 
                           n47557, ZN => n35933);
   U254 : OAI22_X1 port map( A1 => n40618, A2 => n47527, B1 => n42555, B2 => 
                           n47557, ZN => n35934);
   U255 : OAI22_X1 port map( A1 => n40622, A2 => n47523, B1 => n42554, B2 => 
                           n47546, ZN => n35935);
   U256 : OAI22_X1 port map( A1 => n40624, A2 => n47516, B1 => n42553, B2 => 
                           n47556, ZN => n35936);
   U257 : OAI22_X1 port map( A1 => n40624, A2 => n47513, B1 => n42552, B2 => 
                           n47556, ZN => n35937);
   U258 : OAI22_X1 port map( A1 => n40624, A2 => n47517, B1 => n42551, B2 => 
                           n47556, ZN => n35938);
   U259 : OAI22_X1 port map( A1 => n40624, A2 => n47529, B1 => n42550, B2 => 
                           n47556, ZN => n35939);
   U260 : OAI22_X1 port map( A1 => n40624, A2 => n47518, B1 => n42549, B2 => 
                           n47556, ZN => n35940);
   U261 : OAI22_X1 port map( A1 => n40624, A2 => n47514, B1 => n42548, B2 => 
                           n47556, ZN => n35941);
   U262 : OAI22_X1 port map( A1 => n40624, A2 => n47525, B1 => n42547, B2 => 
                           n47556, ZN => n35942);
   U263 : OAI22_X1 port map( A1 => n40624, A2 => n47523, B1 => n42546, B2 => 
                           n47556, ZN => n35943);
   U264 : OAI22_X1 port map( A1 => n40624, A2 => n47515, B1 => n42545, B2 => 
                           n47556, ZN => n35944);
   U265 : OAI22_X1 port map( A1 => n40624, A2 => n47519, B1 => n42544, B2 => 
                           n47556, ZN => n35945);
   U266 : OAI22_X1 port map( A1 => n40622, A2 => n47517, B1 => n42543, B2 => 
                           n47546, ZN => n35946);
   U267 : OAI22_X1 port map( A1 => n40625, A2 => n47523, B1 => n42542, B2 => 
                           n47552, ZN => n35947);
   U268 : OAI22_X1 port map( A1 => n40622, A2 => n47513, B1 => n42541, B2 => 
                           n47546, ZN => n35948);
   U269 : OAI22_X1 port map( A1 => n40622, A2 => n47518, B1 => n42540, B2 => 
                           n47546, ZN => n35949);
   U270 : OAI22_X1 port map( A1 => n40625, A2 => n47525, B1 => n42539, B2 => 
                           n47552, ZN => n35950);
   U271 : OAI22_X1 port map( A1 => n40622, A2 => n47516, B1 => n42538, B2 => 
                           n47546, ZN => n35951);
   U272 : OAI22_X1 port map( A1 => n40622, A2 => n47514, B1 => n42537, B2 => 
                           n47546, ZN => n35952);
   U273 : OAI22_X1 port map( A1 => n40622, A2 => n47519, B1 => n42536, B2 => 
                           n47546, ZN => n35953);
   U274 : OAI22_X1 port map( A1 => n40622, A2 => n47515, B1 => n42535, B2 => 
                           n47546, ZN => n35954);
   U275 : OAI22_X1 port map( A1 => n40626, A2 => n47529, B1 => n42534, B2 => 
                           n47553, ZN => n35955);
   U276 : OAI22_X1 port map( A1 => n40626, A2 => n47523, B1 => n42533, B2 => 
                           n47553, ZN => n35956);
   U277 : OAI22_X1 port map( A1 => n40626, A2 => n47517, B1 => n42532, B2 => 
                           n47553, ZN => n35957);
   U278 : OAI22_X1 port map( A1 => n40625, A2 => n47517, B1 => n42531, B2 => 
                           n47552, ZN => n35958);
   U279 : OAI22_X1 port map( A1 => n40622, A2 => n47522, B1 => n42530, B2 => 
                           n47546, ZN => n35959);
   U280 : OAI22_X1 port map( A1 => n40626, A2 => n47530, B1 => n42529, B2 => 
                           n47553, ZN => n35960);
   U281 : OAI22_X1 port map( A1 => n40620, A2 => n47522, B1 => n42528, B2 => 
                           n47558, ZN => n35961);
   U282 : OAI22_X1 port map( A1 => n40627, A2 => n47527, B1 => n42527, B2 => 
                           n47554, ZN => n35962);
   U283 : OAI22_X1 port map( A1 => n40626, A2 => n47533, B1 => n42526, B2 => 
                           n47553, ZN => n35963);
   U284 : OAI22_X1 port map( A1 => n40627, A2 => n47528, B1 => n42525, B2 => 
                           n47554, ZN => n35964);
   U285 : OAI22_X1 port map( A1 => n40626, A2 => n47527, B1 => n42524, B2 => 
                           n47553, ZN => n35965);
   U286 : OAI22_X1 port map( A1 => n40626, A2 => n47528, B1 => n42523, B2 => 
                           n47553, ZN => n35966);
   U287 : OAI22_X1 port map( A1 => n40627, A2 => n47531, B1 => n42522, B2 => 
                           n47554, ZN => n35967);
   U288 : OAI22_X1 port map( A1 => n40626, A2 => n47531, B1 => n42521, B2 => 
                           n47553, ZN => n35968);
   U289 : OAI22_X1 port map( A1 => n40607, A2 => n47513, B1 => n42520, B2 => 
                           n47550, ZN => n35969);
   U290 : OAI22_X1 port map( A1 => n40609, A2 => n47513, B1 => n42519, B2 => 
                           n47544, ZN => n35970);
   U291 : OAI22_X1 port map( A1 => n40612, A2 => n47522, B1 => n42518, B2 => 
                           n47559, ZN => n35971);
   U292 : OAI22_X1 port map( A1 => n40606, A2 => n47513, B1 => n42517, B2 => 
                           n47551, ZN => n35972);
   U293 : OAI22_X1 port map( A1 => n40608, A2 => n47513, B1 => n42516, B2 => 
                           n47548, ZN => n35973);
   U294 : OAI22_X1 port map( A1 => n40608, A2 => n47534, B1 => n42515, B2 => 
                           n47548, ZN => n35974);
   U295 : OAI22_X1 port map( A1 => n40608, A2 => n47521, B1 => n42514, B2 => 
                           n47548, ZN => n35975);
   U296 : OAI22_X1 port map( A1 => n40627, A2 => n47534, B1 => n42513, B2 => 
                           n47554, ZN => n35976);
   U297 : OAI22_X1 port map( A1 => n40627, A2 => n47521, B1 => n42512, B2 => 
                           n47554, ZN => n35977);
   U298 : OAI22_X1 port map( A1 => n40626, A2 => n47534, B1 => n42511, B2 => 
                           n47553, ZN => n35978);
   U299 : OAI22_X1 port map( A1 => n40626, A2 => n47521, B1 => n42510, B2 => 
                           n47553, ZN => n35979);
   U300 : OAI22_X1 port map( A1 => n40625, A2 => n47534, B1 => n42509, B2 => 
                           n47552, ZN => n35980);
   U301 : OAI22_X1 port map( A1 => n40625, A2 => n47521, B1 => n42508, B2 => 
                           n47552, ZN => n35981);
   U302 : OAI22_X1 port map( A1 => n40607, A2 => n47521, B1 => n42507, B2 => 
                           n47550, ZN => n35982);
   U303 : OAI22_X1 port map( A1 => n40607, A2 => n47525, B1 => n42506, B2 => 
                           n47550, ZN => n35983);
   U304 : OAI22_X1 port map( A1 => n40609, A2 => n47521, B1 => n42505, B2 => 
                           n47544, ZN => n35984);
   U305 : OAI22_X1 port map( A1 => n40606, A2 => n47521, B1 => n42504, B2 => 
                           n47551, ZN => n35985);
   U306 : OAI22_X1 port map( A1 => n40615, A2 => n47522, B1 => n42503, B2 => 
                           n47545, ZN => n35986);
   U307 : OAI22_X1 port map( A1 => n40616, A2 => n47522, B1 => n42502, B2 => 
                           n47560, ZN => n35987);
   U308 : OAI22_X1 port map( A1 => n40609, A2 => n47525, B1 => n42501, B2 => 
                           n47544, ZN => n35988);
   U309 : OAI22_X1 port map( A1 => n40626, A2 => n47537, B1 => n42500, B2 => 
                           n47553, ZN => n35989);
   U310 : OAI22_X1 port map( A1 => n40625, A2 => n47537, B1 => n42499, B2 => 
                           n47552, ZN => n35990);
   U311 : OAI22_X1 port map( A1 => n40627, A2 => n47537, B1 => n42498, B2 => 
                           n47554, ZN => n35991);
   U312 : OAI22_X1 port map( A1 => n40608, A2 => n47525, B1 => n42497, B2 => 
                           n47548, ZN => n35992);
   U313 : OAI22_X1 port map( A1 => n40620, A2 => n47555, B1 => n42496, B2 => 
                           n47558, ZN => n35993);
   U314 : OAI22_X1 port map( A1 => n40632, A2 => n47555, B1 => n42495, B2 => 
                           n47547, ZN => n35994);
   U315 : OAI22_X1 port map( A1 => n40606, A2 => n47534, B1 => n42494, B2 => 
                           n47551, ZN => n35995);
   U316 : OAI22_X1 port map( A1 => n40615, A2 => n47555, B1 => n42493, B2 => 
                           n47545, ZN => n35996);
   U317 : OAI22_X1 port map( A1 => n40624, A2 => n47531, B1 => n42492, B2 => 
                           n47556, ZN => n35997);
   U318 : OAI22_X1 port map( A1 => n40624, A2 => n47537, B1 => n42491, B2 => 
                           n47556, ZN => n35998);
   U319 : OAI22_X1 port map( A1 => n40624, A2 => n47524, B1 => n42490, B2 => 
                           n47556, ZN => n35999);
   U320 : OAI22_X1 port map( A1 => n40632, A2 => n47513, B1 => n42489, B2 => 
                           n47547, ZN => n36000);
   U321 : OAI22_X1 port map( A1 => n40624, A2 => n47521, B1 => n42488, B2 => 
                           n47556, ZN => n36001);
   U322 : OAI22_X1 port map( A1 => n40624, A2 => n47522, B1 => n42487, B2 => 
                           n47556, ZN => n36002);
   U323 : OAI22_X1 port map( A1 => n40624, A2 => n47520, B1 => n42486, B2 => 
                           n47556, ZN => n36003);
   U324 : OAI22_X1 port map( A1 => n40632, A2 => n47525, B1 => n42485, B2 => 
                           n47547, ZN => n36004);
   U325 : OAI22_X1 port map( A1 => n40624, A2 => n47530, B1 => n42484, B2 => 
                           n47556, ZN => n36005);
   U326 : OAI22_X1 port map( A1 => n40624, A2 => n47527, B1 => n42483, B2 => 
                           n47556, ZN => n36006);
   U327 : OAI22_X1 port map( A1 => n40624, A2 => n47534, B1 => n42482, B2 => 
                           n47556, ZN => n36007);
   U328 : OAI22_X1 port map( A1 => n40624, A2 => n47533, B1 => n42481, B2 => 
                           n47556, ZN => n36008);
   U329 : OAI22_X1 port map( A1 => n40624, A2 => n47528, B1 => n42480, B2 => 
                           n47556, ZN => n36009);
   U330 : OAI22_X1 port map( A1 => n40615, A2 => n47528, B1 => n42479, B2 => 
                           n47545, ZN => n36010);
   U331 : OAI22_X1 port map( A1 => n40615, A2 => n47525, B1 => n42478, B2 => 
                           n47545, ZN => n36011);
   U332 : OAI22_X1 port map( A1 => n40616, A2 => n47528, B1 => n42477, B2 => 
                           n47560, ZN => n36012);
   U333 : OAI22_X1 port map( A1 => n40616, A2 => n47525, B1 => n42476, B2 => 
                           n47560, ZN => n36013);
   U334 : OAI22_X1 port map( A1 => n40615, A2 => n47534, B1 => n42475, B2 => 
                           n47545, ZN => n36014);
   U335 : OAI22_X1 port map( A1 => n40616, A2 => n47534, B1 => n42474, B2 => 
                           n47560, ZN => n36015);
   U336 : OAI22_X1 port map( A1 => n40622, A2 => n47534, B1 => n42473, B2 => 
                           n47546, ZN => n36016);
   U337 : OAI22_X1 port map( A1 => n40615, A2 => n47521, B1 => n42472, B2 => 
                           n47545, ZN => n36017);
   U338 : OAI22_X1 port map( A1 => n40632, A2 => n47534, B1 => n42471, B2 => 
                           n47547, ZN => n36018);
   U339 : OAI22_X1 port map( A1 => n40632, A2 => n47521, B1 => n42470, B2 => 
                           n47547, ZN => n36019);
   U340 : OAI22_X1 port map( A1 => n40616, A2 => n47521, B1 => n42469, B2 => 
                           n47560, ZN => n36020);
   U341 : OAI22_X1 port map( A1 => n40615, A2 => n47530, B1 => n42468, B2 => 
                           n47545, ZN => n36021);
   U342 : OAI22_X1 port map( A1 => n40615, A2 => n47527, B1 => n42467, B2 => 
                           n47545, ZN => n36022);
   U343 : OAI22_X1 port map( A1 => n40608, A2 => n47522, B1 => n42466, B2 => 
                           n47548, ZN => n36023);
   U344 : OAI22_X1 port map( A1 => n40616, A2 => n47527, B1 => n42465, B2 => 
                           n47560, ZN => n36024);
   U345 : OAI22_X1 port map( A1 => n40612, A2 => n47528, B1 => n42464, B2 => 
                           n47559, ZN => n36025);
   U346 : OAI22_X1 port map( A1 => n40612, A2 => n47527, B1 => n42463, B2 => 
                           n47559, ZN => n36026);
   U347 : OAI22_X1 port map( A1 => n40612, A2 => n47530, B1 => n42462, B2 => 
                           n47559, ZN => n36027);
   U348 : OAI22_X1 port map( A1 => n40612, A2 => n47525, B1 => n42461, B2 => 
                           n47559, ZN => n36028);
   U349 : OAI22_X1 port map( A1 => n40612, A2 => n47521, B1 => n42460, B2 => 
                           n47559, ZN => n36029);
   U350 : OAI22_X1 port map( A1 => n40612, A2 => n47533, B1 => n42459, B2 => 
                           n47559, ZN => n36030);
   U351 : OAI22_X1 port map( A1 => n40616, A2 => n47529, B1 => n42458, B2 => 
                           n47560, ZN => n36031);
   U352 : OAI22_X1 port map( A1 => n40622, A2 => n47521, B1 => n42457, B2 => 
                           n47546, ZN => n36032);
   U353 : OAI22_X1 port map( A1 => n40615, A2 => n47513, B1 => n42456, B2 => 
                           n47545, ZN => n36033);
   U354 : OAI22_X1 port map( A1 => n40612, A2 => n47514, B1 => n42455, B2 => 
                           n47559, ZN => n36034);
   U355 : OAI22_X1 port map( A1 => n40615, A2 => n47529, B1 => n42454, B2 => 
                           n47545, ZN => n36035);
   U356 : OAI22_X1 port map( A1 => n40618, A2 => n47537, B1 => n42453, B2 => 
                           n47557, ZN => n36036);
   U357 : OAI22_X1 port map( A1 => n40616, A2 => n47515, B1 => n42452, B2 => 
                           n47560, ZN => n36037);
   U358 : OAI22_X1 port map( A1 => n40618, A2 => n47519, B1 => n42451, B2 => 
                           n47557, ZN => n36038);
   U359 : OAI22_X1 port map( A1 => n40616, A2 => n47513, B1 => n42450, B2 => 
                           n47560, ZN => n36039);
   U360 : OAI22_X1 port map( A1 => n40612, A2 => n47517, B1 => n42449, B2 => 
                           n47559, ZN => n36040);
   U361 : OAI22_X1 port map( A1 => n40616, A2 => n47519, B1 => n42448, B2 => 
                           n47560, ZN => n36041);
   U362 : OAI22_X1 port map( A1 => n40615, A2 => n47515, B1 => n42447, B2 => 
                           n47545, ZN => n36042);
   U363 : OAI22_X1 port map( A1 => n40615, A2 => n47519, B1 => n42446, B2 => 
                           n47545, ZN => n36043);
   U364 : OAI22_X1 port map( A1 => n40616, A2 => n47555, B1 => n42445, B2 => 
                           n47560, ZN => n36044);
   U365 : OAI22_X1 port map( A1 => n40612, A2 => n47529, B1 => n42444, B2 => 
                           n47559, ZN => n36045);
   U366 : OAI22_X1 port map( A1 => n40618, A2 => n47518, B1 => n42443, B2 => 
                           n47557, ZN => n36046);
   U367 : OAI22_X1 port map( A1 => n40612, A2 => n47524, B1 => n42442, B2 => 
                           n47559, ZN => n36047);
   U368 : OAI22_X1 port map( A1 => n40618, A2 => n47516, B1 => n42441, B2 => 
                           n47557, ZN => n36048);
   U369 : OAI22_X1 port map( A1 => n40616, A2 => n47516, B1 => n42440, B2 => 
                           n47560, ZN => n36049);
   U370 : OAI22_X1 port map( A1 => n40615, A2 => n47516, B1 => n42439, B2 => 
                           n47545, ZN => n36050);
   U371 : OAI22_X1 port map( A1 => n40612, A2 => n47518, B1 => n42438, B2 => 
                           n47559, ZN => n36051);
   U372 : OAI22_X1 port map( A1 => n40622, A2 => n47525, B1 => n42437, B2 => 
                           n47546, ZN => n36052);
   U373 : OAI22_X1 port map( A1 => n40618, A2 => n47517, B1 => n42436, B2 => 
                           n47557, ZN => n36053);
   U374 : OAI22_X1 port map( A1 => n40620, A2 => n47515, B1 => n42435, B2 => 
                           n47558, ZN => n36054);
   U375 : OAI22_X1 port map( A1 => n40615, A2 => n47537, B1 => n42434, B2 => 
                           n47545, ZN => n36055);
   U376 : OAI22_X1 port map( A1 => n40620, A2 => n47516, B1 => n42433, B2 => 
                           n47558, ZN => n36056);
   U377 : OAI22_X1 port map( A1 => n40620, A2 => n47517, B1 => n42432, B2 => 
                           n47558, ZN => n36057);
   U378 : OAI22_X1 port map( A1 => n40615, A2 => n47524, B1 => n42431, B2 => 
                           n47545, ZN => n36058);
   U379 : OAI22_X1 port map( A1 => n40620, A2 => n47537, B1 => n42430, B2 => 
                           n47558, ZN => n36059);
   U380 : OAI22_X1 port map( A1 => n40612, A2 => n47519, B1 => n42429, B2 => 
                           n47559, ZN => n36060);
   U381 : OAI22_X1 port map( A1 => n40616, A2 => n47524, B1 => n42428, B2 => 
                           n47560, ZN => n36061);
   U382 : OAI22_X1 port map( A1 => n40620, A2 => n47519, B1 => n42427, B2 => 
                           n47558, ZN => n36062);
   U383 : OAI22_X1 port map( A1 => n40615, A2 => n47518, B1 => n42426, B2 => 
                           n47545, ZN => n36063);
   U384 : OAI22_X1 port map( A1 => n40612, A2 => n47531, B1 => n42425, B2 => 
                           n47559, ZN => n36064);
   U385 : OAI22_X1 port map( A1 => n40612, A2 => n47513, B1 => n42424, B2 => 
                           n47559, ZN => n36065);
   U386 : OAI22_X1 port map( A1 => n40615, A2 => n47531, B1 => n42423, B2 => 
                           n47545, ZN => n36066);
   U387 : OAI22_X1 port map( A1 => n40616, A2 => n47518, B1 => n42422, B2 => 
                           n47560, ZN => n36067);
   U388 : OAI22_X1 port map( A1 => n40612, A2 => n47520, B1 => n42421, B2 => 
                           n47559, ZN => n36068);
   U389 : OAI22_X1 port map( A1 => n40615, A2 => n47514, B1 => n42420, B2 => 
                           n47545, ZN => n36069);
   U390 : OAI22_X1 port map( A1 => n40620, A2 => n47518, B1 => n42419, B2 => 
                           n47558, ZN => n36070);
   U391 : OAI22_X1 port map( A1 => n40616, A2 => n47531, B1 => n42418, B2 => 
                           n47560, ZN => n36071);
   U392 : OAI22_X1 port map( A1 => n40616, A2 => n47514, B1 => n42417, B2 => 
                           n47560, ZN => n36072);
   U393 : OAI22_X1 port map( A1 => n40618, A2 => n47513, B1 => n42416, B2 => 
                           n47557, ZN => n36073);
   U394 : OAI22_X1 port map( A1 => n40615, A2 => n47517, B1 => n42415, B2 => 
                           n47545, ZN => n36074);
   U395 : OAI22_X1 port map( A1 => n40612, A2 => n47515, B1 => n42414, B2 => 
                           n47559, ZN => n36075);
   U396 : OAI22_X1 port map( A1 => n40616, A2 => n47520, B1 => n42413, B2 => 
                           n47560, ZN => n36076);
   U397 : OAI22_X1 port map( A1 => n40612, A2 => n47516, B1 => n42412, B2 => 
                           n47559, ZN => n36077);
   U398 : OAI22_X1 port map( A1 => n40620, A2 => n47514, B1 => n42411, B2 => 
                           n47558, ZN => n36078);
   U399 : OAI22_X1 port map( A1 => n40618, A2 => n47515, B1 => n42410, B2 => 
                           n47557, ZN => n36079);
   U400 : OAI22_X1 port map( A1 => n40615, A2 => n47520, B1 => n42409, B2 => 
                           n47545, ZN => n36080);
   U401 : OAI22_X1 port map( A1 => n40616, A2 => n47517, B1 => n42408, B2 => 
                           n47560, ZN => n36081);
   U402 : OAI22_X1 port map( A1 => n40618, A2 => n47514, B1 => n42407, B2 => 
                           n47557, ZN => n36082);
   U403 : OAI22_X1 port map( A1 => n40628, A2 => n47522, B1 => n42406, B2 => 
                           n47512, ZN => n36083);
   U404 : OAI22_X1 port map( A1 => n40637, A2 => n47522, B1 => n42405, B2 => 
                           n47511, ZN => n36084);
   U405 : OAI22_X1 port map( A1 => n40638, A2 => n47522, B1 => n42404, B2 => 
                           n47563, ZN => n36085);
   U406 : OAI22_X1 port map( A1 => n40642, A2 => n47522, B1 => n42403, B2 => 
                           n47561, ZN => n36086);
   U407 : OAI22_X1 port map( A1 => n40646, A2 => n47522, B1 => n42402, B2 => 
                           n47562, ZN => n36087);
   U408 : OAI22_X1 port map( A1 => n40637, A2 => n47524, B1 => n42401, B2 => 
                           n47511, ZN => n36088);
   U409 : OAI22_X1 port map( A1 => n40647, A2 => n47549, B1 => n42400, B2 => 
                           n47567, ZN => n36089);
   U410 : OAI22_X1 port map( A1 => n40638, A2 => n47524, B1 => n42399, B2 => 
                           n47563, ZN => n36090);
   U411 : OAI22_X1 port map( A1 => n40642, A2 => n47524, B1 => n42398, B2 => 
                           n47561, ZN => n36091);
   U412 : OAI22_X1 port map( A1 => n40646, A2 => n47524, B1 => n42397, B2 => 
                           n47562, ZN => n36092);
   U413 : OAI22_X1 port map( A1 => n40647, A2 => n47524, B1 => n42396, B2 => 
                           n47567, ZN => n36093);
   U414 : OAI22_X1 port map( A1 => n40628, A2 => n47524, B1 => n42395, B2 => 
                           n47512, ZN => n36094);
   U415 : OAI22_X1 port map( A1 => n40647, A2 => n47523, B1 => n42394, B2 => 
                           n47567, ZN => n36095);
   U416 : OAI22_X1 port map( A1 => n40637, A2 => n47531, B1 => n42393, B2 => 
                           n47511, ZN => n36096);
   U417 : OAI22_X1 port map( A1 => n40638, A2 => n47531, B1 => n42392, B2 => 
                           n47563, ZN => n36097);
   U418 : OAI22_X1 port map( A1 => n40642, A2 => n47531, B1 => n42391, B2 => 
                           n47561, ZN => n36098);
   U419 : OAI22_X1 port map( A1 => n40647, A2 => n47531, B1 => n42390, B2 => 
                           n47567, ZN => n36099);
   U420 : OAI22_X1 port map( A1 => n40647, A2 => n47530, B1 => n42389, B2 => 
                           n47567, ZN => n36100);
   U421 : OAI22_X1 port map( A1 => n40628, A2 => n47531, B1 => n42388, B2 => 
                           n47512, ZN => n36101);
   U422 : OAI22_X1 port map( A1 => n40637, A2 => n47520, B1 => n42387, B2 => 
                           n47511, ZN => n36102);
   U423 : OAI22_X1 port map( A1 => n40642, A2 => n47520, B1 => n42386, B2 => 
                           n47561, ZN => n36103);
   U424 : OAI22_X1 port map( A1 => n40646, A2 => n47520, B1 => n42385, B2 => 
                           n47562, ZN => n36104);
   U425 : OAI22_X1 port map( A1 => n40647, A2 => n47520, B1 => n42384, B2 => 
                           n47567, ZN => n36105);
   U426 : OAI22_X1 port map( A1 => n40628, A2 => n47520, B1 => n42383, B2 => 
                           n47512, ZN => n36106);
   U427 : OAI22_X1 port map( A1 => n40638, A2 => n47528, B1 => n42382, B2 => 
                           n47563, ZN => n36107);
   U428 : OAI22_X1 port map( A1 => n40637, A2 => n47528, B1 => n42381, B2 => 
                           n47511, ZN => n36108);
   U429 : OAI22_X1 port map( A1 => n40647, A2 => n47529, B1 => n42380, B2 => 
                           n47567, ZN => n36109);
   U430 : OAI22_X1 port map( A1 => n40646, A2 => n47528, B1 => n42379, B2 => 
                           n47562, ZN => n36110);
   U431 : OAI22_X1 port map( A1 => n40642, A2 => n47528, B1 => n42378, B2 => 
                           n47561, ZN => n36111);
   U432 : OAI22_X1 port map( A1 => n40638, A2 => n47527, B1 => n42377, B2 => 
                           n47563, ZN => n36112);
   U433 : OAI22_X1 port map( A1 => n40646, A2 => n47527, B1 => n42376, B2 => 
                           n47562, ZN => n36113);
   U434 : OAI22_X1 port map( A1 => n40647, A2 => n47527, B1 => n42375, B2 => 
                           n47567, ZN => n36114);
   U435 : OAI22_X1 port map( A1 => n40642, A2 => n47527, B1 => n42374, B2 => 
                           n47561, ZN => n36115);
   U436 : OAI22_X1 port map( A1 => n40637, A2 => n47527, B1 => n42373, B2 => 
                           n47511, ZN => n36116);
   U437 : OAI22_X1 port map( A1 => n40628, A2 => n47527, B1 => n42372, B2 => 
                           n47512, ZN => n36117);
   U438 : OAI22_X1 port map( A1 => n40628, A2 => n47533, B1 => n42371, B2 => 
                           n47512, ZN => n36118);
   U439 : OAI22_X1 port map( A1 => n40646, A2 => n47533, B1 => n42370, B2 => 
                           n47562, ZN => n36119);
   U440 : OAI22_X1 port map( A1 => n40637, A2 => n47533, B1 => n42369, B2 => 
                           n47511, ZN => n36120);
   U441 : OAI22_X1 port map( A1 => n40642, A2 => n47533, B1 => n42368, B2 => 
                           n47561, ZN => n36121);
   U442 : OAI22_X1 port map( A1 => n40638, A2 => n47533, B1 => n42367, B2 => 
                           n47563, ZN => n36122);
   U443 : OAI22_X1 port map( A1 => n40647, A2 => n47533, B1 => n42366, B2 => 
                           n47567, ZN => n36123);
   U444 : OAI22_X1 port map( A1 => n40604, A2 => n47527, B1 => n42365, B2 => 
                           n47566, ZN => n36124);
   U445 : OAI22_X1 port map( A1 => n40604, A2 => n47533, B1 => n42364, B2 => 
                           n47566, ZN => n36125);
   U446 : OAI22_X1 port map( A1 => n40604, A2 => n47524, B1 => n42363, B2 => 
                           n47566, ZN => n36126);
   U447 : OAI22_X1 port map( A1 => n40604, A2 => n47520, B1 => n42362, B2 => 
                           n47566, ZN => n36127);
   U448 : OAI22_X1 port map( A1 => n40605, A2 => n47526, B1 => n42361, B2 => 
                           n47565, ZN => n36128);
   U449 : OAI22_X1 port map( A1 => n40605, A2 => n47549, B1 => n42360, B2 => 
                           n47565, ZN => n36129);
   U450 : OAI22_X1 port map( A1 => n40605, A2 => n47530, B1 => n42359, B2 => 
                           n47565, ZN => n36130);
   U451 : OAI22_X1 port map( A1 => n40604, A2 => n47522, B1 => n42358, B2 => 
                           n47566, ZN => n36131);
   U452 : OAI22_X1 port map( A1 => n40605, A2 => n47523, B1 => n42357, B2 => 
                           n47565, ZN => n36132);
   U453 : OAI22_X1 port map( A1 => n40605, A2 => n47522, B1 => n42356, B2 => 
                           n47565, ZN => n36133);
   U454 : OAI22_X1 port map( A1 => n40605, A2 => n47529, B1 => n42355, B2 => 
                           n47565, ZN => n36134);
   U455 : OAI22_X1 port map( A1 => n40605, A2 => n47528, B1 => n42354, B2 => 
                           n47565, ZN => n36135);
   U456 : OAI22_X1 port map( A1 => n40605, A2 => n47520, B1 => n42353, B2 => 
                           n47565, ZN => n36136);
   U457 : OAI22_X1 port map( A1 => n40605, A2 => n47524, B1 => n42352, B2 => 
                           n47565, ZN => n36137);
   U458 : OAI22_X1 port map( A1 => n40605, A2 => n47533, B1 => n42351, B2 => 
                           n47565, ZN => n36138);
   U459 : OAI22_X1 port map( A1 => n40605, A2 => n47527, B1 => n42350, B2 => 
                           n47565, ZN => n36139);
   U460 : OAI22_X1 port map( A1 => n40604, A2 => n47526, B1 => n42349, B2 => 
                           n47566, ZN => n36140);
   U461 : OAI22_X1 port map( A1 => n40604, A2 => n47549, B1 => n42348, B2 => 
                           n47566, ZN => n36141);
   U462 : OAI22_X1 port map( A1 => n40604, A2 => n47530, B1 => n42347, B2 => 
                           n47566, ZN => n36142);
   U463 : OAI22_X1 port map( A1 => n40604, A2 => n47523, B1 => n42346, B2 => 
                           n47566, ZN => n36143);
   U464 : OAI22_X1 port map( A1 => n40604, A2 => n47529, B1 => n42345, B2 => 
                           n47566, ZN => n36144);
   U465 : OAI22_X1 port map( A1 => n40637, A2 => n47534, B1 => n42344, B2 => 
                           n47511, ZN => n36145);
   U466 : OAI22_X1 port map( A1 => n40628, A2 => n47521, B1 => n42343, B2 => 
                           n47512, ZN => n36146);
   U467 : OAI22_X1 port map( A1 => n40642, A2 => n47525, B1 => n42342, B2 => 
                           n47561, ZN => n36147);
   U468 : OAI22_X1 port map( A1 => n40647, A2 => n47513, B1 => n42341, B2 => 
                           n47567, ZN => n36148);
   U469 : OAI22_X1 port map( A1 => n40638, A2 => n47521, B1 => n42340, B2 => 
                           n47563, ZN => n36149);
   U470 : OAI22_X1 port map( A1 => n40647, A2 => n47525, B1 => n42339, B2 => 
                           n47567, ZN => n36150);
   U471 : OAI22_X1 port map( A1 => n40638, A2 => n47525, B1 => n42338, B2 => 
                           n47563, ZN => n36151);
   U472 : OAI22_X1 port map( A1 => n40638, A2 => n47513, B1 => n42337, B2 => 
                           n47563, ZN => n36152);
   U473 : OAI22_X1 port map( A1 => n40642, A2 => n47513, B1 => n42336, B2 => 
                           n47561, ZN => n36153);
   U474 : OAI22_X1 port map( A1 => n40646, A2 => n47521, B1 => n42335, B2 => 
                           n47562, ZN => n36154);
   U475 : OAI22_X1 port map( A1 => n40646, A2 => n47525, B1 => n42334, B2 => 
                           n47562, ZN => n36155);
   U476 : OAI22_X1 port map( A1 => n40628, A2 => n47525, B1 => n42333, B2 => 
                           n47512, ZN => n36156);
   U477 : OAI22_X1 port map( A1 => n40637, A2 => n47525, B1 => n42332, B2 => 
                           n47511, ZN => n36157);
   U478 : OAI22_X1 port map( A1 => n40604, A2 => n47555, B1 => n42331, B2 => 
                           n47566, ZN => n36158);
   U479 : OAI22_X1 port map( A1 => n40605, A2 => n47555, B1 => n42330, B2 => 
                           n47565, ZN => n36159);
   U480 : OAI22_X1 port map( A1 => n40646, A2 => n47513, B1 => n42329, B2 => 
                           n47562, ZN => n36160);
   U481 : OAI22_X1 port map( A1 => n40605, A2 => n47514, B1 => n42328, B2 => 
                           n47565, ZN => n36161);
   U482 : OAI22_X1 port map( A1 => n40628, A2 => n47513, B1 => n42327, B2 => 
                           n47512, ZN => n36162);
   U483 : OAI22_X1 port map( A1 => n40605, A2 => n47518, B1 => n42326, B2 => 
                           n47565, ZN => n36163);
   U484 : OAI22_X1 port map( A1 => n40605, A2 => n47515, B1 => n42325, B2 => 
                           n47565, ZN => n36164);
   U485 : OAI22_X1 port map( A1 => n40605, A2 => n47516, B1 => n42324, B2 => 
                           n47565, ZN => n36165);
   U486 : OAI22_X1 port map( A1 => n40605, A2 => n47517, B1 => n42323, B2 => 
                           n47565, ZN => n36166);
   U487 : OAI22_X1 port map( A1 => n40604, A2 => n47519, B1 => n42322, B2 => 
                           n47566, ZN => n36167);
   U488 : OAI22_X1 port map( A1 => n40604, A2 => n47517, B1 => n42321, B2 => 
                           n47566, ZN => n36168);
   U489 : OAI22_X1 port map( A1 => n40604, A2 => n47516, B1 => n42320, B2 => 
                           n47566, ZN => n36169);
   U490 : OAI22_X1 port map( A1 => n40604, A2 => n47515, B1 => n42319, B2 => 
                           n47566, ZN => n36170);
   U491 : OAI22_X1 port map( A1 => n40604, A2 => n47518, B1 => n42318, B2 => 
                           n47566, ZN => n36171);
   U492 : OAI22_X1 port map( A1 => n40605, A2 => n47519, B1 => n42317, B2 => 
                           n47565, ZN => n36172);
   U493 : OAI22_X1 port map( A1 => n40637, A2 => n47513, B1 => n42316, B2 => 
                           n47511, ZN => n36173);
   U494 : OAI22_X1 port map( A1 => n40604, A2 => n47514, B1 => n42315, B2 => 
                           n47566, ZN => n36174);
   U495 : OAI22_X1 port map( A1 => n40646, A2 => n47555, B1 => n42314, B2 => 
                           n47562, ZN => n36175);
   U496 : OAI22_X1 port map( A1 => n40628, A2 => n47537, B1 => n42313, B2 => 
                           n47512, ZN => n36176);
   U497 : OAI22_X1 port map( A1 => n40637, A2 => n47537, B1 => n42312, B2 => 
                           n47511, ZN => n36177);
   U498 : OAI22_X1 port map( A1 => n40647, A2 => n47555, B1 => n42311, B2 => 
                           n47567, ZN => n36178);
   U499 : OAI22_X1 port map( A1 => n40646, A2 => n47537, B1 => n42310, B2 => 
                           n47562, ZN => n36179);
   U500 : OAI22_X1 port map( A1 => n40642, A2 => n47555, B1 => n42309, B2 => 
                           n47561, ZN => n36180);
   U501 : OAI22_X1 port map( A1 => n40647, A2 => n47537, B1 => n42308, B2 => 
                           n47567, ZN => n36181);
   U502 : OAI22_X1 port map( A1 => n40637, A2 => n47555, B1 => n42307, B2 => 
                           n47511, ZN => n36182);
   U503 : OAI22_X1 port map( A1 => n40642, A2 => n47537, B1 => n42306, B2 => 
                           n47561, ZN => n36183);
   U504 : OAI22_X1 port map( A1 => n40638, A2 => n47555, B1 => n42305, B2 => 
                           n47563, ZN => n36185);
   U505 : OAI22_X1 port map( A1 => n40642, A2 => n47523, B1 => n42304, B2 => 
                           n47561, ZN => n36186);
   U506 : OAI22_X1 port map( A1 => n40646, A2 => n47523, B1 => n42303, B2 => 
                           n47562, ZN => n36187);
   U507 : OAI22_X1 port map( A1 => n40628, A2 => n47555, B1 => n42302, B2 => 
                           n47512, ZN => n36188);
   U508 : OAI22_X1 port map( A1 => n40605, A2 => n47513, B1 => n42301, B2 => 
                           n47565, ZN => n36189);
   U509 : OAI22_X1 port map( A1 => n40604, A2 => n47513, B1 => n42300, B2 => 
                           n47566, ZN => n36190);
   U510 : OAI22_X1 port map( A1 => n40647, A2 => n47519, B1 => n42299, B2 => 
                           n47567, ZN => n36191);
   U511 : OAI22_X1 port map( A1 => n40628, A2 => n47523, B1 => n42298, B2 => 
                           n47512, ZN => n36192);
   U512 : OAI22_X1 port map( A1 => n40647, A2 => n47522, B1 => n42297, B2 => 
                           n47567, ZN => n36193);
   U513 : OAI22_X1 port map( A1 => n40638, A2 => n47515, B1 => n42296, B2 => 
                           n47563, ZN => n36194);
   U514 : OAI22_X1 port map( A1 => n40637, A2 => n47523, B1 => n42295, B2 => 
                           n47511, ZN => n36195);
   U515 : OAI22_X1 port map( A1 => n40628, A2 => n47519, B1 => n42294, B2 => 
                           n47512, ZN => n36196);
   U516 : OAI22_X1 port map( A1 => n40638, A2 => n47523, B1 => n42293, B2 => 
                           n47563, ZN => n36197);
   U517 : OAI22_X1 port map( A1 => n40628, A2 => n47515, B1 => n42292, B2 => 
                           n47512, ZN => n36198);
   U518 : OAI22_X1 port map( A1 => n40647, A2 => n47521, B1 => n42291, B2 => 
                           n47567, ZN => n36199);
   U519 : OAI22_X1 port map( A1 => n40637, A2 => n47517, B1 => n42290, B2 => 
                           n47511, ZN => n36200);
   U520 : OAI22_X1 port map( A1 => n40647, A2 => n47528, B1 => n42289, B2 => 
                           n47567, ZN => n36201);
   U521 : OAI22_X1 port map( A1 => n40638, A2 => n47517, B1 => n42288, B2 => 
                           n47563, ZN => n36202);
   U522 : OAI22_X1 port map( A1 => n40646, A2 => n47519, B1 => n42287, B2 => 
                           n47562, ZN => n36203);
   U523 : OAI22_X1 port map( A1 => n40642, A2 => n47519, B1 => n42286, B2 => 
                           n47561, ZN => n36204);
   U524 : OAI22_X1 port map( A1 => n40638, A2 => n47519, B1 => n42285, B2 => 
                           n47563, ZN => n36205);
   U525 : OAI22_X1 port map( A1 => n40637, A2 => n47519, B1 => n42284, B2 => 
                           n47511, ZN => n36206);
   U526 : OAI22_X1 port map( A1 => n40647, A2 => n47514, B1 => n42283, B2 => 
                           n47567, ZN => n36207);
   U527 : OAI22_X1 port map( A1 => n40637, A2 => n47515, B1 => n42282, B2 => 
                           n47511, ZN => n36208);
   U528 : OAI22_X1 port map( A1 => n40647, A2 => n47516, B1 => n42281, B2 => 
                           n47567, ZN => n36209);
   U529 : OAI22_X1 port map( A1 => n40647, A2 => n47517, B1 => n42280, B2 => 
                           n47567, ZN => n36210);
   U530 : OAI22_X1 port map( A1 => n40642, A2 => n47517, B1 => n42279, B2 => 
                           n47561, ZN => n36211);
   U531 : OAI22_X1 port map( A1 => n40646, A2 => n47515, B1 => n42278, B2 => 
                           n47562, ZN => n36212);
   U532 : OAI22_X1 port map( A1 => n40642, A2 => n47515, B1 => n42277, B2 => 
                           n47561, ZN => n36213);
   U533 : OAI22_X1 port map( A1 => n40637, A2 => n47516, B1 => n42276, B2 => 
                           n47511, ZN => n36214);
   U534 : OAI22_X1 port map( A1 => n40628, A2 => n47516, B1 => n42275, B2 => 
                           n47512, ZN => n36215);
   U535 : OAI22_X1 port map( A1 => n40646, A2 => n47517, B1 => n42274, B2 => 
                           n47562, ZN => n36216);
   U536 : OAI22_X1 port map( A1 => n40642, A2 => n47534, B1 => n42273, B2 => 
                           n47561, ZN => n36217);
   U537 : OAI22_X1 port map( A1 => n40647, A2 => n47515, B1 => n42272, B2 => 
                           n47567, ZN => n36218);
   U538 : OAI22_X1 port map( A1 => n40646, A2 => n47529, B1 => n42271, B2 => 
                           n47562, ZN => n36219);
   U539 : OAI22_X1 port map( A1 => n40628, A2 => n47517, B1 => n42270, B2 => 
                           n47512, ZN => n36220);
   U540 : OAI22_X1 port map( A1 => n40646, A2 => n47516, B1 => n42269, B2 => 
                           n47562, ZN => n36221);
   U541 : OAI22_X1 port map( A1 => n40646, A2 => n47514, B1 => n42268, B2 => 
                           n47562, ZN => n36222);
   U542 : OAI22_X1 port map( A1 => n40646, A2 => n47518, B1 => n42267, B2 => 
                           n47562, ZN => n36223);
   U543 : OAI22_X1 port map( A1 => n40642, A2 => n47516, B1 => n42266, B2 => 
                           n47561, ZN => n36224);
   U544 : OAI22_X1 port map( A1 => n40638, A2 => n47537, B1 => n42265, B2 => 
                           n47563, ZN => n36225);
   U545 : OAI22_X1 port map( A1 => n40605, A2 => n47537, B1 => n42264, B2 => 
                           n47565, ZN => n36226);
   U546 : OAI22_X1 port map( A1 => n40638, A2 => n47516, B1 => n42263, B2 => 
                           n47563, ZN => n36227);
   U547 : OAI22_X1 port map( A1 => n40638, A2 => n47518, B1 => n42262, B2 => 
                           n47563, ZN => n36228);
   U548 : OAI22_X1 port map( A1 => n40628, A2 => n47529, B1 => n42261, B2 => 
                           n47512, ZN => n36229);
   U549 : OAI22_X1 port map( A1 => n40628, A2 => n47526, B1 => n42260, B2 => 
                           n47512, ZN => n36230);
   U550 : OAI22_X1 port map( A1 => n40646, A2 => n47549, B1 => n42259, B2 => 
                           n47562, ZN => n36231);
   U551 : OAI22_X1 port map( A1 => n40642, A2 => n47530, B1 => n42258, B2 => 
                           n47561, ZN => n36232);
   U552 : OAI22_X1 port map( A1 => n40638, A2 => n47530, B1 => n42257, B2 => 
                           n47563, ZN => n36233);
   U553 : OAI22_X1 port map( A1 => n40604, A2 => n47534, B1 => n42256, B2 => 
                           n47566, ZN => n36234);
   U554 : OAI22_X1 port map( A1 => n40637, A2 => n47530, B1 => n42255, B2 => 
                           n47511, ZN => n36235);
   U555 : OAI22_X1 port map( A1 => n40604, A2 => n47525, B1 => n42254, B2 => 
                           n47566, ZN => n36236);
   U556 : OAI22_X1 port map( A1 => n40605, A2 => n47525, B1 => n42253, B2 => 
                           n47565, ZN => n36237);
   U557 : OAI22_X1 port map( A1 => n40646, A2 => n47526, B1 => n42252, B2 => 
                           n47562, ZN => n36238);
   U558 : OAI22_X1 port map( A1 => n40642, A2 => n47526, B1 => n42251, B2 => 
                           n47561, ZN => n36239);
   U559 : OAI22_X1 port map( A1 => n40647, A2 => n47518, B1 => n42250, B2 => 
                           n47567, ZN => n36240);
   U560 : OAI22_X1 port map( A1 => n40628, A2 => n47549, B1 => n42249, B2 => 
                           n47512, ZN => n36241);
   U561 : OAI22_X1 port map( A1 => n40642, A2 => n47529, B1 => n42248, B2 => 
                           n47561, ZN => n36242);
   U562 : OAI22_X1 port map( A1 => n40637, A2 => n47529, B1 => n42247, B2 => 
                           n47511, ZN => n36243);
   U563 : OAI22_X1 port map( A1 => n40638, A2 => n47526, B1 => n42246, B2 => 
                           n47563, ZN => n36244);
   U564 : OAI22_X1 port map( A1 => n40637, A2 => n47514, B1 => n42245, B2 => 
                           n47511, ZN => n36245);
   U565 : OAI22_X1 port map( A1 => n40638, A2 => n47514, B1 => n42244, B2 => 
                           n47563, ZN => n36246);
   U566 : OAI22_X1 port map( A1 => n40642, A2 => n47514, B1 => n42243, B2 => 
                           n47561, ZN => n36247);
   U567 : OAI22_X1 port map( A1 => n40637, A2 => n47526, B1 => n42242, B2 => 
                           n47511, ZN => n36248);
   U568 : OAI22_X1 port map( A1 => n40628, A2 => n47518, B1 => n42241, B2 => 
                           n47512, ZN => n36249);
   U569 : OAI22_X1 port map( A1 => n40642, A2 => n47518, B1 => n42240, B2 => 
                           n47561, ZN => n36250);
   U570 : OAI22_X1 port map( A1 => n40605, A2 => n47534, B1 => n42239, B2 => 
                           n47565, ZN => n36251);
   U571 : OAI22_X1 port map( A1 => n40646, A2 => n47530, B1 => n42238, B2 => 
                           n47562, ZN => n36252);
   U572 : OAI22_X1 port map( A1 => n40628, A2 => n47530, B1 => n42237, B2 => 
                           n47512, ZN => n36253);
   U573 : OAI22_X1 port map( A1 => n40604, A2 => n47521, B1 => n42236, B2 => 
                           n47566, ZN => n36254);
   U574 : OAI22_X1 port map( A1 => n40637, A2 => n47518, B1 => n42235, B2 => 
                           n47511, ZN => n36255);
   U575 : OAI22_X1 port map( A1 => n40628, A2 => n47514, B1 => n42234, B2 => 
                           n47512, ZN => n36256);
   U576 : OAI22_X1 port map( A1 => n40638, A2 => n47534, B1 => n42233, B2 => 
                           n47563, ZN => n36257);
   U577 : OAI22_X1 port map( A1 => n40638, A2 => n47529, B1 => n42232, B2 => 
                           n47563, ZN => n36258);
   U578 : OAI22_X1 port map( A1 => n40623, A2 => n47520, B1 => n42231, B2 => 
                           n47535, ZN => n36259);
   U579 : OAI22_X1 port map( A1 => n40623, A2 => n47528, B1 => n42230, B2 => 
                           n47535, ZN => n36260);
   U580 : OAI22_X1 port map( A1 => n40623, A2 => n47529, B1 => n42229, B2 => 
                           n47535, ZN => n36261);
   U581 : OAI22_X1 port map( A1 => n40623, A2 => n47530, B1 => n42228, B2 => 
                           n47535, ZN => n36262);
   U582 : OAI22_X1 port map( A1 => n40623, A2 => n47549, B1 => n42227, B2 => 
                           n47535, ZN => n36263);
   U583 : OAI22_X1 port map( A1 => n40623, A2 => n47525, B1 => n42226, B2 => 
                           n47535, ZN => n36264);
   U584 : OAI22_X1 port map( A1 => n40623, A2 => n47521, B1 => n42225, B2 => 
                           n47535, ZN => n36265);
   U585 : OAI22_X1 port map( A1 => n40614, A2 => n47513, B1 => n42224, B2 => 
                           n47536, ZN => n36266);
   U586 : OAI22_X1 port map( A1 => n40623, A2 => n47513, B1 => n42223, B2 => 
                           n47535, ZN => n36267);
   U587 : OAI22_X1 port map( A1 => n40617, A2 => n47514, B1 => n42222, B2 => 
                           n47538, ZN => n36268);
   U588 : OAI22_X1 port map( A1 => n40610, A2 => n47513, B1 => n42221, B2 => 
                           n47540, ZN => n36269);
   U589 : OAI22_X1 port map( A1 => n40611, A2 => n47513, B1 => n42220, B2 => 
                           n47543, ZN => n36270);
   U590 : OAI22_X1 port map( A1 => n40619, A2 => n47515, B1 => n42219, B2 => 
                           n47541, ZN => n36271);
   U591 : OAI22_X1 port map( A1 => n40619, A2 => n47516, B1 => n42218, B2 => 
                           n47541, ZN => n36272);
   U592 : OAI22_X1 port map( A1 => n40610, A2 => n47514, B1 => n42217, B2 => 
                           n47540, ZN => n36273);
   U593 : OAI22_X1 port map( A1 => n40611, A2 => n47517, B1 => n42216, B2 => 
                           n47543, ZN => n36274);
   U594 : OAI22_X1 port map( A1 => n40613, A2 => n47517, B1 => n42215, B2 => 
                           n47532, ZN => n36275);
   U595 : OAI22_X1 port map( A1 => n40613, A2 => n47513, B1 => n42214, B2 => 
                           n47532, ZN => n36276);
   U596 : OAI22_X1 port map( A1 => n40614, A2 => n47517, B1 => n42213, B2 => 
                           n47536, ZN => n36277);
   U597 : OAI22_X1 port map( A1 => n40610, A2 => n47517, B1 => n42212, B2 => 
                           n47540, ZN => n36278);
   U598 : OAI22_X1 port map( A1 => n40623, A2 => n47514, B1 => n42211, B2 => 
                           n47535, ZN => n36279);
   U599 : OAI22_X1 port map( A1 => n40619, A2 => n47514, B1 => n42210, B2 => 
                           n47541, ZN => n36281);
   U600 : OAI22_X1 port map( A1 => n40617, A2 => n47517, B1 => n42209, B2 => 
                           n47538, ZN => n36283);
   U601 : OAI22_X1 port map( A1 => n40619, A2 => n47518, B1 => n42208, B2 => 
                           n47541, ZN => n36284);
   U602 : OAI22_X1 port map( A1 => n40619, A2 => n47513, B1 => n42207, B2 => 
                           n47541, ZN => n36285);
   U603 : OAI22_X1 port map( A1 => n40611, A2 => n47514, B1 => n42206, B2 => 
                           n47543, ZN => n36286);
   U604 : OAI22_X1 port map( A1 => n40614, A2 => n47514, B1 => n42205, B2 => 
                           n47536, ZN => n36287);
   U605 : OAI22_X1 port map( A1 => n40621, A2 => n47521, B1 => n42204, B2 => 
                           n47539, ZN => n36288);
   U606 : OAI22_X1 port map( A1 => n40614, A2 => n47518, B1 => n42203, B2 => 
                           n47536, ZN => n36289);
   U607 : OAI22_X1 port map( A1 => n40614, A2 => n47515, B1 => n42202, B2 => 
                           n47536, ZN => n36290);
   U608 : OAI22_X1 port map( A1 => n40613, A2 => n47514, B1 => n42201, B2 => 
                           n47532, ZN => n36291);
   U609 : OAI22_X1 port map( A1 => n40621, A2 => n47534, B1 => n42200, B2 => 
                           n47539, ZN => n36292);
   U610 : OAI22_X1 port map( A1 => n40636, A2 => n47521, B1 => n42199, B2 => 
                           n47542, ZN => n36293);
   U611 : OAI22_X1 port map( A1 => n40611, A2 => n47518, B1 => n42198, B2 => 
                           n47543, ZN => n36294);
   U612 : OAI22_X1 port map( A1 => n40636, A2 => n47534, B1 => n42197, B2 => 
                           n47542, ZN => n36295);
   U613 : OAI22_X1 port map( A1 => n40617, A2 => n47513, B1 => n42196, B2 => 
                           n47538, ZN => n36297);
   U614 : OAI22_X1 port map( A1 => n40614, A2 => n47516, B1 => n42195, B2 => 
                           n47536, ZN => n36298);
   U615 : OAI22_X1 port map( A1 => n40610, A2 => n47518, B1 => n42194, B2 => 
                           n47540, ZN => n36299);
   U616 : OAI22_X1 port map( A1 => n40617, A2 => n47518, B1 => n42193, B2 => 
                           n47538, ZN => n36300);
   U617 : OAI22_X1 port map( A1 => n40617, A2 => n47519, B1 => n42192, B2 => 
                           n47538, ZN => n36301);
   U618 : OAI22_X1 port map( A1 => n40614, A2 => n47519, B1 => n42191, B2 => 
                           n47536, ZN => n36302);
   U619 : OAI22_X1 port map( A1 => n40623, A2 => n47518, B1 => n42190, B2 => 
                           n47535, ZN => n36304);
   U620 : OAI22_X1 port map( A1 => n40623, A2 => n47515, B1 => n42189, B2 => 
                           n47535, ZN => n36305);
   U621 : OAI22_X1 port map( A1 => n40623, A2 => n47516, B1 => n42188, B2 => 
                           n47535, ZN => n36306);
   U622 : OAI22_X1 port map( A1 => n40623, A2 => n47517, B1 => n42187, B2 => 
                           n47535, ZN => n36307);
   U623 : OAI22_X1 port map( A1 => n40623, A2 => n47519, B1 => n42186, B2 => 
                           n47535, ZN => n36308);
   U624 : OAI22_X1 port map( A1 => n40636, A2 => n47525, B1 => n42185, B2 => 
                           n47542, ZN => n36309);
   U625 : OAI22_X1 port map( A1 => n40636, A2 => n47513, B1 => n42184, B2 => 
                           n47542, ZN => n36310);
   U626 : OAI22_X1 port map( A1 => n40613, A2 => n47518, B1 => n42183, B2 => 
                           n47532, ZN => n36311);
   U627 : OAI22_X1 port map( A1 => n40610, A2 => n47515, B1 => n42182, B2 => 
                           n47540, ZN => n36312);
   U628 : OAI22_X1 port map( A1 => n40617, A2 => n47515, B1 => n42181, B2 => 
                           n47538, ZN => n36313);
   U629 : OAI22_X1 port map( A1 => n40613, A2 => n47515, B1 => n42180, B2 => 
                           n47532, ZN => n36314);
   U630 : OAI22_X1 port map( A1 => n40611, A2 => n47515, B1 => n42179, B2 => 
                           n47543, ZN => n36316);
   U631 : OAI22_X1 port map( A1 => n40613, A2 => n47516, B1 => n42178, B2 => 
                           n47532, ZN => n36317);
   U632 : OAI22_X1 port map( A1 => n40611, A2 => n47516, B1 => n42177, B2 => 
                           n47543, ZN => n36318);
   U633 : OAI22_X1 port map( A1 => n40613, A2 => n47519, B1 => n42176, B2 => 
                           n47532, ZN => n36319);
   U634 : OAI22_X1 port map( A1 => n40611, A2 => n47519, B1 => n42175, B2 => 
                           n47543, ZN => n36320);
   U635 : OAI22_X1 port map( A1 => n40610, A2 => n47519, B1 => n42174, B2 => 
                           n47540, ZN => n36322);
   U636 : OAI22_X1 port map( A1 => n40610, A2 => n47516, B1 => n42173, B2 => 
                           n47540, ZN => n36323);
   U637 : OAI22_X1 port map( A1 => n40617, A2 => n47516, B1 => n42172, B2 => 
                           n47538, ZN => n36324);
   U638 : OAI22_X1 port map( A1 => n40619, A2 => n47517, B1 => n42171, B2 => 
                           n47541, ZN => n36325);
   U639 : OAI22_X1 port map( A1 => n40619, A2 => n47519, B1 => n42170, B2 => 
                           n47541, ZN => n36326);
   U640 : OAI22_X1 port map( A1 => n40621, A2 => n47516, B1 => n42169, B2 => 
                           n47539, ZN => n36328);
   U641 : OAI22_X1 port map( A1 => n40621, A2 => n47517, B1 => n42168, B2 => 
                           n47539, ZN => n36329);
   U642 : OAI22_X1 port map( A1 => n40621, A2 => n47519, B1 => n42167, B2 => 
                           n47539, ZN => n36330);
   U643 : OAI22_X1 port map( A1 => n40636, A2 => n47555, B1 => n42166, B2 => 
                           n47542, ZN => n36331);
   U644 : OAI22_X1 port map( A1 => n40621, A2 => n47518, B1 => n42165, B2 => 
                           n47539, ZN => n36332);
   U645 : OAI22_X1 port map( A1 => n40621, A2 => n47515, B1 => n42164, B2 => 
                           n47539, ZN => n36333);
   U646 : OAI22_X1 port map( A1 => n40621, A2 => n47513, B1 => n42163, B2 => 
                           n47539, ZN => n36334);
   U647 : OAI22_X1 port map( A1 => n40617, A2 => n47531, B1 => n42162, B2 => 
                           n47538, ZN => n36335);
   U648 : OAI22_X1 port map( A1 => n40621, A2 => n47514, B1 => n42161, B2 => 
                           n47539, ZN => n36336);
   U649 : OAI22_X1 port map( A1 => n40613, A2 => n47537, B1 => n42160, B2 => 
                           n47532, ZN => n36337);
   U650 : OAI22_X1 port map( A1 => n40617, A2 => n47528, B1 => n42159, B2 => 
                           n47538, ZN => n36338);
   U651 : OAI22_X1 port map( A1 => n40617, A2 => n47520, B1 => n42158, B2 => 
                           n47538, ZN => n36339);
   U652 : OAI22_X1 port map( A1 => n40617, A2 => n47522, B1 => n42157, B2 => 
                           n47538, ZN => n36340);
   U653 : OAI22_X1 port map( A1 => n40617, A2 => n47529, B1 => n42156, B2 => 
                           n47538, ZN => n36341);
   U654 : OAI22_X1 port map( A1 => n40617, A2 => n47530, B1 => n42155, B2 => 
                           n47538, ZN => n36342);
   U655 : CLKBUF_X1 port map( A => n47549, Z => n47564);
   U656 : OAI22_X1 port map( A1 => n40617, A2 => n47564, B1 => n42154, B2 => 
                           n47538, ZN => n36343);
   U657 : OAI22_X1 port map( A1 => n40617, A2 => n47525, B1 => n42153, B2 => 
                           n47538, ZN => n36344);
   U658 : OAI22_X1 port map( A1 => n40617, A2 => n47526, B1 => n42152, B2 => 
                           n47538, ZN => n36345);
   U659 : OAI22_X1 port map( A1 => n40617, A2 => n47521, B1 => n42151, B2 => 
                           n47538, ZN => n36346);
   U660 : OAI22_X1 port map( A1 => n40617, A2 => n47534, B1 => n42150, B2 => 
                           n47538, ZN => n36347);
   U661 : OAI22_X1 port map( A1 => n40610, A2 => n47522, B1 => n42149, B2 => 
                           n47540, ZN => n36348);
   U662 : OAI22_X1 port map( A1 => n40611, A2 => n47522, B1 => n42148, B2 => 
                           n47543, ZN => n36349);
   U663 : OAI22_X1 port map( A1 => n40617, A2 => n47523, B1 => n42147, B2 => 
                           n47538, ZN => n36350);
   U664 : OAI22_X1 port map( A1 => n40614, A2 => n47522, B1 => n42146, B2 => 
                           n47536, ZN => n36351);
   U665 : OAI22_X1 port map( A1 => n40619, A2 => n47522, B1 => n42145, B2 => 
                           n47541, ZN => n36352);
   U666 : OAI22_X1 port map( A1 => n40613, A2 => n47522, B1 => n42144, B2 => 
                           n47532, ZN => n36353);
   U667 : OAI22_X1 port map( A1 => n40621, A2 => n47522, B1 => n42143, B2 => 
                           n47539, ZN => n36354);
   U668 : OAI22_X1 port map( A1 => n40623, A2 => n47522, B1 => n42142, B2 => 
                           n47535, ZN => n36355);
   U669 : OAI22_X1 port map( A1 => n40619, A2 => n47523, B1 => n42141, B2 => 
                           n47541, ZN => n36356);
   U670 : OAI22_X1 port map( A1 => n40621, A2 => n47523, B1 => n42140, B2 => 
                           n47539, ZN => n36357);
   U671 : OAI22_X1 port map( A1 => n40623, A2 => n47523, B1 => n42139, B2 => 
                           n47535, ZN => n36358);
   U672 : OAI22_X1 port map( A1 => n40610, A2 => n47523, B1 => n42138, B2 => 
                           n47540, ZN => n36359);
   U673 : OAI22_X1 port map( A1 => n40611, A2 => n47523, B1 => n42137, B2 => 
                           n47543, ZN => n36360);
   U674 : OAI22_X1 port map( A1 => n40613, A2 => n47523, B1 => n42136, B2 => 
                           n47532, ZN => n36361);
   U675 : OAI22_X1 port map( A1 => n40614, A2 => n47523, B1 => n42135, B2 => 
                           n47536, ZN => n36362);
   U676 : OAI22_X1 port map( A1 => n40617, A2 => n47524, B1 => n42134, B2 => 
                           n47538, ZN => n36363);
   U677 : OAI22_X1 port map( A1 => n40621, A2 => n47525, B1 => n42133, B2 => 
                           n47539, ZN => n36364);
   U678 : OAI22_X1 port map( A1 => n40619, A2 => n47526, B1 => n42132, B2 => 
                           n47541, ZN => n36365);
   U679 : OAI22_X1 port map( A1 => n40621, A2 => n47526, B1 => n42131, B2 => 
                           n47539, ZN => n36366);
   U680 : OAI22_X1 port map( A1 => n40623, A2 => n47526, B1 => n42130, B2 => 
                           n47535, ZN => n36367);
   U681 : OAI22_X1 port map( A1 => n40610, A2 => n47526, B1 => n42129, B2 => 
                           n47540, ZN => n36368);
   U682 : OAI22_X1 port map( A1 => n40611, A2 => n47526, B1 => n42128, B2 => 
                           n47543, ZN => n36369);
   U683 : OAI22_X1 port map( A1 => n40613, A2 => n47526, B1 => n42127, B2 => 
                           n47532, ZN => n36370);
   U684 : OAI22_X1 port map( A1 => n40614, A2 => n47526, B1 => n42126, B2 => 
                           n47536, ZN => n36371);
   U685 : OAI22_X1 port map( A1 => n40621, A2 => n47555, B1 => n42125, B2 => 
                           n47539, ZN => n36372);
   U686 : OAI22_X1 port map( A1 => n40621, A2 => n47533, B1 => n42124, B2 => 
                           n47539, ZN => n36373);
   U687 : OAI22_X1 port map( A1 => n40621, A2 => n47527, B1 => n42123, B2 => 
                           n47539, ZN => n36374);
   U688 : OAI22_X1 port map( A1 => n40621, A2 => n47524, B1 => n42122, B2 => 
                           n47539, ZN => n36375);
   U689 : OAI22_X1 port map( A1 => n40621, A2 => n47531, B1 => n42121, B2 => 
                           n47539, ZN => n36376);
   U690 : OAI22_X1 port map( A1 => n40621, A2 => n47520, B1 => n42120, B2 => 
                           n47539, ZN => n36377);
   U691 : OAI22_X1 port map( A1 => n40621, A2 => n47528, B1 => n42119, B2 => 
                           n47539, ZN => n36378);
   U692 : OAI22_X1 port map( A1 => n40621, A2 => n47529, B1 => n42118, B2 => 
                           n47539, ZN => n36379);
   U693 : OAI22_X1 port map( A1 => n40621, A2 => n47530, B1 => n42117, B2 => 
                           n47539, ZN => n36380);
   U694 : OAI22_X1 port map( A1 => n40621, A2 => n47564, B1 => n42116, B2 => 
                           n47539, ZN => n36381);
   U695 : OAI22_X1 port map( A1 => n40623, A2 => n47527, B1 => n42115, B2 => 
                           n47535, ZN => n36382);
   U696 : OAI22_X1 port map( A1 => n40623, A2 => n47533, B1 => n42114, B2 => 
                           n47535, ZN => n36383);
   U697 : OAI22_X1 port map( A1 => n40623, A2 => n47555, B1 => n42113, B2 => 
                           n47535, ZN => n36384);
   U698 : OAI22_X1 port map( A1 => n40623, A2 => n47524, B1 => n42112, B2 => 
                           n47535, ZN => n36385);
   U699 : OAI22_X1 port map( A1 => n40623, A2 => n47531, B1 => n42111, B2 => 
                           n47535, ZN => n36386);
   U700 : OAI22_X1 port map( A1 => n40619, A2 => n47534, B1 => n42110, B2 => 
                           n47541, ZN => n36387);
   U701 : OAI22_X1 port map( A1 => n40613, A2 => n47527, B1 => n42109, B2 => 
                           n47532, ZN => n36388);
   U702 : OAI22_X1 port map( A1 => n40613, A2 => n47533, B1 => n42108, B2 => 
                           n47532, ZN => n36389);
   U703 : OAI22_X1 port map( A1 => n40610, A2 => n47524, B1 => n42107, B2 => 
                           n47540, ZN => n36390);
   U704 : OAI22_X1 port map( A1 => n40611, A2 => n47524, B1 => n42106, B2 => 
                           n47543, ZN => n36391);
   U705 : OAI22_X1 port map( A1 => n40613, A2 => n47524, B1 => n42105, B2 => 
                           n47532, ZN => n36392);
   U706 : OAI22_X1 port map( A1 => n40614, A2 => n47524, B1 => n42104, B2 => 
                           n47536, ZN => n36393);
   U707 : OAI22_X1 port map( A1 => n40613, A2 => n47531, B1 => n42103, B2 => 
                           n47532, ZN => n36394);
   U708 : OAI22_X1 port map( A1 => n40613, A2 => n47520, B1 => n42102, B2 => 
                           n47532, ZN => n36395);
   U709 : OAI22_X1 port map( A1 => n40613, A2 => n47528, B1 => n42101, B2 => 
                           n47532, ZN => n36396);
   U710 : OAI22_X1 port map( A1 => n40613, A2 => n47529, B1 => n42100, B2 => 
                           n47532, ZN => n36397);
   U711 : OAI22_X1 port map( A1 => n40636, A2 => n47523, B1 => n42099, B2 => 
                           n47542, ZN => n36399);
   U712 : OAI22_X1 port map( A1 => n40613, A2 => n47530, B1 => n42098, B2 => 
                           n47532, ZN => n36400);
   U713 : OAI22_X1 port map( A1 => n40613, A2 => n47549, B1 => n42097, B2 => 
                           n47532, ZN => n36401);
   U714 : OAI22_X1 port map( A1 => n40613, A2 => n47525, B1 => n42096, B2 => 
                           n47532, ZN => n36402);
   U715 : OAI22_X1 port map( A1 => n40636, A2 => n47517, B1 => n42095, B2 => 
                           n47542, ZN => n36404);
   U716 : OAI22_X1 port map( A1 => n40613, A2 => n47555, B1 => n42094, B2 => 
                           n47532, ZN => n36405);
   U717 : OAI22_X1 port map( A1 => n40613, A2 => n47521, B1 => n42093, B2 => 
                           n47532, ZN => n36406);
   U718 : OAI22_X1 port map( A1 => n40610, A2 => n47531, B1 => n42092, B2 => 
                           n47540, ZN => n36407);
   U719 : OAI22_X1 port map( A1 => n40611, A2 => n47531, B1 => n42091, B2 => 
                           n47543, ZN => n36408);
   U720 : OAI22_X1 port map( A1 => n40614, A2 => n47531, B1 => n42090, B2 => 
                           n47536, ZN => n36409);
   U721 : OAI22_X1 port map( A1 => n40613, A2 => n47534, B1 => n42089, B2 => 
                           n47532, ZN => n36410);
   U722 : OAI22_X1 port map( A1 => n40610, A2 => n47520, B1 => n42088, B2 => 
                           n47540, ZN => n36411);
   U723 : OAI22_X1 port map( A1 => n40611, A2 => n47555, B1 => n42087, B2 => 
                           n47543, ZN => n36412);
   U724 : OAI22_X1 port map( A1 => n40611, A2 => n47520, B1 => n42086, B2 => 
                           n47543, ZN => n36413);
   U725 : OAI22_X1 port map( A1 => n40610, A2 => n47555, B1 => n42085, B2 => 
                           n47540, ZN => n36414);
   U726 : OAI22_X1 port map( A1 => n40610, A2 => n47533, B1 => n42084, B2 => 
                           n47540, ZN => n36415);
   U727 : OAI22_X1 port map( A1 => n40614, A2 => n47520, B1 => n42083, B2 => 
                           n47536, ZN => n36416);
   U728 : OAI22_X1 port map( A1 => n40614, A2 => n47527, B1 => n42082, B2 => 
                           n47536, ZN => n36417);
   U729 : OAI22_X1 port map( A1 => n40614, A2 => n47533, B1 => n42081, B2 => 
                           n47536, ZN => n36418);
   U730 : OAI22_X1 port map( A1 => n40614, A2 => n47528, B1 => n42080, B2 => 
                           n47536, ZN => n36419);
   U731 : OAI22_X1 port map( A1 => n40619, A2 => n47527, B1 => n42079, B2 => 
                           n47541, ZN => n36421);
   U732 : OAI22_X1 port map( A1 => n40619, A2 => n47533, B1 => n42078, B2 => 
                           n47541, ZN => n36423);
   U733 : OAI22_X1 port map( A1 => n40619, A2 => n47555, B1 => n42077, B2 => 
                           n47541, ZN => n36424);
   U734 : OAI22_X1 port map( A1 => n40636, A2 => n47519, B1 => n42076, B2 => 
                           n47542, ZN => n36426);
   U735 : OAI22_X1 port map( A1 => n40619, A2 => n47524, B1 => n42075, B2 => 
                           n47541, ZN => n36428);
   U736 : OAI22_X1 port map( A1 => n40619, A2 => n47531, B1 => n42074, B2 => 
                           n47541, ZN => n36430);
   U737 : OAI22_X1 port map( A1 => n40619, A2 => n47520, B1 => n42073, B2 => 
                           n47541, ZN => n36432);
   U738 : OAI22_X1 port map( A1 => n40619, A2 => n47528, B1 => n42072, B2 => 
                           n47541, ZN => n36434);
   U739 : OAI22_X1 port map( A1 => n40614, A2 => n47529, B1 => n42071, B2 => 
                           n47536, ZN => n36435);
   U740 : OAI22_X1 port map( A1 => n40610, A2 => n47529, B1 => n42070, B2 => 
                           n47540, ZN => n36436);
   U741 : OAI22_X1 port map( A1 => n40619, A2 => n47529, B1 => n42069, B2 => 
                           n47541, ZN => n36437);
   U742 : OAI22_X1 port map( A1 => n40619, A2 => n47530, B1 => n42068, B2 => 
                           n47541, ZN => n36438);
   U743 : OAI22_X1 port map( A1 => n40611, A2 => n47529, B1 => n42067, B2 => 
                           n47543, ZN => n36439);
   U744 : OAI22_X1 port map( A1 => n40617, A2 => n47555, B1 => n42066, B2 => 
                           n47538, ZN => n36440);
   U745 : OAI22_X1 port map( A1 => n40636, A2 => n47515, B1 => n42065, B2 => 
                           n47542, ZN => n36442);
   U746 : OAI22_X1 port map( A1 => n40636, A2 => n47533, B1 => n42064, B2 => 
                           n47542, ZN => n36443);
   U747 : OAI22_X1 port map( A1 => n40611, A2 => n47533, B1 => n42063, B2 => 
                           n47543, ZN => n36444);
   U748 : OAI22_X1 port map( A1 => n40617, A2 => n47533, B1 => n42062, B2 => 
                           n47538, ZN => n36445);
   U749 : OAI22_X1 port map( A1 => n40611, A2 => n47527, B1 => n42061, B2 => 
                           n47543, ZN => n36446);
   U750 : OAI22_X1 port map( A1 => n40610, A2 => n47527, B1 => n42060, B2 => 
                           n47540, ZN => n36447);
   U751 : OAI22_X1 port map( A1 => n40614, A2 => n47555, B1 => n42059, B2 => 
                           n47536, ZN => n36448);
   U752 : OAI22_X1 port map( A1 => n40636, A2 => n47529, B1 => n42058, B2 => 
                           n47542, ZN => n36450);
   U753 : OAI22_X1 port map( A1 => n40636, A2 => n47527, B1 => n42057, B2 => 
                           n47542, ZN => n36451);
   U754 : OAI22_X1 port map( A1 => n40611, A2 => n47534, B1 => n42056, B2 => 
                           n47543, ZN => n36452);
   U755 : OAI22_X1 port map( A1 => n40611, A2 => n47521, B1 => n42055, B2 => 
                           n47543, ZN => n36453);
   U756 : OAI22_X1 port map( A1 => n40636, A2 => n47514, B1 => n42054, B2 => 
                           n47542, ZN => n36455);
   U757 : OAI22_X1 port map( A1 => n40636, A2 => n47528, B1 => n42053, B2 => 
                           n47542, ZN => n36456);
   U758 : OAI22_X1 port map( A1 => n40617, A2 => n47527, B1 => n42052, B2 => 
                           n47538, ZN => n36458);
   U759 : OAI22_X1 port map( A1 => n40619, A2 => n47564, B1 => n42051, B2 => 
                           n47541, ZN => n36459);
   U760 : OAI22_X1 port map( A1 => n40611, A2 => n47530, B1 => n42050, B2 => 
                           n47543, ZN => n36460);
   U761 : OAI22_X1 port map( A1 => n40619, A2 => n47525, B1 => n42049, B2 => 
                           n47541, ZN => n36461);
   U762 : OAI22_X1 port map( A1 => n40614, A2 => n47525, B1 => n42048, B2 => 
                           n47536, ZN => n36462);
   U763 : OAI22_X1 port map( A1 => n40611, A2 => n47525, B1 => n42047, B2 => 
                           n47543, ZN => n36463);
   U764 : OAI22_X1 port map( A1 => n40611, A2 => n47549, B1 => n42046, B2 => 
                           n47543, ZN => n36464);
   U765 : OAI22_X1 port map( A1 => n40636, A2 => n47520, B1 => n42045, B2 => 
                           n47542, ZN => n36465);
   U766 : OAI22_X1 port map( A1 => n40610, A2 => n47549, B1 => n42044, B2 => 
                           n47540, ZN => n36466);
   U767 : OAI22_X1 port map( A1 => n40611, A2 => n47528, B1 => n42043, B2 => 
                           n47543, ZN => n36467);
   U768 : OAI22_X1 port map( A1 => n40610, A2 => n47534, B1 => n42042, B2 => 
                           n47540, ZN => n36468);
   U769 : OAI22_X1 port map( A1 => n40636, A2 => n47518, B1 => n42041, B2 => 
                           n47542, ZN => n36470);
   U770 : OAI22_X1 port map( A1 => n40610, A2 => n47521, B1 => n42040, B2 => 
                           n47540, ZN => n36471);
   U771 : OAI22_X1 port map( A1 => n40610, A2 => n47525, B1 => n42039, B2 => 
                           n47540, ZN => n36473);
   U772 : OAI22_X1 port map( A1 => n40636, A2 => n47531, B1 => n42038, B2 => 
                           n47542, ZN => n36474);
   U773 : OAI22_X1 port map( A1 => n40614, A2 => n47521, B1 => n42037, B2 => 
                           n47536, ZN => n36475);
   U774 : OAI22_X1 port map( A1 => n40610, A2 => n47528, B1 => n42036, B2 => 
                           n47540, ZN => n36476);
   U775 : OAI22_X1 port map( A1 => n40636, A2 => n47526, B1 => n42035, B2 => 
                           n47542, ZN => n36478);
   U776 : OAI22_X1 port map( A1 => n40614, A2 => n47530, B1 => n42034, B2 => 
                           n47536, ZN => n36479);
   U777 : OAI22_X1 port map( A1 => n40636, A2 => n47549, B1 => n42033, B2 => 
                           n47542, ZN => n36480);
   U778 : OAI22_X1 port map( A1 => n40614, A2 => n47534, B1 => n42032, B2 => 
                           n47536, ZN => n36481);
   U779 : OAI22_X1 port map( A1 => n40610, A2 => n47530, B1 => n42031, B2 => 
                           n47540, ZN => n36482);
   U780 : OAI22_X1 port map( A1 => n40636, A2 => n47530, B1 => n42030, B2 => 
                           n47542, ZN => n36483);
   U781 : OAI22_X1 port map( A1 => n40636, A2 => n47522, B1 => n42029, B2 => 
                           n47542, ZN => n36484);
   U782 : OAI22_X1 port map( A1 => n40636, A2 => n47524, B1 => n42028, B2 => 
                           n47542, ZN => n36486);
   U783 : OAI22_X1 port map( A1 => n40619, A2 => n47521, B1 => n42027, B2 => 
                           n47541, ZN => n36488);
   U784 : OAI22_X1 port map( A1 => n40636, A2 => n47516, B1 => n42026, B2 => 
                           n47542, ZN => n36490);
   U785 : OAI22_X1 port map( A1 => n40623, A2 => n47534, B1 => n42025, B2 => 
                           n47535, ZN => n36491);
   U786 : OAI22_X1 port map( A1 => n40614, A2 => n47549, B1 => n42024, B2 => 
                           n47536, ZN => n36492);
   U787 : OAI22_X1 port map( A1 => n40623, A2 => n47537, B1 => n42023, B2 => 
                           n47535, ZN => n36494);
   U788 : OAI22_X1 port map( A1 => n40614, A2 => n47537, B1 => n42022, B2 => 
                           n47536, ZN => n36495);
   U789 : OAI22_X1 port map( A1 => n40617, A2 => n47537, B1 => n42021, B2 => 
                           n47538, ZN => n36496);
   U790 : OAI22_X1 port map( A1 => n40621, A2 => n47537, B1 => n42020, B2 => 
                           n47539, ZN => n36497);
   U791 : OAI22_X1 port map( A1 => n40610, A2 => n47537, B1 => n42019, B2 => 
                           n47540, ZN => n36498);
   U792 : OAI22_X1 port map( A1 => n40604, A2 => n47537, B1 => n42018, B2 => 
                           n47566, ZN => n36499);
   U793 : OAI22_X1 port map( A1 => n40619, A2 => n47537, B1 => n42017, B2 => 
                           n47541, ZN => n36500);
   U794 : OAI22_X1 port map( A1 => n40636, A2 => n47537, B1 => n42016, B2 => 
                           n47542, ZN => n36501);
   U795 : OAI22_X1 port map( A1 => n40611, A2 => n47537, B1 => n42015, B2 => 
                           n47543, ZN => n36502);
   U796 : OAI22_X1 port map( A1 => n40607, A2 => n47537, B1 => n42014, B2 => 
                           n47550, ZN => n36504);
   U797 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42753, ZN => n47573);
   U798 : OAI22_X1 port map( A1 => n40615, A2 => n47573, B1 => n42013, B2 => 
                           n47545, ZN => n36506);
   U799 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42750, ZN => n47572);
   U800 : OAI22_X1 port map( A1 => n40615, A2 => n47572, B1 => n42012, B2 => 
                           n47545, ZN => n36507);
   U801 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42748, ZN => n47574);
   U802 : OAI22_X1 port map( A1 => n40622, A2 => n47574, B1 => n42011, B2 => 
                           n47546, ZN => n36509);
   U803 : OAI22_X1 port map( A1 => n40622, A2 => n47573, B1 => n42010, B2 => 
                           n47546, ZN => n36510);
   U804 : OAI22_X1 port map( A1 => n40609, A2 => n47572, B1 => n42009, B2 => 
                           n47544, ZN => n36512);
   U805 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42751, ZN => n47571);
   U806 : OAI22_X1 port map( A1 => n40615, A2 => n47571, B1 => n42008, B2 => 
                           n47545, ZN => n36513);
   U807 : OAI22_X1 port map( A1 => n40620, A2 => n47513, B1 => n42007, B2 => 
                           n47558, ZN => n36516);
   U808 : OAI22_X1 port map( A1 => n40622, A2 => n47571, B1 => n42006, B2 => 
                           n47546, ZN => n36517);
   U809 : OAI22_X1 port map( A1 => n40609, A2 => n47571, B1 => n42005, B2 => 
                           n47544, ZN => n36518);
   U810 : OAI22_X1 port map( A1 => n40632, A2 => n47571, B1 => n42004, B2 => 
                           n47547, ZN => n36520);
   U811 : OAI22_X1 port map( A1 => n40609, A2 => n47526, B1 => n42003, B2 => 
                           n47544, ZN => n36521);
   U812 : OAI22_X1 port map( A1 => n40608, A2 => n47531, B1 => n42002, B2 => 
                           n47548, ZN => n36523);
   U813 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42754, ZN => n47575);
   U814 : OAI22_X1 port map( A1 => n40632, A2 => n47575, B1 => n42001, B2 => 
                           n47547, ZN => n36524);
   U815 : OAI22_X1 port map( A1 => n40626, A2 => n47525, B1 => n42000, B2 => 
                           n47553, ZN => n36526);
   U816 : OAI22_X1 port map( A1 => n40632, A2 => n47574, B1 => n41999, B2 => 
                           n47547, ZN => n36527);
   U817 : OAI22_X1 port map( A1 => n40615, A2 => n47574, B1 => n41998, B2 => 
                           n47545, ZN => n36528);
   U818 : OAI22_X1 port map( A1 => n40609, A2 => n47574, B1 => n41997, B2 => 
                           n47544, ZN => n36529);
   U819 : OAI22_X1 port map( A1 => n40632, A2 => n47572, B1 => n41996, B2 => 
                           n47547, ZN => n36530);
   U820 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42747, ZN => n47568);
   U821 : OAI22_X1 port map( A1 => n40608, A2 => n47568, B1 => n41995, B2 => 
                           n47548, ZN => n36531);
   U822 : OAI22_X1 port map( A1 => n40622, A2 => n47572, B1 => n41994, B2 => 
                           n47546, ZN => n36532);
   U823 : OAI22_X1 port map( A1 => n40608, A2 => n47570, B1 => n41993, B2 => 
                           n47548, ZN => n36533);
   U824 : OAI22_X1 port map( A1 => n40608, A2 => n47549, B1 => n41992, B2 => 
                           n47548, ZN => n36534);
   U825 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n42752, ZN => n47569);
   U826 : OAI22_X1 port map( A1 => n40607, A2 => n47569, B1 => n41991, B2 => 
                           n47550, ZN => n36536);
   U827 : OAI22_X1 port map( A1 => n40608, A2 => n47569, B1 => n41990, B2 => 
                           n47548, ZN => n36537);
   U828 : OAI22_X1 port map( A1 => n40627, A2 => n47525, B1 => n41989, B2 => 
                           n47554, ZN => n36539);
   U829 : OAI22_X1 port map( A1 => n40607, A2 => n47570, B1 => n41988, B2 => 
                           n47550, ZN => n36540);
   U830 : OAI22_X1 port map( A1 => n40607, A2 => n47568, B1 => n41987, B2 => 
                           n47550, ZN => n36541);
   U831 : OAI22_X1 port map( A1 => n40607, A2 => n47572, B1 => n41986, B2 => 
                           n47550, ZN => n36542);
   U832 : OAI22_X1 port map( A1 => n40606, A2 => n47574, B1 => n41985, B2 => 
                           n47551, ZN => n36544);
   U833 : OAI22_X1 port map( A1 => n40606, A2 => n47571, B1 => n41984, B2 => 
                           n47551, ZN => n36545);
   U834 : OAI22_X1 port map( A1 => n40606, A2 => n47573, B1 => n41983, B2 => 
                           n47551, ZN => n36546);
   U835 : OAI22_X1 port map( A1 => n40609, A2 => n47570, B1 => n41982, B2 => 
                           n47544, ZN => n36547);
   U836 : OAI22_X1 port map( A1 => n40609, A2 => n47569, B1 => n41981, B2 => 
                           n47544, ZN => n36548);
   U837 : OAI22_X1 port map( A1 => n40627, A2 => n47571, B1 => n41980, B2 => 
                           n47554, ZN => n36549);
   U838 : OAI22_X1 port map( A1 => n40625, A2 => n47574, B1 => n41979, B2 => 
                           n47552, ZN => n36551);
   U839 : OAI22_X1 port map( A1 => n40606, A2 => n47575, B1 => n41978, B2 => 
                           n47551, ZN => n36552);
   U840 : OAI22_X1 port map( A1 => n40608, A2 => n47573, B1 => n41977, B2 => 
                           n47548, ZN => n36553);
   U841 : OAI22_X1 port map( A1 => n40608, A2 => n47571, B1 => n41976, B2 => 
                           n47548, ZN => n36554);
   U842 : OAI22_X1 port map( A1 => n40608, A2 => n47572, B1 => n41975, B2 => 
                           n47548, ZN => n36555);
   U843 : OAI22_X1 port map( A1 => n40625, A2 => n47572, B1 => n41974, B2 => 
                           n47552, ZN => n36556);
   U844 : OAI22_X1 port map( A1 => n40625, A2 => n47571, B1 => n41973, B2 => 
                           n47552, ZN => n36557);
   U845 : OAI22_X1 port map( A1 => n40625, A2 => n47573, B1 => n41972, B2 => 
                           n47552, ZN => n36558);
   U846 : OAI22_X1 port map( A1 => n40609, A2 => n47534, B1 => n41971, B2 => 
                           n47544, ZN => n36559);
   U847 : OAI22_X1 port map( A1 => n40608, A2 => n47574, B1 => n41970, B2 => 
                           n47548, ZN => n36560);
   U848 : OAI22_X1 port map( A1 => n40626, A2 => n47574, B1 => n41969, B2 => 
                           n47553, ZN => n36561);
   U849 : OAI22_X1 port map( A1 => n40626, A2 => n47572, B1 => n41968, B2 => 
                           n47553, ZN => n36562);
   U850 : OAI22_X1 port map( A1 => n40626, A2 => n47571, B1 => n41967, B2 => 
                           n47553, ZN => n36563);
   U851 : OAI22_X1 port map( A1 => n40626, A2 => n47573, B1 => n41966, B2 => 
                           n47553, ZN => n36564);
   U852 : OAI22_X1 port map( A1 => n40632, A2 => n47531, B1 => n41965, B2 => 
                           n47547, ZN => n36565);
   U853 : OAI22_X1 port map( A1 => n40627, A2 => n47574, B1 => n41964, B2 => 
                           n47554, ZN => n36566);
   U854 : OAI22_X1 port map( A1 => n40627, A2 => n47572, B1 => n41963, B2 => 
                           n47554, ZN => n36567);
   U855 : OAI22_X1 port map( A1 => n40627, A2 => n47573, B1 => n41962, B2 => 
                           n47554, ZN => n36568);
   U856 : OAI22_X1 port map( A1 => n40607, A2 => n47571, B1 => n41961, B2 => 
                           n47550, ZN => n36569);
   U857 : OAI22_X1 port map( A1 => n40608, A2 => n47575, B1 => n41960, B2 => 
                           n47548, ZN => n36570);
   U858 : OAI22_X1 port map( A1 => n40622, A2 => n47555, B1 => n41959, B2 => 
                           n47546, ZN => n36571);
   U859 : OAI22_X1 port map( A1 => n40618, A2 => n47568, B1 => n41958, B2 => 
                           n47557, ZN => n36573);
   U860 : OAI22_X1 port map( A1 => n40607, A2 => n47573, B1 => n41957, B2 => 
                           n47550, ZN => n36574);
   U861 : OAI22_X1 port map( A1 => n40607, A2 => n47534, B1 => n41956, B2 => 
                           n47550, ZN => n36575);
   U862 : OAI22_X1 port map( A1 => n40620, A2 => n47568, B1 => n41955, B2 => 
                           n47558, ZN => n36576);
   U863 : OAI22_X1 port map( A1 => n40626, A2 => n47526, B1 => n41954, B2 => 
                           n47553, ZN => n36577);
   U864 : OAI22_X1 port map( A1 => n40622, A2 => n47568, B1 => n41953, B2 => 
                           n47546, ZN => n36578);
   U865 : OAI22_X1 port map( A1 => n40618, A2 => n47522, B1 => n41952, B2 => 
                           n47557, ZN => n36580);
   U866 : OAI22_X1 port map( A1 => n40607, A2 => n47574, B1 => n41951, B2 => 
                           n47550, ZN => n36581);
   U867 : OAI22_X1 port map( A1 => n40625, A2 => n47575, B1 => n41950, B2 => 
                           n47552, ZN => n36582);
   U868 : OAI22_X1 port map( A1 => n40626, A2 => n47555, B1 => n41949, B2 => 
                           n47553, ZN => n36583);
   U869 : OAI22_X1 port map( A1 => n40606, A2 => n47525, B1 => n41948, B2 => 
                           n47551, ZN => n36585);
   U870 : OAI22_X1 port map( A1 => n40624, A2 => n47573, B1 => n41947, B2 => 
                           n47556, ZN => n36587);
   U871 : OAI22_X1 port map( A1 => n40624, A2 => n47572, B1 => n41946, B2 => 
                           n47556, ZN => n36588);
   U872 : OAI22_X1 port map( A1 => n40626, A2 => n47570, B1 => n41945, B2 => 
                           n47553, ZN => n36589);
   U873 : OAI22_X1 port map( A1 => n40624, A2 => n47564, B1 => n41944, B2 => 
                           n47556, ZN => n36590);
   U874 : OAI22_X1 port map( A1 => n40625, A2 => n47570, B1 => n41943, B2 => 
                           n47552, ZN => n36591);
   U875 : OAI22_X1 port map( A1 => n40625, A2 => n47568, B1 => n41942, B2 => 
                           n47552, ZN => n36592);
   U876 : OAI22_X1 port map( A1 => n40627, A2 => n47555, B1 => n41941, B2 => 
                           n47554, ZN => n36593);
   U877 : OAI22_X1 port map( A1 => n40625, A2 => n47526, B1 => n41940, B2 => 
                           n47552, ZN => n36594);
   U878 : OAI22_X1 port map( A1 => n40624, A2 => n47569, B1 => n41939, B2 => 
                           n47556, ZN => n36595);
   U879 : OAI22_X1 port map( A1 => n40624, A2 => n47574, B1 => n41938, B2 => 
                           n47556, ZN => n36596);
   U880 : OAI22_X1 port map( A1 => n40607, A2 => n47575, B1 => n41937, B2 => 
                           n47550, ZN => n36597);
   U881 : OAI22_X1 port map( A1 => n40627, A2 => n47568, B1 => n41936, B2 => 
                           n47554, ZN => n36598);
   U882 : OAI22_X1 port map( A1 => n40624, A2 => n47526, B1 => n41935, B2 => 
                           n47556, ZN => n36599);
   U883 : OAI22_X1 port map( A1 => n40624, A2 => n47555, B1 => n41934, B2 => 
                           n47556, ZN => n36600);
   U884 : OAI22_X1 port map( A1 => n40624, A2 => n47568, B1 => n41933, B2 => 
                           n47556, ZN => n36601);
   U885 : OAI22_X1 port map( A1 => n40625, A2 => n47522, B1 => n41932, B2 => 
                           n47552, ZN => n36602);
   U886 : OAI22_X1 port map( A1 => n40624, A2 => n47570, B1 => n41931, B2 => 
                           n47556, ZN => n36603);
   U887 : OAI22_X1 port map( A1 => n40624, A2 => n47571, B1 => n41930, B2 => 
                           n47556, ZN => n36604);
   U888 : OAI22_X1 port map( A1 => n40626, A2 => n47575, B1 => n41929, B2 => 
                           n47553, ZN => n36605);
   U889 : OAI22_X1 port map( A1 => n40612, A2 => n47568, B1 => n41928, B2 => 
                           n47559, ZN => n36607);
   U890 : OAI22_X1 port map( A1 => n40626, A2 => n47569, B1 => n41927, B2 => 
                           n47553, ZN => n36608);
   U891 : OAI22_X1 port map( A1 => n40616, A2 => n47568, B1 => n41926, B2 => 
                           n47560, ZN => n36610);
   U892 : OAI22_X1 port map( A1 => n40625, A2 => n47533, B1 => n41925, B2 => 
                           n47552, ZN => n36611);
   U893 : OAI22_X1 port map( A1 => n40627, A2 => n47570, B1 => n41924, B2 => 
                           n47554, ZN => n36612);
   U894 : OAI22_X1 port map( A1 => n40618, A2 => n47523, B1 => n41923, B2 => 
                           n47557, ZN => n36613);
   U895 : OAI22_X1 port map( A1 => n40632, A2 => n47570, B1 => n41922, B2 => 
                           n47547, ZN => n36614);
   U896 : OAI22_X1 port map( A1 => n40625, A2 => n47569, B1 => n41921, B2 => 
                           n47552, ZN => n36615);
   U897 : OAI22_X1 port map( A1 => n40627, A2 => n47569, B1 => n41920, B2 => 
                           n47554, ZN => n36616);
   U898 : OAI22_X1 port map( A1 => n40627, A2 => n47530, B1 => n41919, B2 => 
                           n47554, ZN => n36617);
   U899 : OAI22_X1 port map( A1 => n40620, A2 => n47523, B1 => n41918, B2 => 
                           n47558, ZN => n36619);
   U900 : OAI22_X1 port map( A1 => n40626, A2 => n47568, B1 => n41917, B2 => 
                           n47553, ZN => n36620);
   U901 : OAI22_X1 port map( A1 => n40627, A2 => n47575, B1 => n41916, B2 => 
                           n47554, ZN => n36621);
   U902 : OAI22_X1 port map( A1 => n40607, A2 => n47555, B1 => n41915, B2 => 
                           n47550, ZN => n36622);
   U903 : OAI22_X1 port map( A1 => n40608, A2 => n47555, B1 => n41914, B2 => 
                           n47548, ZN => n36623);
   U904 : OAI22_X1 port map( A1 => n40609, A2 => n47575, B1 => n41913, B2 => 
                           n47544, ZN => n36624);
   U905 : OAI22_X1 port map( A1 => n40609, A2 => n47555, B1 => n41912, B2 => 
                           n47544, ZN => n36625);
   U906 : OAI22_X1 port map( A1 => n40618, A2 => n47555, B1 => n41911, B2 => 
                           n47557, ZN => n36626);
   U907 : OAI22_X1 port map( A1 => n40632, A2 => n47569, B1 => n41910, B2 => 
                           n47547, ZN => n36627);
   U908 : OAI22_X1 port map( A1 => n40620, A2 => n47574, B1 => n41909, B2 => 
                           n47558, ZN => n36628);
   U909 : OAI22_X1 port map( A1 => n40615, A2 => n47526, B1 => n41908, B2 => 
                           n47545, ZN => n36629);
   U910 : OAI22_X1 port map( A1 => n40616, A2 => n47574, B1 => n41907, B2 => 
                           n47560, ZN => n36630);
   U911 : OAI22_X1 port map( A1 => n40618, A2 => n47574, B1 => n41906, B2 => 
                           n47557, ZN => n36631);
   U912 : OAI22_X1 port map( A1 => n40622, A2 => n47570, B1 => n41905, B2 => 
                           n47546, ZN => n36632);
   U913 : OAI22_X1 port map( A1 => n40612, A2 => n47571, B1 => n41904, B2 => 
                           n47559, ZN => n36633);
   U914 : OAI22_X1 port map( A1 => n40622, A2 => n47575, B1 => n41903, B2 => 
                           n47546, ZN => n36634);
   U915 : OAI22_X1 port map( A1 => n40612, A2 => n47574, B1 => n41902, B2 => 
                           n47559, ZN => n36635);
   U916 : OAI22_X1 port map( A1 => n40606, A2 => n47569, B1 => n41901, B2 => 
                           n47551, ZN => n36636);
   U917 : OAI22_X1 port map( A1 => n40618, A2 => n47570, B1 => n41900, B2 => 
                           n47557, ZN => n36637);
   U918 : OAI22_X1 port map( A1 => n40624, A2 => n47575, B1 => n41899, B2 => 
                           n47556, ZN => n36639);
   U919 : OAI22_X1 port map( A1 => n40620, A2 => n47575, B1 => n41898, B2 => 
                           n47558, ZN => n36640);
   U920 : OAI22_X1 port map( A1 => n40620, A2 => n47573, B1 => n41897, B2 => 
                           n47558, ZN => n36641);
   U921 : OAI22_X1 port map( A1 => n40620, A2 => n47569, B1 => n41896, B2 => 
                           n47558, ZN => n36642);
   U922 : OAI22_X1 port map( A1 => n40612, A2 => n47555, B1 => n41895, B2 => 
                           n47559, ZN => n36644);
   U923 : OAI22_X1 port map( A1 => n40620, A2 => n47571, B1 => n41894, B2 => 
                           n47558, ZN => n36645);
   U924 : OAI22_X1 port map( A1 => n40615, A2 => n47564, B1 => n41893, B2 => 
                           n47545, ZN => n36646);
   U925 : OAI22_X1 port map( A1 => n40620, A2 => n47572, B1 => n41892, B2 => 
                           n47558, ZN => n36647);
   U926 : OAI22_X1 port map( A1 => n40609, A2 => n47568, B1 => n41891, B2 => 
                           n47544, ZN => n36648);
   U927 : OAI22_X1 port map( A1 => n40618, A2 => n47575, B1 => n41890, B2 => 
                           n47557, ZN => n36649);
   U928 : OAI22_X1 port map( A1 => n40616, A2 => n47575, B1 => n41889, B2 => 
                           n47560, ZN => n36650);
   U929 : OAI22_X1 port map( A1 => n40615, A2 => n47575, B1 => n41888, B2 => 
                           n47545, ZN => n36651);
   U930 : OAI22_X1 port map( A1 => n40632, A2 => n47568, B1 => n41887, B2 => 
                           n47547, ZN => n36652);
   U931 : OAI22_X1 port map( A1 => n40616, A2 => n47564, B1 => n41886, B2 => 
                           n47560, ZN => n36653);
   U932 : OAI22_X1 port map( A1 => n40632, A2 => n47533, B1 => n41885, B2 => 
                           n47547, ZN => n36654);
   U933 : OAI22_X1 port map( A1 => n40616, A2 => n47570, B1 => n41884, B2 => 
                           n47560, ZN => n36655);
   U934 : OAI22_X1 port map( A1 => n40616, A2 => n47571, B1 => n41883, B2 => 
                           n47560, ZN => n36656);
   U935 : OAI22_X1 port map( A1 => n40618, A2 => n47571, B1 => n41882, B2 => 
                           n47557, ZN => n36657);
   U936 : OAI22_X1 port map( A1 => n40612, A2 => n47575, B1 => n41881, B2 => 
                           n47559, ZN => n36658);
   U937 : OAI22_X1 port map( A1 => n40615, A2 => n47570, B1 => n41880, B2 => 
                           n47545, ZN => n36659);
   U938 : OAI22_X1 port map( A1 => n40620, A2 => n47570, B1 => n41879, B2 => 
                           n47558, ZN => n36660);
   U939 : OAI22_X1 port map( A1 => n40606, A2 => n47533, B1 => n41878, B2 => 
                           n47551, ZN => n36661);
   U940 : OAI22_X1 port map( A1 => n40616, A2 => n47530, B1 => n41877, B2 => 
                           n47560, ZN => n36663);
   U941 : OAI22_X1 port map( A1 => n40606, A2 => n47568, B1 => n41876, B2 => 
                           n47551, ZN => n36664);
   U942 : OAI22_X1 port map( A1 => n40612, A2 => n47570, B1 => n41875, B2 => 
                           n47559, ZN => n36665);
   U943 : OAI22_X1 port map( A1 => n40607, A2 => n47529, B1 => n41874, B2 => 
                           n47550, ZN => n36666);
   U944 : OAI22_X1 port map( A1 => n40632, A2 => n47573, B1 => n41873, B2 => 
                           n47547, ZN => n36667);
   U945 : OAI22_X1 port map( A1 => n40616, A2 => n47533, B1 => n41872, B2 => 
                           n47560, ZN => n36668);
   U946 : OAI22_X1 port map( A1 => n40609, A2 => n47573, B1 => n41871, B2 => 
                           n47544, ZN => n36669);
   U947 : OAI22_X1 port map( A1 => n40612, A2 => n47564, B1 => n41870, B2 => 
                           n47559, ZN => n36670);
   U948 : OAI22_X1 port map( A1 => n40616, A2 => n47572, B1 => n41869, B2 => 
                           n47560, ZN => n36671);
   U949 : OAI22_X1 port map( A1 => n40618, A2 => n47573, B1 => n41868, B2 => 
                           n47557, ZN => n36672);
   U950 : OAI22_X1 port map( A1 => n40622, A2 => n47569, B1 => n41867, B2 => 
                           n47546, ZN => n36673);
   U951 : OAI22_X1 port map( A1 => n40615, A2 => n47533, B1 => n41866, B2 => 
                           n47545, ZN => n36675);
   U952 : OAI22_X1 port map( A1 => n40620, A2 => n47529, B1 => n41865, B2 => 
                           n47558, ZN => n36678);
   U953 : OAI22_X1 port map( A1 => n40606, A2 => n47570, B1 => n41864, B2 => 
                           n47551, ZN => n36679);
   U954 : OAI22_X1 port map( A1 => n40615, A2 => n47568, B1 => n41863, B2 => 
                           n47545, ZN => n36680);
   U955 : OAI22_X1 port map( A1 => n40606, A2 => n47572, B1 => n41862, B2 => 
                           n47551, ZN => n36681);
   U956 : OAI22_X1 port map( A1 => n40618, A2 => n47572, B1 => n41861, B2 => 
                           n47557, ZN => n36682);
   U957 : OAI22_X1 port map( A1 => n40606, A2 => n47522, B1 => n41860, B2 => 
                           n47551, ZN => n36684);
   U958 : OAI22_X1 port map( A1 => n40632, A2 => n47526, B1 => n41859, B2 => 
                           n47547, ZN => n36685);
   U959 : OAI22_X1 port map( A1 => n40612, A2 => n47572, B1 => n41858, B2 => 
                           n47559, ZN => n36686);
   U960 : OAI22_X1 port map( A1 => n40618, A2 => n47569, B1 => n41857, B2 => 
                           n47557, ZN => n36688);
   U961 : OAI22_X1 port map( A1 => n40616, A2 => n47569, B1 => n41856, B2 => 
                           n47560, ZN => n36689);
   U962 : OAI22_X1 port map( A1 => n40612, A2 => n47573, B1 => n41855, B2 => 
                           n47559, ZN => n36690);
   U963 : OAI22_X1 port map( A1 => n40612, A2 => n47534, B1 => n41854, B2 => 
                           n47559, ZN => n36691);
   U964 : OAI22_X1 port map( A1 => n40622, A2 => n47530, B1 => n41853, B2 => 
                           n47546, ZN => n36693);
   U965 : OAI22_X1 port map( A1 => n40616, A2 => n47573, B1 => n41852, B2 => 
                           n47560, ZN => n36695);
   U966 : OAI22_X1 port map( A1 => n40612, A2 => n47569, B1 => n41851, B2 => 
                           n47559, ZN => n36697);
   U967 : OAI22_X1 port map( A1 => n40615, A2 => n47569, B1 => n41850, B2 => 
                           n47545, ZN => n36699);
   U968 : OAI22_X1 port map( A1 => n40622, A2 => n47564, B1 => n41849, B2 => 
                           n47546, ZN => n36702);
   U969 : OAI22_X1 port map( A1 => n40646, A2 => n47568, B1 => n41848, B2 => 
                           n47562, ZN => n36704);
   U970 : OAI22_X1 port map( A1 => n40642, A2 => n47564, B1 => n41847, B2 => 
                           n47561, ZN => n36706);
   U971 : OAI22_X1 port map( A1 => n40646, A2 => n47531, B1 => n41846, B2 => 
                           n47562, ZN => n36707);
   U972 : OAI22_X1 port map( A1 => n40638, A2 => n47564, B1 => n41845, B2 => 
                           n47563, ZN => n36709);
   U973 : OAI22_X1 port map( A1 => n40604, A2 => n47575, B1 => n41844, B2 => 
                           n47566, ZN => n36711);
   U974 : OAI22_X1 port map( A1 => n40638, A2 => n47520, B1 => n41843, B2 => 
                           n47563, ZN => n36713);
   U975 : OAI22_X1 port map( A1 => n40647, A2 => n47526, B1 => n41842, B2 => 
                           n47567, ZN => n36716);
   U976 : OAI22_X1 port map( A1 => n40637, A2 => n47564, B1 => n41841, B2 => 
                           n47511, ZN => n36719);
   U977 : OAI22_X1 port map( A1 => n40638, A2 => n47568, B1 => n41840, B2 => 
                           n47563, ZN => n36720);
   U978 : OAI22_X1 port map( A1 => n40638, A2 => n47571, B1 => n41839, B2 => 
                           n47563, ZN => n36721);
   U979 : OAI22_X1 port map( A1 => n40642, A2 => n47571, B1 => n41838, B2 => 
                           n47561, ZN => n36722);
   U980 : OAI22_X1 port map( A1 => n40642, A2 => n47568, B1 => n41837, B2 => 
                           n47561, ZN => n36723);
   U981 : OAI22_X1 port map( A1 => n40637, A2 => n47571, B1 => n41836, B2 => 
                           n47511, ZN => n36724);
   U982 : OAI22_X1 port map( A1 => n40642, A2 => n47574, B1 => n41835, B2 => 
                           n47561, ZN => n36725);
   U983 : OAI22_X1 port map( A1 => n40628, A2 => n47568, B1 => n41834, B2 => 
                           n47512, ZN => n36727);
   U984 : OAI22_X1 port map( A1 => n40637, A2 => n47521, B1 => n41833, B2 => 
                           n47511, ZN => n36728);
   U985 : OAI22_X1 port map( A1 => n40637, A2 => n47568, B1 => n41832, B2 => 
                           n47511, ZN => n36729);
   U986 : OAI22_X1 port map( A1 => n40628, A2 => n47534, B1 => n41831, B2 => 
                           n47512, ZN => n36731);
   U987 : OAI22_X1 port map( A1 => n40628, A2 => n47569, B1 => n41830, B2 => 
                           n47512, ZN => n36732);
   U988 : OAI22_X1 port map( A1 => n40628, A2 => n47573, B1 => n41829, B2 => 
                           n47512, ZN => n36733);
   U989 : OAI22_X1 port map( A1 => n40642, A2 => n47521, B1 => n41828, B2 => 
                           n47561, ZN => n36734);
   U990 : OAI22_X1 port map( A1 => n40628, A2 => n47572, B1 => n41827, B2 => 
                           n47512, ZN => n36735);
   U991 : OAI22_X1 port map( A1 => n40605, A2 => n47575, B1 => n41826, B2 => 
                           n47565, ZN => n36737);
   U992 : OAI22_X1 port map( A1 => n40637, A2 => n47569, B1 => n41825, B2 => 
                           n47511, ZN => n36738);
   U993 : OAI22_X1 port map( A1 => n40605, A2 => n47570, B1 => n41824, B2 => 
                           n47565, ZN => n36739);
   U994 : OAI22_X1 port map( A1 => n40638, A2 => n47569, B1 => n41823, B2 => 
                           n47563, ZN => n36740);
   U995 : OAI22_X1 port map( A1 => n40642, A2 => n47569, B1 => n41822, B2 => 
                           n47561, ZN => n36741);
   U996 : OAI22_X1 port map( A1 => n40628, A2 => n47570, B1 => n41821, B2 => 
                           n47512, ZN => n36742);
   U997 : OAI22_X1 port map( A1 => n40638, A2 => n47574, B1 => n41820, B2 => 
                           n47563, ZN => n36743);
   U998 : OAI22_X1 port map( A1 => n40604, A2 => n47569, B1 => n41819, B2 => 
                           n47566, ZN => n36744);
   U999 : CLKBUF_X1 port map( A => n47570, Z => n47576);
   U1000 : OAI22_X1 port map( A1 => n40604, A2 => n47576, B1 => n41818, B2 => 
                           n47566, ZN => n36745);
   U1001 : OAI22_X1 port map( A1 => n40604, A2 => n47568, B1 => n41817, B2 => 
                           n47566, ZN => n36746);
   U1002 : OAI22_X1 port map( A1 => n40628, A2 => n47528, B1 => n41816, B2 => 
                           n47512, ZN => n36747);
   U1003 : OAI22_X1 port map( A1 => n40604, A2 => n47528, B1 => n41815, B2 => 
                           n47566, ZN => n36749);
   U1004 : OAI22_X1 port map( A1 => n40647, A2 => n47534, B1 => n41814, B2 => 
                           n47567, ZN => n36750);
   U1005 : OAI22_X1 port map( A1 => n40646, A2 => n47534, B1 => n41813, B2 => 
                           n47562, ZN => n36752);
   U1006 : OAI22_X1 port map( A1 => n40637, A2 => n47572, B1 => n41812, B2 => 
                           n47511, ZN => n36753);
   U1007 : OAI22_X1 port map( A1 => n40647, A2 => n47575, B1 => n41811, B2 => 
                           n47567, ZN => n36754);
   U1008 : OAI22_X1 port map( A1 => n40637, A2 => n47574, B1 => n41810, B2 => 
                           n47511, ZN => n36755);
   U1009 : OAI22_X1 port map( A1 => n40604, A2 => n47531, B1 => n41809, B2 => 
                           n47566, ZN => n36756);
   U1010 : OAI22_X1 port map( A1 => n40646, A2 => n47576, B1 => n41808, B2 => 
                           n47562, ZN => n36757);
   U1011 : OAI22_X1 port map( A1 => n40642, A2 => n47572, B1 => n41807, B2 => 
                           n47561, ZN => n36758);
   U1012 : OAI22_X1 port map( A1 => n40647, A2 => n47568, B1 => n41806, B2 => 
                           n47567, ZN => n36759);
   U1013 : OAI22_X1 port map( A1 => n40605, A2 => n47569, B1 => n41805, B2 => 
                           n47565, ZN => n36760);
   U1014 : OAI22_X1 port map( A1 => n40628, A2 => n47574, B1 => n41804, B2 => 
                           n47512, ZN => n36761);
   U1015 : OAI22_X1 port map( A1 => n40638, A2 => n47575, B1 => n41803, B2 => 
                           n47563, ZN => n36762);
   U1016 : OAI22_X1 port map( A1 => n40638, A2 => n47572, B1 => n41802, B2 => 
                           n47563, ZN => n36763);
   U1017 : OAI22_X1 port map( A1 => n40604, A2 => n47574, B1 => n41801, B2 => 
                           n47566, ZN => n36764);
   U1018 : OAI22_X1 port map( A1 => n40642, A2 => n47570, B1 => n41800, B2 => 
                           n47561, ZN => n36765);
   U1019 : OAI22_X1 port map( A1 => n40638, A2 => n47570, B1 => n41799, B2 => 
                           n47563, ZN => n36766);
   U1020 : OAI22_X1 port map( A1 => n40646, A2 => n47575, B1 => n41798, B2 => 
                           n47562, ZN => n36767);
   U1021 : OAI22_X1 port map( A1 => n40642, A2 => n47575, B1 => n41797, B2 => 
                           n47561, ZN => n36768);
   U1022 : OAI22_X1 port map( A1 => n40642, A2 => n47573, B1 => n41796, B2 => 
                           n47561, ZN => n36769);
   U1023 : OAI22_X1 port map( A1 => n40605, A2 => n47573, B1 => n41795, B2 => 
                           n47565, ZN => n36770);
   U1024 : OAI22_X1 port map( A1 => n40646, A2 => n47573, B1 => n41794, B2 => 
                           n47562, ZN => n36771);
   U1025 : OAI22_X1 port map( A1 => n40647, A2 => n47569, B1 => n41793, B2 => 
                           n47567, ZN => n36772);
   U1026 : OAI22_X1 port map( A1 => n40646, A2 => n47569, B1 => n41792, B2 => 
                           n47562, ZN => n36773);
   U1027 : OAI22_X1 port map( A1 => n40647, A2 => n47570, B1 => n41791, B2 => 
                           n47567, ZN => n36774);
   U1028 : OAI22_X1 port map( A1 => n40637, A2 => n47570, B1 => n41790, B2 => 
                           n47511, ZN => n36775);
   U1029 : OAI22_X1 port map( A1 => n40647, A2 => n47574, B1 => n41789, B2 => 
                           n47567, ZN => n36776);
   U1030 : OAI22_X1 port map( A1 => n40628, A2 => n47575, B1 => n41788, B2 => 
                           n47512, ZN => n36777);
   U1031 : OAI22_X1 port map( A1 => n40604, A2 => n47571, B1 => n41787, B2 => 
                           n47566, ZN => n36778);
   U1032 : OAI22_X1 port map( A1 => n40605, A2 => n47572, B1 => n41786, B2 => 
                           n47565, ZN => n36779);
   U1033 : OAI22_X1 port map( A1 => n40637, A2 => n47575, B1 => n41785, B2 => 
                           n47511, ZN => n36780);
   U1034 : OAI22_X1 port map( A1 => n40647, A2 => n47572, B1 => n41784, B2 => 
                           n47567, ZN => n36781);
   U1035 : OAI22_X1 port map( A1 => n40646, A2 => n47571, B1 => n41783, B2 => 
                           n47562, ZN => n36782);
   U1036 : OAI22_X1 port map( A1 => n40605, A2 => n47531, B1 => n41782, B2 => 
                           n47565, ZN => n36784);
   U1037 : OAI22_X1 port map( A1 => n40605, A2 => n47571, B1 => n41781, B2 => 
                           n47565, ZN => n36785);
   U1038 : OAI22_X1 port map( A1 => n40628, A2 => n47571, B1 => n41780, B2 => 
                           n47512, ZN => n36786);
   U1039 : OAI22_X1 port map( A1 => n40604, A2 => n47573, B1 => n41779, B2 => 
                           n47566, ZN => n36787);
   U1040 : OAI22_X1 port map( A1 => n40605, A2 => n47521, B1 => n41778, B2 => 
                           n47565, ZN => n36789);
   U1041 : OAI22_X1 port map( A1 => n40638, A2 => n47573, B1 => n41777, B2 => 
                           n47563, ZN => n36790);
   U1042 : OAI22_X1 port map( A1 => n40605, A2 => n47568, B1 => n41776, B2 => 
                           n47565, ZN => n36791);
   U1043 : OAI22_X1 port map( A1 => n40647, A2 => n47571, B1 => n41775, B2 => 
                           n47567, ZN => n36792);
   U1044 : OAI22_X1 port map( A1 => n40637, A2 => n47573, B1 => n41774, B2 => 
                           n47511, ZN => n36793);
   U1045 : OAI22_X1 port map( A1 => n40646, A2 => n47574, B1 => n41773, B2 => 
                           n47562, ZN => n36794);
   U1046 : OAI22_X1 port map( A1 => n40646, A2 => n47572, B1 => n41772, B2 => 
                           n47562, ZN => n36795);
   U1047 : OAI22_X1 port map( A1 => n40604, A2 => n47572, B1 => n41771, B2 => 
                           n47566, ZN => n36796);
   U1048 : OAI22_X1 port map( A1 => n40605, A2 => n47574, B1 => n41770, B2 => 
                           n47565, ZN => n36797);
   U1049 : OAI22_X1 port map( A1 => n40647, A2 => n47573, B1 => n41769, B2 => 
                           n47567, ZN => n36798);
   U1050 : OAI22_X1 port map( A1 => n40636, A2 => n47568, B1 => n41768, B2 => 
                           n47542, ZN => n36800);
   U1051 : OAI22_X1 port map( A1 => n40611, A2 => n47569, B1 => n41767, B2 => 
                           n47543, ZN => n36802);
   U1052 : OAI22_X1 port map( A1 => n40610, A2 => n47569, B1 => n41766, B2 => 
                           n47540, ZN => n36804);
   U1053 : OAI22_X1 port map( A1 => n40619, A2 => n47569, B1 => n41765, B2 => 
                           n47541, ZN => n36806);
   U1054 : OAI22_X1 port map( A1 => n40614, A2 => n47569, B1 => n41764, B2 => 
                           n47536, ZN => n36808);
   U1055 : OAI22_X1 port map( A1 => n40610, A2 => n47570, B1 => n41763, B2 => 
                           n47540, ZN => n36809);
   U1056 : OAI22_X1 port map( A1 => n40611, A2 => n47576, B1 => n41762, B2 => 
                           n47543, ZN => n36810);
   U1057 : OAI22_X1 port map( A1 => n40623, A2 => n47571, B1 => n41761, B2 => 
                           n47535, ZN => n36812);
   U1058 : OAI22_X1 port map( A1 => n40613, A2 => n47576, B1 => n41760, B2 => 
                           n47532, ZN => n36814);
   U1059 : OAI22_X1 port map( A1 => n40610, A2 => n47571, B1 => n41759, B2 => 
                           n47540, ZN => n36815);
   U1060 : OAI22_X1 port map( A1 => n40614, A2 => n47576, B1 => n41758, B2 => 
                           n47536, ZN => n36816);
   U1061 : OAI22_X1 port map( A1 => n40613, A2 => n47569, B1 => n41757, B2 => 
                           n47532, ZN => n36817);
   U1062 : OAI22_X1 port map( A1 => n40614, A2 => n47572, B1 => n41756, B2 => 
                           n47536, ZN => n36818);
   U1063 : OAI22_X1 port map( A1 => n40619, A2 => n47572, B1 => n41755, B2 => 
                           n47541, ZN => n36819);
   U1064 : OAI22_X1 port map( A1 => n40619, A2 => n47573, B1 => n41754, B2 => 
                           n47541, ZN => n36820);
   U1065 : OAI22_X1 port map( A1 => n40610, A2 => n47573, B1 => n41753, B2 => 
                           n47540, ZN => n36821);
   U1066 : OAI22_X1 port map( A1 => n40614, A2 => n47571, B1 => n41752, B2 => 
                           n47536, ZN => n36822);
   U1067 : OAI22_X1 port map( A1 => n40619, A2 => n47571, B1 => n41751, B2 => 
                           n47541, ZN => n36823);
   U1068 : OAI22_X1 port map( A1 => n40623, A2 => n47572, B1 => n41750, B2 => 
                           n47535, ZN => n36824);
   U1069 : OAI22_X1 port map( A1 => n40610, A2 => n47572, B1 => n41749, B2 => 
                           n47540, ZN => n36825);
   U1070 : OAI22_X1 port map( A1 => n40613, A2 => n47571, B1 => n41748, B2 => 
                           n47532, ZN => n36826);
   U1071 : OAI22_X1 port map( A1 => n40614, A2 => n47573, B1 => n41747, B2 => 
                           n47536, ZN => n36827);
   U1072 : OAI22_X1 port map( A1 => n40613, A2 => n47573, B1 => n41746, B2 => 
                           n47532, ZN => n36828);
   U1073 : OAI22_X1 port map( A1 => n40623, A2 => n47574, B1 => n41745, B2 => 
                           n47535, ZN => n36829);
   U1074 : OAI22_X1 port map( A1 => n40623, A2 => n47573, B1 => n41744, B2 => 
                           n47535, ZN => n36830);
   U1075 : OAI22_X1 port map( A1 => n40613, A2 => n47572, B1 => n41743, B2 => 
                           n47532, ZN => n36831);
   U1076 : OAI22_X1 port map( A1 => n40610, A2 => n47575, B1 => n41742, B2 => 
                           n47540, ZN => n36832);
   U1077 : OAI22_X1 port map( A1 => n40617, A2 => n47568, B1 => n41741, B2 => 
                           n47538, ZN => n36834);
   U1078 : OAI22_X1 port map( A1 => n40621, A2 => n47573, B1 => n41740, B2 => 
                           n47539, ZN => n36836);
   U1079 : OAI22_X1 port map( A1 => n40621, A2 => n47569, B1 => n41739, B2 => 
                           n47539, ZN => n36837);
   U1080 : OAI22_X1 port map( A1 => n40636, A2 => n47575, B1 => n41738, B2 => 
                           n47542, ZN => n36838);
   U1081 : OAI22_X1 port map( A1 => n40621, A2 => n47571, B1 => n41737, B2 => 
                           n47539, ZN => n36839);
   U1082 : OAI22_X1 port map( A1 => n40623, A2 => n47576, B1 => n41736, B2 => 
                           n47535, ZN => n36840);
   U1083 : OAI22_X1 port map( A1 => n40621, A2 => n47572, B1 => n41735, B2 => 
                           n47539, ZN => n36841);
   U1084 : OAI22_X1 port map( A1 => n40621, A2 => n47576, B1 => n41734, B2 => 
                           n47539, ZN => n36842);
   U1085 : OAI22_X1 port map( A1 => n40623, A2 => n47569, B1 => n41733, B2 => 
                           n47535, ZN => n36843);
   U1086 : OAI22_X1 port map( A1 => n40617, A2 => n47576, B1 => n41732, B2 => 
                           n47538, ZN => n36844);
   U1087 : OAI22_X1 port map( A1 => n40614, A2 => n47574, B1 => n41731, B2 => 
                           n47536, ZN => n36845);
   U1088 : OAI22_X1 port map( A1 => n40613, A2 => n47574, B1 => n41730, B2 => 
                           n47532, ZN => n36846);
   U1089 : OAI22_X1 port map( A1 => n40619, A2 => n47568, B1 => n41729, B2 => 
                           n47541, ZN => n36847);
   U1090 : OAI22_X1 port map( A1 => n40621, A2 => n47575, B1 => n41728, B2 => 
                           n47539, ZN => n36848);
   U1091 : OAI22_X1 port map( A1 => n40623, A2 => n47575, B1 => n41727, B2 => 
                           n47535, ZN => n36849);
   U1092 : OAI22_X1 port map( A1 => n40610, A2 => n47574, B1 => n41726, B2 => 
                           n47540, ZN => n36850);
   U1093 : OAI22_X1 port map( A1 => n40636, A2 => n47569, B1 => n41725, B2 => 
                           n47542, ZN => n36852);
   U1094 : OAI22_X1 port map( A1 => n40613, A2 => n47568, B1 => n41724, B2 => 
                           n47532, ZN => n36853);
   U1095 : OAI22_X1 port map( A1 => n40611, A2 => n47575, B1 => n41723, B2 => 
                           n47543, ZN => n36854);
   U1096 : OAI22_X1 port map( A1 => n40613, A2 => n47575, B1 => n41722, B2 => 
                           n47532, ZN => n36856);
   U1097 : OAI22_X1 port map( A1 => n40619, A2 => n47576, B1 => n41721, B2 => 
                           n47541, ZN => n36858);
   U1098 : OAI22_X1 port map( A1 => n40614, A2 => n47575, B1 => n41720, B2 => 
                           n47536, ZN => n36859);
   U1099 : OAI22_X1 port map( A1 => n40621, A2 => n47574, B1 => n41719, B2 => 
                           n47539, ZN => n36860);
   U1100 : OAI22_X1 port map( A1 => n40611, A2 => n47572, B1 => n41718, B2 => 
                           n47543, ZN => n36861);
   U1101 : OAI22_X1 port map( A1 => n40621, A2 => n47568, B1 => n41717, B2 => 
                           n47539, ZN => n36862);
   U1102 : OAI22_X1 port map( A1 => n40636, A2 => n47576, B1 => n41716, B2 => 
                           n47542, ZN => n36864);
   U1103 : OAI22_X1 port map( A1 => n40611, A2 => n47573, B1 => n41715, B2 => 
                           n47543, ZN => n36865);
   U1104 : OAI22_X1 port map( A1 => n40636, A2 => n47573, B1 => n41714, B2 => 
                           n47542, ZN => n36867);
   U1105 : OAI22_X1 port map( A1 => n40623, A2 => n47568, B1 => n41713, B2 => 
                           n47535, ZN => n36868);
   U1106 : OAI22_X1 port map( A1 => n40636, A2 => n47571, B1 => n41712, B2 => 
                           n47542, ZN => n36869);
   U1107 : OAI22_X1 port map( A1 => n40610, A2 => n47568, B1 => n41711, B2 => 
                           n47540, ZN => n36871);
   U1108 : OAI22_X1 port map( A1 => n40617, A2 => n47572, B1 => n41710, B2 => 
                           n47538, ZN => n36873);
   U1109 : OAI22_X1 port map( A1 => n40617, A2 => n47574, B1 => n41709, B2 => 
                           n47538, ZN => n36874);
   U1110 : OAI22_X1 port map( A1 => n40619, A2 => n47574, B1 => n41708, B2 => 
                           n47541, ZN => n36876);
   U1111 : OAI22_X1 port map( A1 => n40611, A2 => n47574, B1 => n41707, B2 => 
                           n47543, ZN => n36877);
   U1112 : OAI22_X1 port map( A1 => n40611, A2 => n47571, B1 => n41706, B2 => 
                           n47543, ZN => n36879);
   U1113 : OAI22_X1 port map( A1 => n40617, A2 => n47573, B1 => n41705, B2 => 
                           n47538, ZN => n36881);
   U1114 : OAI22_X1 port map( A1 => n40619, A2 => n47575, B1 => n41704, B2 => 
                           n47541, ZN => n36883);
   U1115 : OAI22_X1 port map( A1 => n40617, A2 => n47575, B1 => n41703, B2 => 
                           n47538, ZN => n36885);
   U1116 : OAI22_X1 port map( A1 => n40614, A2 => n47568, B1 => n41702, B2 => 
                           n47536, ZN => n36886);
   U1117 : OAI22_X1 port map( A1 => n40617, A2 => n47571, B1 => n41701, B2 => 
                           n47538, ZN => n36888);
   U1118 : OAI22_X1 port map( A1 => n40611, A2 => n47568, B1 => n41700, B2 => 
                           n47543, ZN => n36890);
   U1119 : OAI22_X1 port map( A1 => n40617, A2 => n47569, B1 => n41699, B2 => 
                           n47538, ZN => n36893);
   U1120 : OAI22_X1 port map( A1 => n40636, A2 => n47572, B1 => n41698, B2 => 
                           n47542, ZN => n36895);
   U1121 : OAI22_X1 port map( A1 => n40636, A2 => n47574, B1 => n41697, B2 => 
                           n47542, ZN => n36897);
   U1122 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1),
                           ZN => n30048);
   U1123 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n41694, ZN => 
                           n47583);
   U1124 : NOR2_X1 port map( A1 => n40660, A2 => n47583, ZN => n47581);
   U1125 : NAND2_X1 port map( A1 => n40561, A2 => n47581, ZN => n30124);
   U1126 : INV_X1 port map( A => ADD_WR(0), ZN => n47577);
   U1127 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n47577, ZN
                           => n30046);
   U1128 : NAND2_X1 port map( A1 => n47581, A2 => n40558, ZN => n30123);
   U1129 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n47577, ZN => n47578);
   U1130 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n47578, ZN => n30121);
   U1131 : NAND2_X1 port map( A1 => n47581, A2 => n40643, ZN => n30120);
   U1132 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n47579);
   U1133 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n47579, ZN => n30118);
   U1134 : NAND2_X1 port map( A1 => n47581, A2 => n40639, ZN => n30117);
   U1135 : INV_X1 port map( A => ADD_WR(2), ZN => n47580);
   U1136 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n47580, ZN
                           => n30044);
   U1137 : NAND2_X1 port map( A1 => n47581, A2 => n40555, ZN => n30116);
   U1138 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n47577, A3 => n47580, ZN =>
                           n30042);
   U1139 : NAND2_X1 port map( A1 => n47581, A2 => n40552, ZN => n30115);
   U1140 : NOR2_X1 port map( A1 => n47580, A2 => n47578, ZN => n30113);
   U1141 : NAND2_X1 port map( A1 => n47581, A2 => n40633, ZN => n30112);
   U1142 : NOR2_X1 port map( A1 => n47580, A2 => n47579, ZN => n30110);
   U1143 : NAND2_X1 port map( A1 => n47581, A2 => n40629, ZN => n30109);
   U1144 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n40658, ZN => 
                           n47585);
   U1145 : NOR2_X1 port map( A1 => n40660, A2 => n47585, ZN => n47582);
   U1146 : NAND2_X1 port map( A1 => n40561, A2 => n47582, ZN => n30108);
   U1147 : NAND2_X1 port map( A1 => n40558, A2 => n47582, ZN => n30107);
   U1148 : NAND2_X1 port map( A1 => n40643, A2 => n47582, ZN => n30106);
   U1149 : NAND2_X1 port map( A1 => n40639, A2 => n47582, ZN => n30105);
   U1150 : NAND2_X1 port map( A1 => n40555, A2 => n47582, ZN => n30104);
   U1151 : NAND2_X1 port map( A1 => n40552, A2 => n47582, ZN => n30103);
   U1152 : NAND2_X1 port map( A1 => n40633, A2 => n47582, ZN => n30102);
   U1153 : NAND2_X1 port map( A1 => n40629, A2 => n47582, ZN => n30101);
   U1154 : NOR2_X1 port map( A1 => n40662, A2 => n47583, ZN => n47584);
   U1155 : NAND2_X1 port map( A1 => n40561, A2 => n47584, ZN => n30100);
   U1156 : NAND2_X1 port map( A1 => n40558, A2 => n47584, ZN => n30099);
   U1157 : NAND2_X1 port map( A1 => n40643, A2 => n47584, ZN => n30098);
   U1158 : NAND2_X1 port map( A1 => n40639, A2 => n47584, ZN => n30097);
   U1159 : NAND2_X1 port map( A1 => n40555, A2 => n47584, ZN => n30096);
   U1160 : NAND2_X1 port map( A1 => n40552, A2 => n47584, ZN => n30095);
   U1161 : NAND2_X1 port map( A1 => n40633, A2 => n47584, ZN => n30094);
   U1162 : NAND2_X1 port map( A1 => n40629, A2 => n47584, ZN => n30093);
   U1163 : NOR2_X1 port map( A1 => n40662, A2 => n47585, ZN => n47586);
   U1164 : NAND2_X1 port map( A1 => n40561, A2 => n47586, ZN => n30092);
   U1165 : NAND2_X1 port map( A1 => n40558, A2 => n47586, ZN => n30091);
   U1166 : NAND2_X1 port map( A1 => n40643, A2 => n47586, ZN => n30090);
   U1167 : NAND2_X1 port map( A1 => n40639, A2 => n47586, ZN => n30089);
   U1168 : NAND2_X1 port map( A1 => n40555, A2 => n47586, ZN => n30088);
   U1169 : NAND2_X1 port map( A1 => n40552, A2 => n47586, ZN => n30087);
   U1170 : NAND2_X1 port map( A1 => n40633, A2 => n47586, ZN => n30086);
   U1171 : NAND2_X1 port map( A1 => n40629, A2 => n47586, ZN => n30085);
   U1172 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), ZN => n47589);
   U1173 : NAND2_X1 port map( A1 => ADD_RD2(2), A2 => n47589, ZN => n47495);
   U1174 : INV_X1 port map( A => ADD_RD2(3), ZN => n47587);
   U1175 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n47587, ZN => n47592);
   U1176 : NOR2_X1 port map( A1 => n47592, A2 => n47495, ZN => n30084);
   U1177 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n47591)
                           ;
   U1178 : NOR2_X1 port map( A1 => n47496, A2 => n47591, ZN => n30083);
   U1179 : NOR2_X1 port map( A1 => n47591, A2 => n1533, ZN => n30082);
   U1180 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => 
                           ADD_RD2(1), ZN => n47503);
   U1181 : NOR2_X1 port map( A1 => n47591, A2 => n47503, ZN => n30081);
   U1182 : NOR2_X1 port map( A1 => n47592, A2 => n1533, ZN => n30080);
   U1183 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n47588,
                           ZN => n47502);
   U1184 : NOR2_X1 port map( A1 => n47591, A2 => n47502, ZN => n30079);
   U1185 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n47588, A3 => n47590, ZN 
                           => n47498);
   U1186 : NOR2_X1 port map( A1 => n47591, A2 => n47498, ZN => n30078);
   U1187 : NOR2_X1 port map( A1 => n47592, A2 => n47503, ZN => n30077);
   U1188 : NAND2_X1 port map( A1 => n47589, A2 => n47588, ZN => n47500);
   U1189 : NOR2_X1 port map( A1 => n47592, A2 => n47500, ZN => n30076);
   U1190 : NOR2_X1 port map( A1 => n47495, A2 => n47591, ZN => n30075);
   U1191 : NOR2_X1 port map( A1 => n47591, A2 => n47500, ZN => n30074);
   U1192 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n47590,
                           ZN => n47497);
   U1193 : NOR2_X1 port map( A1 => n47591, A2 => n47497, ZN => n30073);
   U1194 : NOR2_X1 port map( A1 => n47592, A2 => n47497, ZN => n30072);
   U1195 : NOR2_X1 port map( A1 => n47592, A2 => n47502, ZN => n30071);
   U1196 : NOR2_X1 port map( A1 => n47592, A2 => n47496, ZN => n30070);
   U1197 : NOR2_X1 port map( A1 => n47592, A2 => n47498, ZN => n30069);
   U1198 : CLKBUF_X1 port map( A => n40589, Z => n48304);
   U1199 : AOI22_X1 port map( A1 => n40803, A2 => n49088, B1 => n41328, B2 => 
                           n48304, ZN => n47596);
   U1200 : AOI22_X1 port map( A1 => n41393, A2 => n49087, B1 => n40831, B2 => 
                           n49093, ZN => n47595);
   U1201 : AOI22_X1 port map( A1 => n40812, A2 => n40592, B1 => n40823, B2 => 
                           n49094, ZN => n47594);
   U1202 : CLKBUF_X1 port map( A => n40588, Z => n48205);
   U1203 : AOI22_X1 port map( A1 => n41332, A2 => n48205, B1 => n41329, B2 => 
                           n40591, ZN => n47593);
   U1204 : NAND4_X1 port map( A1 => n47596, A2 => n47595, A3 => n47594, A4 => 
                           n47593, ZN => n47602);
   U1205 : AOI22_X1 port map( A1 => n41331, A2 => n49085, B1 => n41326, B2 => 
                           n47428, ZN => n47600);
   U1206 : CLKBUF_X1 port map( A => n49092, Z => n47839);
   U1207 : CLKBUF_X1 port map( A => n47429, Z => n48228);
   U1208 : AOI22_X1 port map( A1 => n40789, A2 => n47839, B1 => n41330, B2 => 
                           n48228, ZN => n47599);
   U1209 : CLKBUF_X1 port map( A => n49090, Z => n48299);
   U1210 : AOI22_X1 port map( A1 => n41327, A2 => n48299, B1 => n41333, B2 => 
                           n49086, ZN => n47598);
   U1211 : AOI22_X1 port map( A1 => n41325, A2 => n49091, B1 => n40808, B2 => 
                           n49089, ZN => n47597);
   U1212 : NAND4_X1 port map( A1 => n47600, A2 => n47599, A3 => n47598, A4 => 
                           n47597, ZN => n47601);
   U1213 : NOR2_X1 port map( A1 => n47602, A2 => n47601, ZN => n47614);
   U1214 : NOR3_X1 port map( A1 => n40657, A2 => n42755, A3 => n48133, ZN => 
                           n48062);
   U1215 : CLKBUF_X1 port map( A => n48062, Z => n48108);
   U1216 : CLKBUF_X1 port map( A => n49076, Z => n48314);
   U1217 : AOI22_X1 port map( A1 => n40664, A2 => n49082, B1 => n40676, B2 => 
                           n48314, ZN => n47606);
   U1218 : CLKBUF_X1 port map( A => n40565, Z => n48316);
   U1219 : AOI22_X1 port map( A1 => n40663, A2 => n49079, B1 => n40670, B2 => 
                           n48316, ZN => n47605);
   U1220 : CLKBUF_X1 port map( A => n49078, Z => n48322);
   U1221 : AOI22_X1 port map( A1 => n40665, A2 => n49077, B1 => n40672, B2 => 
                           n48322, ZN => n47604);
   U1222 : INV_X1 port map( A => n47449, ZN => n48312);
   U1223 : INV_X1 port map( A => n47432, ZN => n48313);
   U1224 : AOI22_X1 port map( A1 => n40673, A2 => n48312, B1 => n40671, B2 => 
                           n48313, ZN => n47603);
   U1225 : NAND4_X1 port map( A1 => n47606, A2 => n47605, A3 => n47604, A4 => 
                           n47603, ZN => n47612);
   U1226 : NOR3_X1 port map( A1 => n42755, A2 => n42721, A3 => n48133, ZN => 
                           n47835);
   U1227 : CLKBUF_X1 port map( A => n47835, Z => n48329);
   U1228 : CLKBUF_X1 port map( A => n48313, Z => n48259);
   U1229 : AOI22_X1 port map( A1 => n41008, A2 => n48259, B1 => n41322, B2 => 
                           n49082, ZN => n47610);
   U1230 : CLKBUF_X1 port map( A => n49079, Z => n48323);
   U1231 : AOI22_X1 port map( A1 => n41320, A2 => n48322, B1 => n41321, B2 => 
                           n48323, ZN => n47609);
   U1232 : CLKBUF_X1 port map( A => n49077, Z => n48315);
   U1233 : AOI22_X1 port map( A1 => n41691, A2 => n41027, B1 => n41338, B2 => 
                           n48315, ZN => n47608);
   U1234 : AOI22_X1 port map( A1 => n41123, A2 => n49080, B1 => n40989, B2 => 
                           n49076, ZN => n47607);
   U1235 : NAND4_X1 port map( A1 => n47610, A2 => n47609, A3 => n47608, A4 => 
                           n47607, ZN => n47611);
   U1236 : AOI22_X1 port map( A1 => n48108, A2 => n47612, B1 => n48329, B2 => 
                           n47611, ZN => n47613);
   U1237 : OAI21_X1 port map( B1 => n48133, B2 => n47614, A => n47613, ZN => 
                           OUT2(31));
   U1238 : CLKBUF_X1 port map( A => n49088, Z => n48273);
   U1239 : AOI22_X1 port map( A1 => n47429, A2 => n41508, B1 => n41091, B2 => 
                           n48273, ZN => n47618);
   U1240 : AOI22_X1 port map( A1 => n48205, A2 => n41281, B1 => n40591, B2 => 
                           n41279, ZN => n47617);
   U1241 : CLKBUF_X1 port map( A => n47428, Z => n48252);
   U1242 : CLKBUF_X1 port map( A => n49094, Z => n48087);
   U1243 : AOI22_X1 port map( A1 => n48252, A2 => n41496, B1 => n41103, B2 => 
                           n48087, ZN => n47616);
   U1244 : CLKBUF_X1 port map( A => n49089, Z => n47769);
   U1245 : AOI22_X1 port map( A1 => n41062, A2 => n40592, B1 => n41075, B2 => 
                           n47769, ZN => n47615);
   U1246 : NAND4_X1 port map( A1 => n47618, A2 => n47617, A3 => n47616, A4 => 
                           n47615, ZN => n47624);
   U1247 : AOI22_X1 port map( A1 => n41394, A2 => n49087, B1 => n41098, B2 => 
                           n47839, ZN => n47622);
   U1248 : CLKBUF_X1 port map( A => n49086, Z => n48041);
   U1249 : AOI22_X1 port map( A1 => n41278, A2 => n48304, B1 => n41284, B2 => 
                           n48041, ZN => n47621);
   U1250 : AOI22_X1 port map( A1 => n41493, A2 => n49093, B1 => n41280, B2 => 
                           n49085, ZN => n47620);
   U1251 : AOI22_X1 port map( A1 => n41276, A2 => n49090, B1 => n41283, B2 => 
                           n49091, ZN => n47619);
   U1252 : NAND4_X1 port map( A1 => n47622, A2 => n47621, A3 => n47620, A4 => 
                           n47619, ZN => n47623);
   U1253 : NOR2_X1 port map( A1 => n47624, A2 => n47623, ZN => n47636);
   U1254 : AOI22_X1 port map( A1 => n41500, A2 => n49078, B1 => n41066, B2 => 
                           n49076, ZN => n47628);
   U1255 : AOI22_X1 port map( A1 => n41087, A2 => n49081, B1 => n41503, B2 => 
                           n48315, ZN => n47627);
   U1256 : AOI22_X1 port map( A1 => n41497, A2 => n49080, B1 => n41498, B2 => 
                           n49082, ZN => n47626);
   U1257 : CLKBUF_X1 port map( A => n49079, Z => n48285);
   U1258 : AOI22_X1 port map( A1 => n41523, A2 => n41691, B1 => n41499, B2 => 
                           n48285, ZN => n47625);
   U1259 : NAND4_X1 port map( A1 => n47628, A2 => n47627, A3 => n47626, A4 => 
                           n47625, ZN => n47634);
   U1260 : AOI22_X1 port map( A1 => n41104, A2 => n49080, B1 => n41040, B2 => 
                           n49076, ZN => n47632);
   U1261 : AOI22_X1 port map( A1 => n41047, A2 => n48259, B1 => n41275, B2 => 
                           n49082, ZN => n47631);
   U1262 : CLKBUF_X1 port map( A => n49078, Z => n48290);
   U1263 : AOI22_X1 port map( A1 => n40565, A2 => n41054, B1 => n41309, B2 => 
                           n48290, ZN => n47630);
   U1264 : AOI22_X1 port map( A1 => n41337, A2 => n49077, B1 => n41513, B2 => 
                           n48285, ZN => n47629);
   U1265 : NAND4_X1 port map( A1 => n47632, A2 => n47631, A3 => n47630, A4 => 
                           n47629, ZN => n47633);
   U1266 : AOI22_X1 port map( A1 => n48108, A2 => n47634, B1 => n48329, B2 => 
                           n47633, ZN => n47635);
   U1267 : OAI21_X1 port map( B1 => n48133, B2 => n47636, A => n47635, ZN => 
                           OUT2(30));
   U1268 : AOI22_X1 port map( A1 => n40693, A2 => n49094, B1 => n40746, B2 => 
                           n47839, ZN => n47640);
   U1269 : CLKBUF_X1 port map( A => n49091, Z => n47792);
   U1270 : AOI22_X1 port map( A1 => n41395, A2 => n49087, B1 => n41301, B2 => 
                           n47792, ZN => n47639);
   U1271 : AOI22_X1 port map( A1 => n48304, A2 => n41289, B1 => n40588, B2 => 
                           n41293, ZN => n47638);
   U1272 : CLKBUF_X1 port map( A => n40592, Z => n48305);
   U1273 : AOI22_X1 port map( A1 => n48228, A2 => n41291, B1 => n48305, B2 => 
                           n40759, ZN => n47637);
   U1274 : NAND4_X1 port map( A1 => n47640, A2 => n47639, A3 => n47638, A4 => 
                           n47637, ZN => n47646);
   U1275 : AOI22_X1 port map( A1 => n41295, A2 => n49086, B1 => n40682, B2 => 
                           n47769, ZN => n47644);
   U1276 : AOI22_X1 port map( A1 => n47428, A2 => n41302, B1 => n40591, B2 => 
                           n41290, ZN => n47643);
   U1277 : AOI22_X1 port map( A1 => n40814, A2 => n49093, B1 => n41288, B2 => 
                           n49090, ZN => n47642);
   U1278 : CLKBUF_X1 port map( A => n49085, Z => n47819);
   U1279 : AOI22_X1 port map( A1 => n40719, A2 => n49088, B1 => n41292, B2 => 
                           n47819, ZN => n47641);
   U1280 : NAND4_X1 port map( A1 => n47644, A2 => n47643, A3 => n47642, A4 => 
                           n47641, ZN => n47645);
   U1281 : NOR2_X1 port map( A1 => n47646, A2 => n47645, ZN => n47658);
   U1282 : AOI22_X1 port map( A1 => n40787, A2 => n49078, B1 => n40788, B2 => 
                           n48285, ZN => n47650);
   U1283 : CLKBUF_X1 port map( A => n48312, Z => n48192);
   U1284 : AOI22_X1 port map( A1 => n40792, A2 => n41691, B1 => n40791, B2 => 
                           n48192, ZN => n47649);
   U1285 : AOI22_X1 port map( A1 => n40668, A2 => n48259, B1 => n40669, B2 => 
                           n49076, ZN => n47648);
   U1286 : AOI22_X1 port map( A1 => n40786, A2 => n48315, B1 => n40790, B2 => 
                           n49082, ZN => n47647);
   U1287 : NAND4_X1 port map( A1 => n47650, A2 => n47649, A3 => n47648, A4 => 
                           n47647, ZN => n47656);
   U1288 : AOI22_X1 port map( A1 => n41336, A2 => n48315, B1 => n41296, B2 => 
                           n48285, ZN => n47654);
   U1289 : AOI22_X1 port map( A1 => n40995, A2 => n48314, B1 => n41421, B2 => 
                           n49082, ZN => n47653);
   U1290 : AOI22_X1 port map( A1 => n40565, A2 => n40996, B1 => n41310, B2 => 
                           n48290, ZN => n47652);
   U1291 : AOI22_X1 port map( A1 => n41006, A2 => n49081, B1 => n41107, B2 => 
                           n48312, ZN => n47651);
   U1292 : NAND4_X1 port map( A1 => n47654, A2 => n47653, A3 => n47652, A4 => 
                           n47651, ZN => n47655);
   U1293 : AOI22_X1 port map( A1 => n48108, A2 => n47656, B1 => n48329, B2 => 
                           n47655, ZN => n47657);
   U1294 : OAI21_X1 port map( B1 => n48133, B2 => n47658, A => n47657, ZN => 
                           OUT2(29));
   U1295 : AOI22_X1 port map( A1 => n41265, A2 => n49090, B1 => n41263, B2 => 
                           n47792, ZN => n47662);
   U1296 : AOI22_X1 port map( A1 => n41253, A2 => n40591, B1 => n41076, B2 => 
                           n47769, ZN => n47661);
   U1297 : AOI22_X1 port map( A1 => n47428, A2 => n41519, B1 => n41402, B2 => 
                           n49087, ZN => n47660);
   U1298 : AOI22_X1 port map( A1 => n48228, A2 => n41516, B1 => n41084, B2 => 
                           n48273, ZN => n47659);
   U1299 : NAND4_X1 port map( A1 => n47662, A2 => n47661, A3 => n47660, A4 => 
                           n47659, ZN => n47668);
   U1300 : AOI22_X1 port map( A1 => n41252, A2 => n40589, B1 => n41282, B2 => 
                           n48041, ZN => n47666);
   U1301 : AOI22_X1 port map( A1 => n41259, A2 => n40588, B1 => n41258, B2 => 
                           n47819, ZN => n47665);
   U1302 : AOI22_X1 port map( A1 => n41063, A2 => n48305, B1 => n41518, B2 => 
                           n49093, ZN => n47664);
   U1303 : AOI22_X1 port map( A1 => n41094, A2 => n49094, B1 => n41083, B2 => 
                           n47839, ZN => n47663);
   U1304 : NAND4_X1 port map( A1 => n47666, A2 => n47665, A3 => n47664, A4 => 
                           n47663, ZN => n47667);
   U1305 : NOR2_X1 port map( A1 => n47668, A2 => n47667, ZN => n47680);
   U1306 : AOI22_X1 port map( A1 => n41088, A2 => n49081, B1 => n41506, B2 => 
                           n49082, ZN => n47672);
   U1307 : AOI22_X1 port map( A1 => n41511, A2 => n49080, B1 => n41502, B2 => 
                           n48315, ZN => n47671);
   U1308 : AOI22_X1 port map( A1 => n41512, A2 => n40565, B1 => n41067, B2 => 
                           n48314, ZN => n47670);
   U1309 : AOI22_X1 port map( A1 => n41504, A2 => n48290, B1 => n41505, B2 => 
                           n49079, ZN => n47669);
   U1310 : NAND4_X1 port map( A1 => n47672, A2 => n47671, A3 => n47670, A4 => 
                           n47669, ZN => n47678);
   U1311 : AOI22_X1 port map( A1 => n41055, A2 => n41691, B1 => n41311, B2 => 
                           n48290, ZN => n47676);
   U1312 : AOI22_X1 port map( A1 => n41048, A2 => n49081, B1 => n41335, B2 => 
                           n48315, ZN => n47675);
   U1313 : AOI22_X1 port map( A1 => n41119, A2 => n49080, B1 => n41261, B2 => 
                           n49082, ZN => n47674);
   U1314 : CLKBUF_X1 port map( A => n49076, Z => n48321);
   U1315 : AOI22_X1 port map( A1 => n41517, A2 => n48285, B1 => n41070, B2 => 
                           n48321, ZN => n47673);
   U1316 : NAND4_X1 port map( A1 => n47676, A2 => n47675, A3 => n47674, A4 => 
                           n47673, ZN => n47677);
   U1317 : AOI22_X1 port map( A1 => n48108, A2 => n47678, B1 => n48329, B2 => 
                           n47677, ZN => n47679);
   U1318 : OAI21_X1 port map( B1 => n48133, B2 => n47680, A => n47679, ZN => 
                           OUT2(28));
   U1319 : CLKBUF_X1 port map( A => n40591, Z => n48274);
   U1320 : CLKBUF_X1 port map( A => n49087, Z => n47884);
   U1321 : AOI22_X1 port map( A1 => n41266, A2 => n48274, B1 => n41403, B2 => 
                           n47884, ZN => n47684);
   U1322 : AOI22_X1 port map( A1 => n41514, A2 => n48252, B1 => n41079, B2 => 
                           n47839, ZN => n47683);
   U1323 : AOI22_X1 port map( A1 => n41268, A2 => n48205, B1 => n41267, B2 => 
                           n47819, ZN => n47682);
   U1324 : AOI22_X1 port map( A1 => n41085, A2 => n49094, B1 => n41077, B2 => 
                           n47769, ZN => n47681);
   U1325 : NAND4_X1 port map( A1 => n47684, A2 => n47683, A3 => n47682, A4 => 
                           n47681, ZN => n47690);
   U1326 : AOI22_X1 port map( A1 => n40589, A2 => n41273, B1 => n40592, B2 => 
                           n41064, ZN => n47688);
   U1327 : AOI22_X1 port map( A1 => n47429, A2 => n41509, B1 => n41269, B2 => 
                           n48041, ZN => n47687);
   U1328 : AOI22_X1 port map( A1 => n41096, A2 => n49088, B1 => n41271, B2 => 
                           n47792, ZN => n47686);
   U1329 : AOI22_X1 port map( A1 => n41515, A2 => n49093, B1 => n41272, B2 => 
                           n49090, ZN => n47685);
   U1330 : NAND4_X1 port map( A1 => n47688, A2 => n47687, A3 => n47686, A4 => 
                           n47685, ZN => n47689);
   U1331 : NOR2_X1 port map( A1 => n47690, A2 => n47689, ZN => n47702);
   U1332 : AOI22_X1 port map( A1 => n41522, A2 => n49078, B1 => n41525, B2 => 
                           n49082, ZN => n47694);
   U1333 : AOI22_X1 port map( A1 => n41071, A2 => n49081, B1 => n41524, B2 => 
                           n49079, ZN => n47693);
   U1334 : AOI22_X1 port map( A1 => n41535, A2 => n49080, B1 => n41068, B2 => 
                           n48321, ZN => n47692);
   U1335 : AOI22_X1 port map( A1 => n41527, A2 => n41691, B1 => n41520, B2 => 
                           n49077, ZN => n47691);
   U1336 : NAND4_X1 port map( A1 => n47694, A2 => n47693, A3 => n47692, A4 => 
                           n47691, ZN => n47700);
   U1337 : AOI22_X1 port map( A1 => n41056, A2 => n40565, B1 => n41041, B2 => 
                           n48314, ZN => n47698);
   U1338 : AOI22_X1 port map( A1 => n41521, A2 => n48323, B1 => n41270, B2 => 
                           n49082, ZN => n47697);
   U1339 : AOI22_X1 port map( A1 => n41049, A2 => n49081, B1 => n41312, B2 => 
                           n49078, ZN => n47696);
   U1340 : CLKBUF_X1 port map( A => n49077, Z => n48235);
   U1341 : AOI22_X1 port map( A1 => n41105, A2 => n49080, B1 => n41334, B2 => 
                           n48235, ZN => n47695);
   U1342 : NAND4_X1 port map( A1 => n47698, A2 => n47697, A3 => n47696, A4 => 
                           n47695, ZN => n47699);
   U1343 : AOI22_X1 port map( A1 => n48108, A2 => n47700, B1 => n47835, B2 => 
                           n47699, ZN => n47701);
   U1344 : OAI21_X1 port map( B1 => n48133, B2 => n47702, A => n47701, ZN => 
                           OUT2(27));
   U1345 : AOI22_X1 port map( A1 => n41404, A2 => n49087, B1 => n41239, B2 => 
                           n47819, ZN => n47706);
   U1346 : AOI22_X1 port map( A1 => n40739, A2 => n40592, B1 => n40720, B2 => 
                           n48273, ZN => n47705);
   U1347 : AOI22_X1 port map( A1 => n47428, A2 => n41234, B1 => n40591, B2 => 
                           n41237, ZN => n47704);
   U1348 : AOI22_X1 port map( A1 => n41249, A2 => n49086, B1 => n40681, B2 => 
                           n47769, ZN => n47703);
   U1349 : NAND4_X1 port map( A1 => n47706, A2 => n47705, A3 => n47704, A4 => 
                           n47703, ZN => n47712);
   U1350 : CLKBUF_X1 port map( A => n49093, Z => n47907);
   U1351 : AOI22_X1 port map( A1 => n41236, A2 => n40589, B1 => n40813, B2 => 
                           n47907, ZN => n47710);
   U1352 : AOI22_X1 port map( A1 => n40687, A2 => n49094, B1 => n40758, B2 => 
                           n47839, ZN => n47709);
   U1353 : AOI22_X1 port map( A1 => n41235, A2 => n49090, B1 => n41233, B2 => 
                           n47792, ZN => n47708);
   U1354 : AOI22_X1 port map( A1 => n47429, A2 => n41238, B1 => n48205, B2 => 
                           n41241, ZN => n47707);
   U1355 : NAND4_X1 port map( A1 => n47710, A2 => n47709, A3 => n47708, A4 => 
                           n47707, ZN => n47711);
   U1356 : NOR2_X1 port map( A1 => n47712, A2 => n47711, ZN => n47724);
   U1357 : AOI22_X1 port map( A1 => n40805, A2 => n49080, B1 => n40794, B2 => 
                           n48235, ZN => n47716);
   U1358 : AOI22_X1 port map( A1 => n40804, A2 => n40565, B1 => n40667, B2 => 
                           n48314, ZN => n47715);
   U1359 : AOI22_X1 port map( A1 => n40793, A2 => n49078, B1 => n40806, B2 => 
                           n49082, ZN => n47714);
   U1360 : AOI22_X1 port map( A1 => n40675, A2 => n49081, B1 => n40807, B2 => 
                           n49079, ZN => n47713);
   U1361 : NAND4_X1 port map( A1 => n47716, A2 => n47715, A3 => n47714, A4 => 
                           n47713, ZN => n47722);
   U1362 : AOI22_X1 port map( A1 => n41020, A2 => n41691, B1 => n41115, B2 => 
                           n48312, ZN => n47720);
   U1363 : AOI22_X1 port map( A1 => n41313, A2 => n48322, B1 => n41230, B2 => 
                           n49082, ZN => n47719);
   U1364 : AOI22_X1 port map( A1 => n41021, A2 => n49081, B1 => n40998, B2 => 
                           n48314, ZN => n47718);
   U1365 : AOI22_X1 port map( A1 => n41324, A2 => n48235, B1 => n41274, B2 => 
                           n49079, ZN => n47717);
   U1366 : NAND4_X1 port map( A1 => n47720, A2 => n47719, A3 => n47718, A4 => 
                           n47717, ZN => n47721);
   U1367 : AOI22_X1 port map( A1 => n48108, A2 => n47722, B1 => n47835, B2 => 
                           n47721, ZN => n47723);
   U1368 : OAI21_X1 port map( B1 => n48133, B2 => n47724, A => n47723, ZN => 
                           OUT2(26));
   U1369 : AOI22_X1 port map( A1 => n41097, A2 => n49088, B1 => n41080, B2 => 
                           n47839, ZN => n47728);
   U1370 : AOI22_X1 port map( A1 => n47429, A2 => n41533, B1 => n48305, B2 => 
                           n41065, ZN => n47727);
   U1371 : AOI22_X1 port map( A1 => n41350, A2 => n49086, B1 => n41220, B2 => 
                           n49090, ZN => n47726);
   U1372 : AOI22_X1 port map( A1 => n48252, A2 => n41532, B1 => n48274, B2 => 
                           n41222, ZN => n47725);
   U1373 : NAND4_X1 port map( A1 => n47728, A2 => n47727, A3 => n47726, A4 => 
                           n47725, ZN => n47734);
   U1374 : AOI22_X1 port map( A1 => n41405, A2 => n49087, B1 => n41351, B2 => 
                           n47819, ZN => n47732);
   U1375 : AOI22_X1 port map( A1 => n41102, A2 => n49094, B1 => n41078, B2 => 
                           n47769, ZN => n47731);
   U1376 : AOI22_X1 port map( A1 => n41349, A2 => n40588, B1 => n41531, B2 => 
                           n47907, ZN => n47730);
   U1377 : AOI22_X1 port map( A1 => n41221, A2 => n48304, B1 => n41219, B2 => 
                           n47792, ZN => n47729);
   U1378 : NAND4_X1 port map( A1 => n47732, A2 => n47731, A3 => n47730, A4 => 
                           n47729, ZN => n47733);
   U1379 : NOR2_X1 port map( A1 => n47734, A2 => n47733, ZN => n47746);
   U1380 : INV_X1 port map( A => n47453, ZN => n48264);
   U1381 : CLKBUF_X1 port map( A => n48264, Z => n47984);
   U1382 : AOI22_X1 port map( A1 => n41479, A2 => n41691, B1 => n41526, B2 => 
                           n47984, ZN => n47738);
   U1383 : AOI22_X1 port map( A1 => n41090, A2 => n49081, B1 => n41489, B2 => 
                           n48192, ZN => n47737);
   U1384 : AOI22_X1 port map( A1 => n41528, A2 => n49079, B1 => n41069, B2 => 
                           n49076, ZN => n47736);
   U1385 : AOI22_X1 port map( A1 => n41534, A2 => n49078, B1 => n41529, B2 => 
                           n48235, ZN => n47735);
   U1386 : NAND4_X1 port map( A1 => n47738, A2 => n47737, A3 => n47736, A4 => 
                           n47735, ZN => n47744);
   U1387 : AOI22_X1 port map( A1 => n41050, A2 => n49081, B1 => n41424, B2 => 
                           n48290, ZN => n47742);
   U1388 : AOI22_X1 port map( A1 => n41510, A2 => n48323, B1 => n41043, B2 => 
                           n48321, ZN => n47741);
   U1389 : AOI22_X1 port map( A1 => n40565, A2 => n41057, B1 => n41108, B2 => 
                           n48312, ZN => n47740);
   U1390 : AOI22_X1 port map( A1 => n41372, A2 => n48235, B1 => n41277, B2 => 
                           n47984, ZN => n47739);
   U1391 : NAND4_X1 port map( A1 => n47742, A2 => n47741, A3 => n47740, A4 => 
                           n47739, ZN => n47743);
   U1392 : AOI22_X1 port map( A1 => n48108, A2 => n47744, B1 => n47835, B2 => 
                           n47743, ZN => n47745);
   U1393 : OAI21_X1 port map( B1 => n48133, B2 => n47746, A => n47745, ZN => 
                           OUT2(25));
   U1394 : AOI22_X1 port map( A1 => n41418, A2 => n49086, B1 => n41399, B2 => 
                           n49090, ZN => n47750);
   U1395 : AOI22_X1 port map( A1 => n40591, A2 => n41397, B1 => n40592, B2 => 
                           n40751, ZN => n47749);
   U1396 : AOI22_X1 port map( A1 => n40773, A2 => n49093, B1 => n40679, B2 => 
                           n47769, ZN => n47748);
   U1397 : AOI22_X1 port map( A1 => n40686, A2 => n49094, B1 => n40721, B2 => 
                           n49088, ZN => n47747);
   U1398 : NAND4_X1 port map( A1 => n47750, A2 => n47749, A3 => n47748, A4 => 
                           n47747, ZN => n47756);
   U1399 : AOI22_X1 port map( A1 => n41396, A2 => n49085, B1 => n40743, B2 => 
                           n47839, ZN => n47754);
   U1400 : AOI22_X1 port map( A1 => n48252, A2 => n41400, B1 => n40589, B2 => 
                           n41398, ZN => n47753);
   U1401 : AOI22_X1 port map( A1 => n48228, A2 => n41148, B1 => n41426, B2 => 
                           n47884, ZN => n47752);
   U1402 : AOI22_X1 port map( A1 => n41419, A2 => n40588, B1 => n41401, B2 => 
                           n47792, ZN => n47751);
   U1403 : NAND4_X1 port map( A1 => n47754, A2 => n47753, A3 => n47752, A4 => 
                           n47751, ZN => n47755);
   U1404 : NOR2_X1 port map( A1 => n47756, A2 => n47755, ZN => n47768);
   U1405 : AOI22_X1 port map( A1 => n48316, A2 => n40775, B1 => n40666, B2 => 
                           n48259, ZN => n47760);
   U1406 : AOI22_X1 port map( A1 => n40774, A2 => n49080, B1 => n40771, B2 => 
                           n48290, ZN => n47759);
   U1407 : AOI22_X1 port map( A1 => n40776, A2 => n49077, B1 => n40772, B2 => 
                           n49079, ZN => n47758);
   U1408 : AOI22_X1 port map( A1 => n40674, A2 => n49076, B1 => n40777, B2 => 
                           n47984, ZN => n47757);
   U1409 : NAND4_X1 port map( A1 => n47760, A2 => n47759, A3 => n47758, A4 => 
                           n47757, ZN => n47766);
   U1410 : AOI22_X1 port map( A1 => n41415, A2 => n48322, B1 => n41414, B2 => 
                           n49079, ZN => n47764);
   U1411 : AOI22_X1 port map( A1 => n48316, A2 => n41018, B1 => n40990, B2 => 
                           n48259, ZN => n47763);
   U1412 : AOI22_X1 port map( A1 => n41416, A2 => n49077, B1 => n41406, B2 => 
                           n47984, ZN => n47762);
   U1413 : AOI22_X1 port map( A1 => n41114, A2 => n49080, B1 => n41010, B2 => 
                           n48321, ZN => n47761);
   U1414 : NAND4_X1 port map( A1 => n47764, A2 => n47763, A3 => n47762, A4 => 
                           n47761, ZN => n47765);
   U1415 : AOI22_X1 port map( A1 => n48108, A2 => n47766, B1 => n47835, B2 => 
                           n47765, ZN => n47767);
   U1416 : OAI21_X1 port map( B1 => n48133, B2 => n47768, A => n47767, ZN => 
                           OUT2(24));
   U1417 : AOI22_X1 port map( A1 => n48304, A2 => n41188, B1 => n41093, B2 => 
                           n48087, ZN => n47773);
   U1418 : AOI22_X1 port map( A1 => n41092, A2 => n49088, B1 => n41147, B2 => 
                           n47792, ZN => n47772);
   U1419 : AOI22_X1 port map( A1 => n47429, A2 => n41134, B1 => n41042, B2 => 
                           n47769, ZN => n47771);
   U1420 : AOI22_X1 port map( A1 => n41166, A2 => n49090, B1 => n41081, B2 => 
                           n47839, ZN => n47770);
   U1421 : NAND4_X1 port map( A1 => n47773, A2 => n47772, A3 => n47771, A4 => 
                           n47770, ZN => n47779);
   U1422 : AOI22_X1 port map( A1 => n47428, A2 => n41154, B1 => n41053, B2 => 
                           n47907, ZN => n47777);
   U1423 : AOI22_X1 port map( A1 => n41095, A2 => n40592, B1 => n41245, B2 => 
                           n48041, ZN => n47776);
   U1424 : AOI22_X1 port map( A1 => n41133, A2 => n48274, B1 => n41135, B2 => 
                           n47819, ZN => n47775);
   U1425 : AOI22_X1 port map( A1 => n41358, A2 => n48205, B1 => n41427, B2 => 
                           n47884, ZN => n47774);
   U1426 : NAND4_X1 port map( A1 => n47777, A2 => n47776, A3 => n47775, A4 => 
                           n47774, ZN => n47778);
   U1427 : NOR2_X1 port map( A1 => n47779, A2 => n47778, ZN => n47791);
   U1428 : AOI22_X1 port map( A1 => n41474, A2 => n49078, B1 => n41490, B2 => 
                           n49076, ZN => n47783);
   U1429 : AOI22_X1 port map( A1 => n41495, A2 => n41691, B1 => n41507, B2 => 
                           n48192, ZN => n47782);
   U1430 : AOI22_X1 port map( A1 => n41494, A2 => n49081, B1 => n41476, B2 => 
                           n48323, ZN => n47781);
   U1431 : AOI22_X1 port map( A1 => n41471, A2 => n49077, B1 => n41477, B2 => 
                           n47984, ZN => n47780);
   U1432 : NAND4_X1 port map( A1 => n47783, A2 => n47782, A3 => n47781, A4 => 
                           n47780, ZN => n47789);
   U1433 : AOI22_X1 port map( A1 => n41051, A2 => n49081, B1 => n41481, B2 => 
                           n48290, ZN => n47787);
   U1434 : AOI22_X1 port map( A1 => n41058, A2 => n41691, B1 => n41472, B2 => 
                           n49079, ZN => n47786);
   U1435 : AOI22_X1 port map( A1 => n41045, A2 => n48321, B1 => n41240, B2 => 
                           n47984, ZN => n47785);
   U1436 : AOI22_X1 port map( A1 => n41121, A2 => n49080, B1 => n41323, B2 => 
                           n48235, ZN => n47784);
   U1437 : NAND4_X1 port map( A1 => n47787, A2 => n47786, A3 => n47785, A4 => 
                           n47784, ZN => n47788);
   U1438 : AOI22_X1 port map( A1 => n48108, A2 => n47789, B1 => n47835, B2 => 
                           n47788, ZN => n47790);
   U1439 : OAI21_X1 port map( B1 => n48334, B2 => n47791, A => n47790, ZN => 
                           OUT2(23));
   U1440 : AOI22_X1 port map( A1 => n41073, A2 => n40592, B1 => n41060, B2 => 
                           n49088, ZN => n47796);
   U1441 : AOI22_X1 port map( A1 => n41089, A2 => n49094, B1 => n41146, B2 => 
                           n47792, ZN => n47795);
   U1442 : AOI22_X1 port map( A1 => n40589, A2 => n41195, B1 => n40591, B2 => 
                           n41138, ZN => n47794);
   U1443 : AOI22_X1 port map( A1 => n41244, A2 => n49086, B1 => n41082, B2 => 
                           n47839, ZN => n47793);
   U1444 : NAND4_X1 port map( A1 => n47796, A2 => n47795, A3 => n47794, A4 => 
                           n47793, ZN => n47802);
   U1445 : AOI22_X1 port map( A1 => n41044, A2 => n49089, B1 => n41137, B2 => 
                           n47819, ZN => n47800);
   U1446 : AOI22_X1 port map( A1 => n47428, A2 => n41153, B1 => n41428, B2 => 
                           n47884, ZN => n47799);
   U1447 : AOI22_X1 port map( A1 => n47429, A2 => n41136, B1 => n48205, B2 => 
                           n41359, ZN => n47798);
   U1448 : AOI22_X1 port map( A1 => n41072, A2 => n49093, B1 => n41165, B2 => 
                           n49090, ZN => n47797);
   U1449 : NAND4_X1 port map( A1 => n47800, A2 => n47799, A3 => n47798, A4 => 
                           n47797, ZN => n47801);
   U1450 : NOR2_X1 port map( A1 => n47802, A2 => n47801, ZN => n47814);
   U1451 : AOI22_X1 port map( A1 => n41473, A2 => n49077, B1 => n41480, B2 => 
                           n47984, ZN => n47806);
   U1452 : AOI22_X1 port map( A1 => n41483, A2 => n41691, B1 => n41484, B2 => 
                           n48259, ZN => n47805);
   U1453 : AOI22_X1 port map( A1 => n41475, A2 => n49078, B1 => n41478, B2 => 
                           n49079, ZN => n47804);
   U1454 : AOI22_X1 port map( A1 => n41482, A2 => n49080, B1 => n41485, B2 => 
                           n48321, ZN => n47803);
   U1455 : NAND4_X1 port map( A1 => n47806, A2 => n47805, A3 => n47804, A4 => 
                           n47803, ZN => n47812);
   U1456 : AOI22_X1 port map( A1 => n41113, A2 => n49080, B1 => n41488, B2 => 
                           n49079, ZN => n47810);
   U1457 : AOI22_X1 port map( A1 => n48316, A2 => n41059, B1 => n41052, B2 => 
                           n48259, ZN => n47809);
   U1458 : AOI22_X1 port map( A1 => n41319, A2 => n48315, B1 => n41046, B2 => 
                           n48314, ZN => n47808);
   U1459 : AOI22_X1 port map( A1 => n41486, A2 => n48322, B1 => n41246, B2 => 
                           n47984, ZN => n47807);
   U1460 : NAND4_X1 port map( A1 => n47810, A2 => n47809, A3 => n47808, A4 => 
                           n47807, ZN => n47811);
   U1461 : AOI22_X1 port map( A1 => n48108, A2 => n47812, B1 => n47835, B2 => 
                           n47811, ZN => n47813);
   U1462 : OAI21_X1 port map( B1 => n48334, B2 => n47814, A => n47813, ZN => 
                           OUT2(22));
   U1463 : AOI22_X1 port map( A1 => n41353, A2 => n48274, B1 => n40722, B2 => 
                           n49088, ZN => n47818);
   U1464 : AOI22_X1 port map( A1 => n41354, A2 => n48304, B1 => n40704, B2 => 
                           n47907, ZN => n47817);
   U1465 : AOI22_X1 port map( A1 => n40685, A2 => n49094, B1 => n41429, B2 => 
                           n47884, ZN => n47816);
   U1466 : AOI22_X1 port map( A1 => n47428, A2 => n41356, B1 => n40588, B2 => 
                           n41367, ZN => n47815);
   U1467 : NAND4_X1 port map( A1 => n47818, A2 => n47817, A3 => n47816, A4 => 
                           n47815, ZN => n47825);
   U1468 : AOI22_X1 port map( A1 => n47429, A2 => n41352, B1 => n41355, B2 => 
                           n49090, ZN => n47823);
   U1469 : AOI22_X1 port map( A1 => n41366, A2 => n49086, B1 => n40715, B2 => 
                           n49089, ZN => n47822);
   U1470 : AOI22_X1 port map( A1 => n40757, A2 => n48305, B1 => n41368, B2 => 
                           n47819, ZN => n47821);
   U1471 : AOI22_X1 port map( A1 => n41357, A2 => n49091, B1 => n40737, B2 => 
                           n47839, ZN => n47820);
   U1472 : NAND4_X1 port map( A1 => n47823, A2 => n47822, A3 => n47821, A4 => 
                           n47820, ZN => n47824);
   U1473 : NOR2_X1 port map( A1 => n47825, A2 => n47824, ZN => n47838);
   U1474 : AOI22_X1 port map( A1 => n40850, A2 => n49081, B1 => n40855, B2 => 
                           n49079, ZN => n47829);
   U1475 : AOI22_X1 port map( A1 => n40857, A2 => n48235, B1 => n40848, B2 => 
                           n48321, ZN => n47828);
   U1476 : AOI22_X1 port map( A1 => n40851, A2 => n48316, B1 => n40854, B2 => 
                           n47984, ZN => n47827);
   U1477 : AOI22_X1 port map( A1 => n40853, A2 => n49080, B1 => n40856, B2 => 
                           n48290, ZN => n47826);
   U1478 : NAND4_X1 port map( A1 => n47829, A2 => n47828, A3 => n47827, A4 => 
                           n47826, ZN => n47836);
   U1479 : AOI22_X1 port map( A1 => n41364, A2 => n48322, B1 => n41363, B2 => 
                           n49079, ZN => n47833);
   U1480 : AOI22_X1 port map( A1 => n41004, A2 => n48314, B1 => n41362, B2 => 
                           n47984, ZN => n47832);
   U1481 : AOI22_X1 port map( A1 => n41015, A2 => n41691, B1 => n41031, B2 => 
                           n48259, ZN => n47831);
   U1482 : AOI22_X1 port map( A1 => n41111, A2 => n49080, B1 => n41365, B2 => 
                           n48235, ZN => n47830);
   U1483 : NAND4_X1 port map( A1 => n47833, A2 => n47832, A3 => n47831, A4 => 
                           n47830, ZN => n47834);
   U1484 : AOI22_X1 port map( A1 => n48108, A2 => n47836, B1 => n47835, B2 => 
                           n47834, ZN => n47837);
   U1485 : OAI21_X1 port map( B1 => n48334, B2 => n47838, A => n47837, ZN => 
                           OUT2(21));
   U1486 : AOI22_X1 port map( A1 => n41243, A2 => n49086, B1 => n41086, B2 => 
                           n49089, ZN => n47843);
   U1487 : AOI22_X1 port map( A1 => n41164, A2 => n49090, B1 => n41100, B2 => 
                           n47839, ZN => n47842);
   U1488 : AOI22_X1 port map( A1 => n41196, A2 => n40589, B1 => n41074, B2 => 
                           n47907, ZN => n47841);
   U1489 : AOI22_X1 port map( A1 => n41099, A2 => n49094, B1 => n41145, B2 => 
                           n49091, ZN => n47840);
   U1490 : NAND4_X1 port map( A1 => n47843, A2 => n47842, A3 => n47841, A4 => 
                           n47840, ZN => n47849);
   U1491 : AOI22_X1 port map( A1 => n41360, A2 => n40588, B1 => n41061, B2 => 
                           n49088, ZN => n47847);
   U1492 : AOI22_X1 port map( A1 => n41126, A2 => n40591, B1 => n41430, B2 => 
                           n47884, ZN => n47846);
   U1493 : AOI22_X1 port map( A1 => n48228, A2 => n41127, B1 => n41132, B2 => 
                           n49085, ZN => n47845);
   U1494 : AOI22_X1 port map( A1 => n48252, A2 => n41152, B1 => n48305, B2 => 
                           n41101, ZN => n47844);
   U1495 : NAND4_X1 port map( A1 => n47847, A2 => n47846, A3 => n47845, A4 => 
                           n47844, ZN => n47848);
   U1496 : NOR2_X1 port map( A1 => n47849, A2 => n47848, ZN => n47861);
   U1497 : AOI22_X1 port map( A1 => n41470, A2 => n41691, B1 => n41460, B2 => 
                           n48290, ZN => n47853);
   U1498 : AOI22_X1 port map( A1 => n41462, A2 => n49081, B1 => n41467, B2 => 
                           n48192, ZN => n47852);
   U1499 : AOI22_X1 port map( A1 => n41461, A2 => n48235, B1 => n41464, B2 => 
                           n49079, ZN => n47851);
   U1500 : AOI22_X1 port map( A1 => n41468, A2 => n49076, B1 => n41459, B2 => 
                           n47984, ZN => n47850);
   U1501 : NAND4_X1 port map( A1 => n47853, A2 => n47852, A3 => n47851, A4 => 
                           n47850, ZN => n47859);
   U1502 : AOI22_X1 port map( A1 => n41583, A2 => n49080, B1 => n41545, B2 => 
                           n48321, ZN => n47857);
   U1503 : AOI22_X1 port map( A1 => n41538, A2 => n49081, B1 => n41530, B2 => 
                           n48290, ZN => n47856);
   U1504 : AOI22_X1 port map( A1 => n41491, A2 => n48323, B1 => n41247, B2 => 
                           n47984, ZN => n47855);
   U1505 : AOI22_X1 port map( A1 => n40565, A2 => n41541, B1 => n41318, B2 => 
                           n48235, ZN => n47854);
   U1506 : NAND4_X1 port map( A1 => n47857, A2 => n47856, A3 => n47855, A4 => 
                           n47854, ZN => n47858);
   U1507 : AOI22_X1 port map( A1 => n48108, A2 => n47859, B1 => n48329, B2 => 
                           n47858, ZN => n47860);
   U1508 : OAI21_X1 port map( B1 => n48334, B2 => n47861, A => n47860, ZN => 
                           OUT2(20));
   U1509 : AOI22_X1 port map( A1 => n41129, A2 => n48274, B1 => n40731, B2 => 
                           n49092, ZN => n47865);
   U1510 : AOI22_X1 port map( A1 => n41197, A2 => n40589, B1 => n41431, B2 => 
                           n47884, ZN => n47864);
   U1511 : AOI22_X1 port map( A1 => n41163, A2 => n48299, B1 => n40712, B2 => 
                           n49089, ZN => n47863);
   U1512 : AOI22_X1 port map( A1 => n48228, A2 => n41130, B1 => n40683, B2 => 
                           n48087, ZN => n47862);
   U1513 : NAND4_X1 port map( A1 => n47865, A2 => n47864, A3 => n47863, A4 => 
                           n47862, ZN => n47871);
   U1514 : AOI22_X1 port map( A1 => n41242, A2 => n49086, B1 => n41131, B2 => 
                           n49085, ZN => n47869);
   U1515 : AOI22_X1 port map( A1 => n40723, A2 => n49088, B1 => n40700, B2 => 
                           n47907, ZN => n47868);
   U1516 : AOI22_X1 port map( A1 => n41361, A2 => n48205, B1 => n41144, B2 => 
                           n49091, ZN => n47867);
   U1517 : AOI22_X1 port map( A1 => n47428, A2 => n41151, B1 => n40592, B2 => 
                           n40750, ZN => n47866);
   U1518 : NAND4_X1 port map( A1 => n47869, A2 => n47868, A3 => n47867, A4 => 
                           n47866, ZN => n47870);
   U1519 : NOR2_X1 port map( A1 => n47871, A2 => n47870, ZN => n47883);
   U1520 : AOI22_X1 port map( A1 => n40865, A2 => n48316, B1 => n40837, B2 => 
                           n48321, ZN => n47875);
   U1521 : AOI22_X1 port map( A1 => n40866, A2 => n49080, B1 => n40867, B2 => 
                           n48235, ZN => n47874);
   U1522 : AOI22_X1 port map( A1 => n40868, A2 => n49079, B1 => n40852, B2 => 
                           n49082, ZN => n47873);
   U1523 : AOI22_X1 port map( A1 => n40849, A2 => n49081, B1 => n40869, B2 => 
                           n48290, ZN => n47872);
   U1524 : NAND4_X1 port map( A1 => n47875, A2 => n47874, A3 => n47873, A4 => 
                           n47872, ZN => n47881);
   U1525 : AOI22_X1 port map( A1 => n41106, A2 => n49080, B1 => n41248, B2 => 
                           n49082, ZN => n47879);
   U1526 : AOI22_X1 port map( A1 => n41285, A2 => n49079, B1 => n41012, B2 => 
                           n48321, ZN => n47878);
   U1527 : AOI22_X1 port map( A1 => n40565, A2 => n41014, B1 => n41317, B2 => 
                           n48235, ZN => n47877);
   U1528 : AOI22_X1 port map( A1 => n41017, A2 => n49081, B1 => n41339, B2 => 
                           n48290, ZN => n47876);
   U1529 : NAND4_X1 port map( A1 => n47879, A2 => n47878, A3 => n47877, A4 => 
                           n47876, ZN => n47880);
   U1530 : AOI22_X1 port map( A1 => n48108, A2 => n47881, B1 => n48329, B2 => 
                           n47880, ZN => n47882);
   U1531 : OAI21_X1 port map( B1 => n48334, B2 => n47883, A => n47882, ZN => 
                           OUT2(19));
   U1532 : AOI22_X1 port map( A1 => n41162, A2 => n48299, B1 => n41143, B2 => 
                           n49091, ZN => n47888);
   U1533 : AOI22_X1 port map( A1 => n41198, A2 => n40589, B1 => n40708, B2 => 
                           n49089, ZN => n47887);
   U1534 : AOI22_X1 port map( A1 => n47428, A2 => n41150, B1 => n41432, B2 => 
                           n47884, ZN => n47886);
   U1535 : AOI22_X1 port map( A1 => n40747, A2 => n48305, B1 => n40699, B2 => 
                           n47907, ZN => n47885);
   U1536 : NAND4_X1 port map( A1 => n47888, A2 => n47887, A3 => n47886, A4 => 
                           n47885, ZN => n47894);
   U1537 : AOI22_X1 port map( A1 => n41140, A2 => n49085, B1 => n40729, B2 => 
                           n49092, ZN => n47892);
   U1538 : AOI22_X1 port map( A1 => n40588, A2 => n41369, B1 => n40680, B2 => 
                           n48087, ZN => n47891);
   U1539 : AOI22_X1 port map( A1 => n41141, A2 => n40591, B1 => n41232, B2 => 
                           n48041, ZN => n47890);
   U1540 : AOI22_X1 port map( A1 => n47429, A2 => n41139, B1 => n40724, B2 => 
                           n49088, ZN => n47889);
   U1541 : NAND4_X1 port map( A1 => n47892, A2 => n47891, A3 => n47890, A4 => 
                           n47889, ZN => n47893);
   U1542 : NOR2_X1 port map( A1 => n47894, A2 => n47893, ZN => n47906);
   U1543 : CLKBUF_X1 port map( A => n48062, Z => n48331);
   U1544 : AOI22_X1 port map( A1 => n40860, A2 => n49080, B1 => n40862, B2 => 
                           n48323, ZN => n47898);
   U1545 : AOI22_X1 port map( A1 => n40858, A2 => n49081, B1 => n40861, B2 => 
                           n48264, ZN => n47897);
   U1546 : AOI22_X1 port map( A1 => n40863, A2 => n48290, B1 => n40864, B2 => 
                           n48235, ZN => n47896);
   U1547 : AOI22_X1 port map( A1 => n40859, A2 => n48316, B1 => n40822, B2 => 
                           n48321, ZN => n47895);
   U1548 : NAND4_X1 port map( A1 => n47898, A2 => n47897, A3 => n47896, A4 => 
                           n47895, ZN => n47904);
   U1549 : AOI22_X1 port map( A1 => n40565, A2 => n41013, B1 => n41118, B2 => 
                           n48192, ZN => n47902);
   U1550 : AOI22_X1 port map( A1 => n40993, A2 => n48321, B1 => n41250, B2 => 
                           n49082, ZN => n47901);
   U1551 : AOI22_X1 port map( A1 => n41023, A2 => n49081, B1 => n41340, B2 => 
                           n48290, ZN => n47900);
   U1552 : AOI22_X1 port map( A1 => n41316, A2 => n48235, B1 => n41286, B2 => 
                           n48323, ZN => n47899);
   U1553 : NAND4_X1 port map( A1 => n47902, A2 => n47901, A3 => n47900, A4 => 
                           n47899, ZN => n47903);
   U1554 : AOI22_X1 port map( A1 => n48331, A2 => n47904, B1 => n48329, B2 => 
                           n47903, ZN => n47905);
   U1555 : OAI21_X1 port map( B1 => n48334, B2 => n47906, A => n47905, ZN => 
                           OUT2(18));
   U1556 : AOI22_X1 port map( A1 => n40678, A2 => n49094, B1 => n40727, B2 => 
                           n49092, ZN => n47911);
   U1557 : AOI22_X1 port map( A1 => n47428, A2 => n41383, B1 => n41384, B2 => 
                           n49091, ZN => n47910);
   U1558 : AOI22_X1 port map( A1 => n40734, A2 => n49088, B1 => n41377, B2 => 
                           n49085, ZN => n47909);
   U1559 : AOI22_X1 port map( A1 => n41380, A2 => n40591, B1 => n40698, B2 => 
                           n47907, ZN => n47908);
   U1560 : NAND4_X1 port map( A1 => n47911, A2 => n47910, A3 => n47909, A4 => 
                           n47908, ZN => n47917);
   U1561 : AOI22_X1 port map( A1 => n41391, A2 => n49086, B1 => n41382, B2 => 
                           n49090, ZN => n47915);
   U1562 : AOI22_X1 port map( A1 => n48304, A2 => n41381, B1 => n40592, B2 => 
                           n40695, ZN => n47914);
   U1563 : AOI22_X1 port map( A1 => n47429, A2 => n41379, B1 => n41420, B2 => 
                           n49087, ZN => n47913);
   U1564 : AOI22_X1 port map( A1 => n41392, A2 => n40588, B1 => n40702, B2 => 
                           n49089, ZN => n47912);
   U1565 : NAND4_X1 port map( A1 => n47915, A2 => n47914, A3 => n47913, A4 => 
                           n47912, ZN => n47916);
   U1566 : NOR2_X1 port map( A1 => n47917, A2 => n47916, ZN => n47929);
   U1567 : AOI22_X1 port map( A1 => n40935, A2 => n49077, B1 => n40939, B2 => 
                           n48323, ZN => n47921);
   U1568 : AOI22_X1 port map( A1 => n48316, A2 => n40938, B1 => n40929, B2 => 
                           n48192, ZN => n47920);
   U1569 : AOI22_X1 port map( A1 => n40830, A2 => n49076, B1 => n40931, B2 => 
                           n49082, ZN => n47919);
   U1570 : AOI22_X1 port map( A1 => n40937, A2 => n49081, B1 => n40933, B2 => 
                           n48290, ZN => n47918);
   U1571 : NAND4_X1 port map( A1 => n47921, A2 => n47920, A3 => n47919, A4 => 
                           n47918, ZN => n47927);
   U1572 : AOI22_X1 port map( A1 => n41390, A2 => n49077, B1 => n41387, B2 => 
                           n49082, ZN => n47925);
   U1573 : AOI22_X1 port map( A1 => n41584, A2 => n49080, B1 => n41557, B2 => 
                           n48321, ZN => n47924);
   U1574 : AOI22_X1 port map( A1 => n41539, A2 => n49081, B1 => n41389, B2 => 
                           n48290, ZN => n47923);
   U1575 : AOI22_X1 port map( A1 => n41542, A2 => n40565, B1 => n41388, B2 => 
                           n48323, ZN => n47922);
   U1576 : NAND4_X1 port map( A1 => n47925, A2 => n47924, A3 => n47923, A4 => 
                           n47922, ZN => n47926);
   U1577 : AOI22_X1 port map( A1 => n48331, A2 => n47927, B1 => n48329, B2 => 
                           n47926, ZN => n47928);
   U1578 : OAI21_X1 port map( B1 => n48334, B2 => n47929, A => n47928, ZN => 
                           OUT2(17));
   U1579 : AOI22_X1 port map( A1 => n40697, A2 => n49093, B1 => n41438, B2 => 
                           n49085, ZN => n47933);
   U1580 : AOI22_X1 port map( A1 => n41437, A2 => n47429, B1 => n40726, B2 => 
                           n49092, ZN => n47932);
   U1581 : AOI22_X1 port map( A1 => n41422, A2 => n48299, B1 => n41425, B2 => 
                           n49091, ZN => n47931);
   U1582 : AOI22_X1 port map( A1 => n40592, A2 => n40754, B1 => n40728, B2 => 
                           n48087, ZN => n47930);
   U1583 : NAND4_X1 port map( A1 => n47933, A2 => n47932, A3 => n47931, A4 => 
                           n47930, ZN => n47939);
   U1584 : AOI22_X1 port map( A1 => n41413, A2 => n48205, B1 => n40736, B2 => 
                           n49088, ZN => n47937);
   U1585 : AOI22_X1 port map( A1 => n41417, A2 => n40591, B1 => n40694, B2 => 
                           n49089, ZN => n47936);
   U1586 : AOI22_X1 port map( A1 => n48252, A2 => n41423, B1 => n48304, B2 => 
                           n41411, ZN => n47935);
   U1587 : AOI22_X1 port map( A1 => n41434, A2 => n49087, B1 => n41412, B2 => 
                           n48041, ZN => n47934);
   U1588 : NAND4_X1 port map( A1 => n47937, A2 => n47936, A3 => n47935, A4 => 
                           n47934, ZN => n47938);
   U1589 : NOR2_X1 port map( A1 => n47939, A2 => n47938, ZN => n47951);
   U1590 : AOI22_X1 port map( A1 => n40841, A2 => n41691, B1 => n40934, B2 => 
                           n48321, ZN => n47943);
   U1591 : AOI22_X1 port map( A1 => n40847, A2 => n49077, B1 => n40843, B2 => 
                           n49082, ZN => n47942);
   U1592 : AOI22_X1 port map( A1 => n40840, A2 => n49081, B1 => n40844, B2 => 
                           n48323, ZN => n47941);
   U1593 : AOI22_X1 port map( A1 => n40842, A2 => n49080, B1 => n40845, B2 => 
                           n48290, ZN => n47940);
   U1594 : NAND4_X1 port map( A1 => n47943, A2 => n47942, A3 => n47941, A4 => 
                           n47940, ZN => n47949);
   U1595 : AOI22_X1 port map( A1 => n41409, A2 => n49078, B1 => n41410, B2 => 
                           n48235, ZN => n47947);
   U1596 : AOI22_X1 port map( A1 => n41116, A2 => n49080, B1 => n41005, B2 => 
                           n48321, ZN => n47946);
   U1597 : AOI22_X1 port map( A1 => n41009, A2 => n48316, B1 => n41408, B2 => 
                           n48323, ZN => n47945);
   U1598 : AOI22_X1 port map( A1 => n41022, A2 => n49081, B1 => n41407, B2 => 
                           n49082, ZN => n47944);
   U1599 : NAND4_X1 port map( A1 => n47947, A2 => n47946, A3 => n47945, A4 => 
                           n47944, ZN => n47948);
   U1600 : AOI22_X1 port map( A1 => n48108, A2 => n47949, B1 => n48329, B2 => 
                           n47948, ZN => n47950);
   U1601 : OAI21_X1 port map( B1 => n48334, B2 => n47951, A => n47950, ZN => 
                           OUT2(16));
   U1602 : AOI22_X1 port map( A1 => n47429, A2 => n41174, B1 => n40589, B2 => 
                           n41199, ZN => n47955);
   U1603 : AOI22_X1 port map( A1 => n48205, A2 => n41370, B1 => n48274, B2 => 
                           n41178, ZN => n47954);
   U1604 : AOI22_X1 port map( A1 => n40677, A2 => n49094, B1 => n41173, B2 => 
                           n49085, ZN => n47953);
   U1605 : AOI22_X1 port map( A1 => n40696, A2 => n49093, B1 => n40725, B2 => 
                           n49092, ZN => n47952);
   U1606 : NAND4_X1 port map( A1 => n47955, A2 => n47954, A3 => n47953, A4 => 
                           n47952, ZN => n47961);
   U1607 : AOI22_X1 port map( A1 => n40738, A2 => n49088, B1 => n41433, B2 => 
                           n49087, ZN => n47959);
   U1608 : AOI22_X1 port map( A1 => n40749, A2 => n40592, B1 => n40701, B2 => 
                           n49089, ZN => n47958);
   U1609 : AOI22_X1 port map( A1 => n48252, A2 => n41176, B1 => n41177, B2 => 
                           n49091, ZN => n47957);
   U1610 : AOI22_X1 port map( A1 => n41231, A2 => n49086, B1 => n41175, B2 => 
                           n49090, ZN => n47956);
   U1611 : NAND4_X1 port map( A1 => n47959, A2 => n47958, A3 => n47957, A4 => 
                           n47956, ZN => n47960);
   U1612 : NOR2_X1 port map( A1 => n47961, A2 => n47960, ZN => n47973);
   U1613 : AOI22_X1 port map( A1 => n40888, A2 => n49078, B1 => n40892, B2 => 
                           n47984, ZN => n47965);
   U1614 : AOI22_X1 port map( A1 => n40904, A2 => n48313, B1 => n40882, B2 => 
                           n48192, ZN => n47964);
   U1615 : AOI22_X1 port map( A1 => n40887, A2 => n48315, B1 => n40891, B2 => 
                           n48323, ZN => n47963);
   U1616 : AOI22_X1 port map( A1 => n40893, A2 => n40565, B1 => n40799, B2 => 
                           n48321, ZN => n47962);
   U1617 : NAND4_X1 port map( A1 => n47965, A2 => n47964, A3 => n47963, A4 => 
                           n47962, ZN => n47971);
   U1618 : AOI22_X1 port map( A1 => n41540, A2 => n48259, B1 => n41554, B2 => 
                           n48321, ZN => n47969);
   U1619 : AOI22_X1 port map( A1 => n41580, A2 => n49080, B1 => n41251, B2 => 
                           n49082, ZN => n47968);
   U1620 : AOI22_X1 port map( A1 => n41341, A2 => n48290, B1 => n41315, B2 => 
                           n48235, ZN => n47967);
   U1621 : AOI22_X1 port map( A1 => n41556, A2 => n40565, B1 => n41287, B2 => 
                           n48323, ZN => n47966);
   U1622 : NAND4_X1 port map( A1 => n47969, A2 => n47968, A3 => n47967, A4 => 
                           n47966, ZN => n47970);
   U1623 : AOI22_X1 port map( A1 => n48108, A2 => n47971, B1 => n48329, B2 => 
                           n47970, ZN => n47972);
   U1624 : OAI21_X1 port map( B1 => n48334, B2 => n47973, A => n47972, ZN => 
                           OUT2(15));
   U1625 : AOI22_X1 port map( A1 => n40761, A2 => n40592, B1 => n40717, B2 => 
                           n49092, ZN => n47977);
   U1626 : AOI22_X1 port map( A1 => n41200, A2 => n48304, B1 => n41436, B2 => 
                           n49087, ZN => n47976);
   U1627 : AOI22_X1 port map( A1 => n40684, A2 => n49094, B1 => n41142, B2 => 
                           n49091, ZN => n47975);
   U1628 : AOI22_X1 port map( A1 => n48228, A2 => n41125, B1 => n41128, B2 => 
                           n49085, ZN => n47974);
   U1629 : NAND4_X1 port map( A1 => n47977, A2 => n47976, A3 => n47975, A4 => 
                           n47974, ZN => n47983);
   U1630 : AOI22_X1 port map( A1 => n41229, A2 => n49086, B1 => n40703, B2 => 
                           n49089, ZN => n47981);
   U1631 : AOI22_X1 port map( A1 => n47428, A2 => n41149, B1 => n41158, B2 => 
                           n49090, ZN => n47980);
   U1632 : AOI22_X1 port map( A1 => n40740, A2 => n48273, B1 => n40692, B2 => 
                           n49093, ZN => n47979);
   U1633 : AOI22_X1 port map( A1 => n40588, A2 => n41371, B1 => n40591, B2 => 
                           n41179, ZN => n47978);
   U1634 : NAND4_X1 port map( A1 => n47981, A2 => n47980, A3 => n47979, A4 => 
                           n47978, ZN => n47982);
   U1635 : NOR2_X1 port map( A1 => n47983, A2 => n47982, ZN => n47996);
   U1636 : AOI22_X1 port map( A1 => n40925, A2 => n48314, B1 => n40801, B2 => 
                           n47984, ZN => n47988);
   U1637 : AOI22_X1 port map( A1 => n40798, A2 => n49078, B1 => n40800, B2 => 
                           n48323, ZN => n47987);
   U1638 : AOI22_X1 port map( A1 => n40796, A2 => n48259, B1 => n40797, B2 => 
                           n48235, ZN => n47986);
   U1639 : AOI22_X1 port map( A1 => n40565, A2 => n40795, B1 => n40802, B2 => 
                           n48192, ZN => n47985);
   U1640 : NAND4_X1 port map( A1 => n47988, A2 => n47987, A3 => n47986, A4 => 
                           n47985, ZN => n47994);
   U1641 : AOI22_X1 port map( A1 => n41124, A2 => n48192, B1 => n41028, B2 => 
                           n48321, ZN => n47992);
   U1642 : AOI22_X1 port map( A1 => n41342, A2 => n49078, B1 => n41254, B2 => 
                           n49082, ZN => n47991);
   U1643 : AOI22_X1 port map( A1 => n41030, A2 => n49081, B1 => n41314, B2 => 
                           n48315, ZN => n47990);
   U1644 : AOI22_X1 port map( A1 => n41007, A2 => n40565, B1 => n41294, B2 => 
                           n48323, ZN => n47989);
   U1645 : NAND4_X1 port map( A1 => n47992, A2 => n47991, A3 => n47990, A4 => 
                           n47989, ZN => n47993);
   U1646 : AOI22_X1 port map( A1 => n48108, A2 => n47994, B1 => n48329, B2 => 
                           n47993, ZN => n47995);
   U1647 : OAI21_X1 port map( B1 => n48334, B2 => n47996, A => n47995, ZN => 
                           OUT2(14));
   U1648 : AOI22_X1 port map( A1 => n47428, A2 => n41186, B1 => n40691, B2 => 
                           n49093, ZN => n48000);
   U1649 : AOI22_X1 port map( A1 => n41228, A2 => n49086, B1 => n41187, B2 => 
                           n49091, ZN => n47999);
   U1650 : AOI22_X1 port map( A1 => n41373, A2 => n40588, B1 => n41182, B2 => 
                           n49085, ZN => n47998);
   U1651 : AOI22_X1 port map( A1 => n41201, A2 => n48304, B1 => n41435, B2 => 
                           n49087, ZN => n47997);
   U1652 : NAND4_X1 port map( A1 => n48000, A2 => n47999, A3 => n47998, A4 => 
                           n47997, ZN => n48006);
   U1653 : AOI22_X1 port map( A1 => n40762, A2 => n40592, B1 => n41185, B2 => 
                           n49090, ZN => n48004);
   U1654 : AOI22_X1 port map( A1 => n40742, A2 => n48273, B1 => n40705, B2 => 
                           n49089, ZN => n48003);
   U1655 : AOI22_X1 port map( A1 => n47429, A2 => n41183, B1 => n48274, B2 => 
                           n41184, ZN => n48002);
   U1656 : AOI22_X1 port map( A1 => n40745, A2 => n49094, B1 => n40716, B2 => 
                           n49092, ZN => n48001);
   U1657 : NAND4_X1 port map( A1 => n48004, A2 => n48003, A3 => n48002, A4 => 
                           n48001, ZN => n48005);
   U1658 : NOR2_X1 port map( A1 => n48006, A2 => n48005, ZN => n48018);
   U1659 : AOI22_X1 port map( A1 => n48316, A2 => n40817, B1 => n40810, B2 => 
                           n48322, ZN => n48010);
   U1660 : AOI22_X1 port map( A1 => n40809, A2 => n49079, B1 => n40815, B2 => 
                           n49076, ZN => n48009);
   U1661 : AOI22_X1 port map( A1 => n40818, A2 => n48312, B1 => n40819, B2 => 
                           n48264, ZN => n48008);
   U1662 : AOI22_X1 port map( A1 => n40816, A2 => n48313, B1 => n40811, B2 => 
                           n49077, ZN => n48007);
   U1663 : NAND4_X1 port map( A1 => n48010, A2 => n48009, A3 => n48008, A4 => 
                           n48007, ZN => n48016);
   U1664 : AOI22_X1 port map( A1 => n41308, A2 => n48315, B1 => n41255, B2 => 
                           n48264, ZN => n48014);
   U1665 : AOI22_X1 port map( A1 => n40994, A2 => n40565, B1 => n41011, B2 => 
                           n48321, ZN => n48013);
   U1666 : AOI22_X1 port map( A1 => n41117, A2 => n49080, B1 => n41343, B2 => 
                           n48322, ZN => n48012);
   U1667 : AOI22_X1 port map( A1 => n41001, A2 => n48313, B1 => n41297, B2 => 
                           n48285, ZN => n48011);
   U1668 : NAND4_X1 port map( A1 => n48014, A2 => n48013, A3 => n48012, A4 => 
                           n48011, ZN => n48015);
   U1669 : AOI22_X1 port map( A1 => n48108, A2 => n48016, B1 => n48329, B2 => 
                           n48015, ZN => n48017);
   U1670 : OAI21_X1 port map( B1 => n48334, B2 => n48018, A => n48017, ZN => 
                           OUT2(13));
   U1671 : AOI22_X1 port map( A1 => n41194, A2 => n49091, B1 => n40714, B2 => 
                           n49092, ZN => n48022);
   U1672 : AOI22_X1 port map( A1 => n41191, A2 => n40591, B1 => n40706, B2 => 
                           n49089, ZN => n48021);
   U1673 : AOI22_X1 port map( A1 => n41374, A2 => n48205, B1 => n41439, B2 => 
                           n49087, ZN => n48020);
   U1674 : AOI22_X1 port map( A1 => n40589, A2 => n41202, B1 => n40748, B2 => 
                           n48087, ZN => n48019);
   U1675 : NAND4_X1 port map( A1 => n48022, A2 => n48021, A3 => n48020, A4 => 
                           n48019, ZN => n48028);
   U1676 : AOI22_X1 port map( A1 => n40744, A2 => n48305, B1 => n41227, B2 => 
                           n48041, ZN => n48026);
   U1677 : AOI22_X1 port map( A1 => n48228, A2 => n41190, B1 => n41189, B2 => 
                           n49085, ZN => n48025);
   U1678 : AOI22_X1 port map( A1 => n40756, A2 => n48273, B1 => n40690, B2 => 
                           n49093, ZN => n48024);
   U1679 : AOI22_X1 port map( A1 => n47428, A2 => n41193, B1 => n41192, B2 => 
                           n49090, ZN => n48023);
   U1680 : NAND4_X1 port map( A1 => n48026, A2 => n48025, A3 => n48024, A4 => 
                           n48023, ZN => n48027);
   U1681 : NOR2_X1 port map( A1 => n48028, A2 => n48027, ZN => n48040);
   U1682 : AOI22_X1 port map( A1 => n40826, A2 => n48316, B1 => n40824, B2 => 
                           n49076, ZN => n48032);
   U1683 : AOI22_X1 port map( A1 => n40829, A2 => n48323, B1 => n40828, B2 => 
                           n48264, ZN => n48031);
   U1684 : AOI22_X1 port map( A1 => n40825, A2 => n48313, B1 => n40827, B2 => 
                           n48192, ZN => n48030);
   U1685 : AOI22_X1 port map( A1 => n40820, A2 => n49078, B1 => n40821, B2 => 
                           n49077, ZN => n48029);
   U1686 : NAND4_X1 port map( A1 => n48032, A2 => n48031, A3 => n48030, A4 => 
                           n48029, ZN => n48038);
   U1687 : AOI22_X1 port map( A1 => n41033, A2 => n48313, B1 => n41344, B2 => 
                           n48322, ZN => n48036);
   U1688 : AOI22_X1 port map( A1 => n41109, A2 => n48312, B1 => n41307, B2 => 
                           n49077, ZN => n48035);
   U1689 : AOI22_X1 port map( A1 => n41003, A2 => n48316, B1 => n41298, B2 => 
                           n48285, ZN => n48034);
   U1690 : AOI22_X1 port map( A1 => n41032, A2 => n49076, B1 => n41256, B2 => 
                           n48264, ZN => n48033);
   U1691 : NAND4_X1 port map( A1 => n48036, A2 => n48035, A3 => n48034, A4 => 
                           n48033, ZN => n48037);
   U1692 : AOI22_X1 port map( A1 => n48108, A2 => n48038, B1 => n48329, B2 => 
                           n48037, ZN => n48039);
   U1693 : OAI21_X1 port map( B1 => n48334, B2 => n48040, A => n48039, ZN => 
                           OUT2(12));
   U1694 : AOI22_X1 port map( A1 => n41206, A2 => n40589, B1 => n40732, B2 => 
                           n49088, ZN => n48045);
   U1695 : AOI22_X1 port map( A1 => n41205, A2 => n48274, B1 => n41693, B2 => 
                           n49093, ZN => n48044);
   U1696 : AOI22_X1 port map( A1 => n41378, A2 => n49087, B1 => n41226, B2 => 
                           n48041, ZN => n48043);
   U1697 : AOI22_X1 port map( A1 => n40592, A2 => n40760, B1 => n40752, B2 => 
                           n48087, ZN => n48042);
   U1698 : NAND4_X1 port map( A1 => n48045, A2 => n48044, A3 => n48043, A4 => 
                           n48042, ZN => n48051);
   U1699 : AOI22_X1 port map( A1 => n41207, A2 => n48299, B1 => n41209, B2 => 
                           n49091, ZN => n48049);
   U1700 : AOI22_X1 port map( A1 => n40707, A2 => n49089, B1 => n40713, B2 => 
                           n49092, ZN => n48048);
   U1701 : AOI22_X1 port map( A1 => n41375, A2 => n40588, B1 => n41203, B2 => 
                           n49085, ZN => n48047);
   U1702 : AOI22_X1 port map( A1 => n47429, A2 => n41204, B1 => n48252, B2 => 
                           n41208, ZN => n48046);
   U1703 : NAND4_X1 port map( A1 => n48049, A2 => n48048, A3 => n48047, A4 => 
                           n48046, ZN => n48050);
   U1704 : NOR2_X1 port map( A1 => n48051, A2 => n48050, ZN => n48064);
   U1705 : AOI22_X1 port map( A1 => n40836, A2 => n48312, B1 => n40846, B2 => 
                           n48322, ZN => n48055);
   U1706 : AOI22_X1 port map( A1 => n40832, A2 => n48315, B1 => n40839, B2 => 
                           n48285, ZN => n48054);
   U1707 : AOI22_X1 port map( A1 => n48316, A2 => n40835, B1 => n40834, B2 => 
                           n48259, ZN => n48053);
   U1708 : AOI22_X1 port map( A1 => n40833, A2 => n48314, B1 => n40838, B2 => 
                           n48264, ZN => n48052);
   U1709 : NAND4_X1 port map( A1 => n48055, A2 => n48054, A3 => n48053, A4 => 
                           n48052, ZN => n48061);
   U1710 : AOI22_X1 port map( A1 => n41110, A2 => n48312, B1 => n41257, B2 => 
                           n48264, ZN => n48059);
   U1711 : AOI22_X1 port map( A1 => n41303, A2 => n48323, B1 => n41019, B2 => 
                           n49076, ZN => n48058);
   U1712 : AOI22_X1 port map( A1 => n48316, A2 => n41002, B1 => n40999, B2 => 
                           n48259, ZN => n48057);
   U1713 : AOI22_X1 port map( A1 => n41345, A2 => n49078, B1 => n41306, B2 => 
                           n49077, ZN => n48056);
   U1714 : NAND4_X1 port map( A1 => n48059, A2 => n48058, A3 => n48057, A4 => 
                           n48056, ZN => n48060);
   U1715 : AOI22_X1 port map( A1 => n48062, A2 => n48061, B1 => n48329, B2 => 
                           n48060, ZN => n48063);
   U1716 : OAI21_X1 port map( B1 => n48133, B2 => n48064, A => n48063, ZN => 
                           OUT2(11));
   U1717 : AOI22_X1 port map( A1 => n48252, A2 => n41216, B1 => n40588, B2 => 
                           n41376, ZN => n48068);
   U1718 : AOI22_X1 port map( A1 => n40985, A2 => n49094, B1 => n40986, B2 => 
                           n49089, ZN => n48067);
   U1719 : AOI22_X1 port map( A1 => n40987, A2 => n40592, B1 => n40983, B2 => 
                           n49093, ZN => n48066);
   U1720 : AOI22_X1 port map( A1 => n41215, A2 => n48299, B1 => n41212, B2 => 
                           n49085, ZN => n48065);
   U1721 : NAND4_X1 port map( A1 => n48068, A2 => n48067, A3 => n48066, A4 => 
                           n48065, ZN => n48074);
   U1722 : AOI22_X1 port map( A1 => n41225, A2 => n49086, B1 => n41217, B2 => 
                           n49091, ZN => n48072);
   U1723 : AOI22_X1 port map( A1 => n41172, A2 => n49087, B1 => n40984, B2 => 
                           n49092, ZN => n48071);
   U1724 : AOI22_X1 port map( A1 => n48228, A2 => n41451, B1 => n40589, B2 => 
                           n41214, ZN => n48070);
   U1725 : AOI22_X1 port map( A1 => n41213, A2 => n40591, B1 => n40988, B2 => 
                           n49088, ZN => n48069);
   U1726 : NAND4_X1 port map( A1 => n48072, A2 => n48071, A3 => n48070, A4 => 
                           n48069, ZN => n48073);
   U1727 : NOR2_X1 port map( A1 => n48074, A2 => n48073, ZN => n48086);
   U1728 : AOI22_X1 port map( A1 => n48316, A2 => n41450, B1 => n41446, B2 => 
                           n48192, ZN => n48078);
   U1729 : AOI22_X1 port map( A1 => n41453, A2 => n48313, B1 => n41452, B2 => 
                           n49076, ZN => n48077);
   U1730 : AOI22_X1 port map( A1 => n41445, A2 => n49077, B1 => n41443, B2 => 
                           n48285, ZN => n48076);
   U1731 : AOI22_X1 port map( A1 => n41448, A2 => n49078, B1 => n41449, B2 => 
                           n48264, ZN => n48075);
   U1732 : NAND4_X1 port map( A1 => n48078, A2 => n48077, A3 => n48076, A4 => 
                           n48075, ZN => n48084);
   U1733 : AOI22_X1 port map( A1 => n41348, A2 => n49078, B1 => n41016, B2 => 
                           n49076, ZN => n48082);
   U1734 : AOI22_X1 port map( A1 => n41112, A2 => n48192, B1 => n41444, B2 => 
                           n48285, ZN => n48081);
   U1735 : AOI22_X1 port map( A1 => n41026, A2 => n48313, B1 => n41260, B2 => 
                           n48264, ZN => n48080);
   U1736 : AOI22_X1 port map( A1 => n40565, A2 => n40992, B1 => n41447, B2 => 
                           n49077, ZN => n48079);
   U1737 : NAND4_X1 port map( A1 => n48082, A2 => n48081, A3 => n48080, A4 => 
                           n48079, ZN => n48083);
   U1738 : AOI22_X1 port map( A1 => n48108, A2 => n48084, B1 => n48329, B2 => 
                           n48083, ZN => n48085);
   U1739 : OAI21_X1 port map( B1 => n48133, B2 => n48086, A => n48085, ZN => 
                           OUT2(10));
   U1740 : AOI22_X1 port map( A1 => n41180, A2 => n48274, B1 => n40733, B2 => 
                           n48273, ZN => n48091);
   U1741 : AOI22_X1 port map( A1 => n47428, A2 => n41169, B1 => n40753, B2 => 
                           n48087, ZN => n48090);
   U1742 : AOI22_X1 port map( A1 => n41170, A2 => n48299, B1 => n40711, B2 => 
                           n49092, ZN => n48089);
   U1743 : AOI22_X1 port map( A1 => n41218, A2 => n49091, B1 => n41167, B2 => 
                           n49085, ZN => n48088);
   U1744 : NAND4_X1 port map( A1 => n48091, A2 => n48090, A3 => n48089, A4 => 
                           n48088, ZN => n48097);
   U1745 : AOI22_X1 port map( A1 => n40741, A2 => n40592, B1 => n40689, B2 => 
                           n49093, ZN => n48095);
   U1746 : AOI22_X1 port map( A1 => n41224, A2 => n49086, B1 => n40709, B2 => 
                           n49089, ZN => n48094);
   U1747 : AOI22_X1 port map( A1 => n48228, A2 => n41171, B1 => n40588, B2 => 
                           n41385, ZN => n48093);
   U1748 : AOI22_X1 port map( A1 => n41210, A2 => n40589, B1 => n41168, B2 => 
                           n49087, ZN => n48092);
   U1749 : NAND4_X1 port map( A1 => n48095, A2 => n48094, A3 => n48093, A4 => 
                           n48092, ZN => n48096);
   U1750 : NOR2_X1 port map( A1 => n48097, A2 => n48096, ZN => n48110);
   U1751 : AOI22_X1 port map( A1 => n40764, A2 => n48312, B1 => n40770, B2 => 
                           n48322, ZN => n48101);
   U1752 : AOI22_X1 port map( A1 => n40765, A2 => n48316, B1 => n40766, B2 => 
                           n48264, ZN => n48100);
   U1753 : AOI22_X1 port map( A1 => n40767, A2 => n48313, B1 => n40769, B2 => 
                           n49077, ZN => n48099);
   U1754 : AOI22_X1 port map( A1 => n40768, A2 => n49079, B1 => n40763, B2 => 
                           n49076, ZN => n48098);
   U1755 : NAND4_X1 port map( A1 => n48101, A2 => n48100, A3 => n48099, A4 => 
                           n48098, ZN => n48107);
   U1756 : AOI22_X1 port map( A1 => n40565, A2 => n41000, B1 => n41347, B2 => 
                           n48322, ZN => n48105);
   U1757 : AOI22_X1 port map( A1 => n41300, A2 => n48315, B1 => n41262, B2 => 
                           n48264, ZN => n48104);
   U1758 : AOI22_X1 port map( A1 => n41122, A2 => n48312, B1 => n40991, B2 => 
                           n49076, ZN => n48103);
   U1759 : AOI22_X1 port map( A1 => n41025, A2 => n48313, B1 => n41304, B2 => 
                           n48285, ZN => n48102);
   U1760 : NAND4_X1 port map( A1 => n48105, A2 => n48104, A3 => n48103, A4 => 
                           n48102, ZN => n48106);
   U1761 : AOI22_X1 port map( A1 => n48108, A2 => n48107, B1 => n48329, B2 => 
                           n48106, ZN => n48109);
   U1762 : OAI21_X1 port map( B1 => n48133, B2 => n48110, A => n48109, ZN => 
                           OUT2(9));
   U1763 : AOI22_X1 port map( A1 => n41211, A2 => n40589, B1 => n40735, B2 => 
                           n48273, ZN => n48114);
   U1764 : AOI22_X1 port map( A1 => n40688, A2 => n49093, B1 => n40710, B2 => 
                           n49092, ZN => n48113);
   U1765 : AOI22_X1 port map( A1 => n41386, A2 => n40588, B1 => n41157, B2 => 
                           n49087, ZN => n48112);
   U1766 : AOI22_X1 port map( A1 => n47429, A2 => n41155, B1 => n40718, B2 => 
                           n49089, ZN => n48111);
   U1767 : NAND4_X1 port map( A1 => n48114, A2 => n48113, A3 => n48112, A4 => 
                           n48111, ZN => n48120);
   U1768 : AOI22_X1 port map( A1 => n40730, A2 => n40592, B1 => n41159, B2 => 
                           n49091, ZN => n48118);
   U1769 : AOI22_X1 port map( A1 => n40755, A2 => n49094, B1 => n41161, B2 => 
                           n49090, ZN => n48117);
   U1770 : AOI22_X1 port map( A1 => n47428, A2 => n41160, B1 => n41223, B2 => 
                           n49086, ZN => n48116);
   U1771 : AOI22_X1 port map( A1 => n41181, A2 => n40591, B1 => n41156, B2 => 
                           n49085, ZN => n48115);
   U1772 : NAND4_X1 port map( A1 => n48118, A2 => n48117, A3 => n48116, A4 => 
                           n48115, ZN => n48119);
   U1773 : NOR2_X1 port map( A1 => n48120, A2 => n48119, ZN => n48132);
   U1774 : AOI22_X1 port map( A1 => n40785, A2 => n49078, B1 => n40779, B2 => 
                           n48264, ZN => n48124);
   U1775 : AOI22_X1 port map( A1 => n40782, A2 => n48313, B1 => n40781, B2 => 
                           n49076, ZN => n48123);
   U1776 : AOI22_X1 port map( A1 => n40783, A2 => n48312, B1 => n40778, B2 => 
                           n49077, ZN => n48122);
   U1777 : AOI22_X1 port map( A1 => n40780, A2 => n40565, B1 => n40784, B2 => 
                           n48285, ZN => n48121);
   U1778 : NAND4_X1 port map( A1 => n48124, A2 => n48123, A3 => n48122, A4 => 
                           n48121, ZN => n48130);
   U1779 : AOI22_X1 port map( A1 => n41299, A2 => n48235, B1 => n41264, B2 => 
                           n48264, ZN => n48128);
   U1780 : AOI22_X1 port map( A1 => n40997, A2 => n41691, B1 => n41024, B2 => 
                           n49076, ZN => n48127);
   U1781 : AOI22_X1 port map( A1 => n41029, A2 => n48313, B1 => n41305, B2 => 
                           n48285, ZN => n48126);
   U1782 : AOI22_X1 port map( A1 => n41120, A2 => n48312, B1 => n41346, B2 => 
                           n48322, ZN => n48125);
   U1783 : NAND4_X1 port map( A1 => n48128, A2 => n48127, A3 => n48126, A4 => 
                           n48125, ZN => n48129);
   U1784 : AOI22_X1 port map( A1 => n48331, A2 => n48130, B1 => n48329, B2 => 
                           n48129, ZN => n48131);
   U1785 : OAI21_X1 port map( B1 => n48133, B2 => n48132, A => n48131, ZN => 
                           OUT2(8));
   U1786 : AOI22_X1 port map( A1 => n41683, A2 => n48274, B1 => n41682, B2 => 
                           n49087, ZN => n48137);
   U1787 : AOI22_X1 port map( A1 => n41664, A2 => n40588, B1 => n41655, B2 => 
                           n49086, ZN => n48136);
   U1788 : AOI22_X1 port map( A1 => n41034, A2 => n49088, B1 => n41039, B2 => 
                           n49089, ZN => n48135);
   U1789 : AOI22_X1 port map( A1 => n41684, A2 => n47429, B1 => n41036, B2 => 
                           n49092, ZN => n48134);
   U1790 : NAND4_X1 port map( A1 => n48137, A2 => n48136, A3 => n48135, A4 => 
                           n48134, ZN => n48143);
   U1791 : AOI22_X1 port map( A1 => n40589, A2 => n41667, B1 => n41037, B2 => 
                           n49094, ZN => n48141);
   U1792 : AOI22_X1 port map( A1 => n47428, A2 => n41678, B1 => n41035, B2 => 
                           n49093, ZN => n48140);
   U1793 : AOI22_X1 port map( A1 => n41038, A2 => n48305, B1 => n41679, B2 => 
                           n49091, ZN => n48139);
   U1794 : AOI22_X1 port map( A1 => n41669, A2 => n48299, B1 => n41674, B2 => 
                           n49085, ZN => n48138);
   U1795 : NAND4_X1 port map( A1 => n48141, A2 => n48140, A3 => n48139, A4 => 
                           n48138, ZN => n48142);
   U1796 : NOR2_X1 port map( A1 => n48143, A2 => n48142, ZN => n48155);
   U1797 : AOI22_X1 port map( A1 => n41466, A2 => n48312, B1 => n41456, B2 => 
                           n48322, ZN => n48147);
   U1798 : AOI22_X1 port map( A1 => n41465, A2 => n41691, B1 => n41463, B2 => 
                           n48285, ZN => n48146);
   U1799 : AOI22_X1 port map( A1 => n41469, A2 => n49076, B1 => n41455, B2 => 
                           n48264, ZN => n48145);
   U1800 : AOI22_X1 port map( A1 => n41458, A2 => n48313, B1 => n41457, B2 => 
                           n49077, ZN => n48144);
   U1801 : NAND4_X1 port map( A1 => n48147, A2 => n48146, A3 => n48145, A4 => 
                           n48144, ZN => n48153);
   U1802 : AOI22_X1 port map( A1 => n40565, A2 => n41552, B1 => n41578, B2 => 
                           n48192, ZN => n48151);
   U1803 : AOI22_X1 port map( A1 => n41550, A2 => n48313, B1 => n41547, B2 => 
                           n48314, ZN => n48150);
   U1804 : AOI22_X1 port map( A1 => n41616, A2 => n49077, B1 => n41591, B2 => 
                           n48323, ZN => n48149);
   U1805 : AOI22_X1 port map( A1 => n41588, A2 => n48322, B1 => n41681, B2 => 
                           n48264, ZN => n48148);
   U1806 : NAND4_X1 port map( A1 => n48151, A2 => n48150, A3 => n48149, A4 => 
                           n48148, ZN => n48152);
   U1807 : AOI22_X1 port map( A1 => n48331, A2 => n48153, B1 => n48329, B2 => 
                           n48152, ZN => n48154);
   U1808 : OAI21_X1 port map( B1 => n48334, B2 => n48155, A => n48154, ZN => 
                           OUT2(7));
   U1809 : AOI22_X1 port map( A1 => n41651, A2 => n40591, B1 => n40958, B2 => 
                           n48273, ZN => n48159);
   U1810 : AOI22_X1 port map( A1 => n41658, A2 => n40588, B1 => n40974, B2 => 
                           n49093, ZN => n48158);
   U1811 : AOI22_X1 port map( A1 => n40589, A2 => n41648, B1 => n40948, B2 => 
                           n49094, ZN => n48157);
   U1812 : AOI22_X1 port map( A1 => n41652, A2 => n47428, B1 => n40966, B2 => 
                           n49092, ZN => n48156);
   U1813 : NAND4_X1 port map( A1 => n48159, A2 => n48158, A3 => n48157, A4 => 
                           n48156, ZN => n48165);
   U1814 : AOI22_X1 port map( A1 => n47429, A2 => n41653, B1 => n48305, B2 => 
                           n40957, ZN => n48163);
   U1815 : AOI22_X1 port map( A1 => n41680, A2 => n49087, B1 => n41654, B2 => 
                           n49085, ZN => n48162);
   U1816 : AOI22_X1 port map( A1 => n41661, A2 => n49086, B1 => n41673, B2 => 
                           n49091, ZN => n48161);
   U1817 : AOI22_X1 port map( A1 => n41676, A2 => n48299, B1 => n40976, B2 => 
                           n49089, ZN => n48160);
   U1818 : NAND4_X1 port map( A1 => n48163, A2 => n48162, A3 => n48161, A4 => 
                           n48160, ZN => n48164);
   U1819 : NOR2_X1 port map( A1 => n48165, A2 => n48164, ZN => n48177);
   U1820 : AOI22_X1 port map( A1 => n40884, A2 => n49078, B1 => n40885, B2 => 
                           n49077, ZN => n48169);
   U1821 : AOI22_X1 port map( A1 => n40883, A2 => n48285, B1 => n40881, B2 => 
                           n48264, ZN => n48168);
   U1822 : AOI22_X1 port map( A1 => n40565, A2 => n40890, B1 => n40898, B2 => 
                           n48259, ZN => n48167);
   U1823 : AOI22_X1 port map( A1 => n40880, A2 => n48312, B1 => n40919, B2 => 
                           n49076, ZN => n48166);
   U1824 : NAND4_X1 port map( A1 => n48169, A2 => n48168, A3 => n48167, A4 => 
                           n48166, ZN => n48175);
   U1825 : AOI22_X1 port map( A1 => n41561, A2 => n48313, B1 => n41597, B2 => 
                           n48285, ZN => n48173);
   U1826 : AOI22_X1 port map( A1 => n41562, A2 => n41691, B1 => n41587, B2 => 
                           n48322, ZN => n48172);
   U1827 : AOI22_X1 port map( A1 => n41662, A2 => n48235, B1 => n41546, B2 => 
                           n49076, ZN => n48171);
   U1828 : AOI22_X1 port map( A1 => n41582, A2 => n48312, B1 => n41663, B2 => 
                           n48264, ZN => n48170);
   U1829 : NAND4_X1 port map( A1 => n48173, A2 => n48172, A3 => n48171, A4 => 
                           n48170, ZN => n48174);
   U1830 : AOI22_X1 port map( A1 => n48331, A2 => n48175, B1 => n48329, B2 => 
                           n48174, ZN => n48176);
   U1831 : OAI21_X1 port map( B1 => n48334, B2 => n48177, A => n48176, ZN => 
                           OUT2(6));
   U1832 : AOI22_X1 port map( A1 => n41644, A2 => n47428, B1 => n40965, B2 => 
                           n49092, ZN => n48181);
   U1833 : AOI22_X1 port map( A1 => n47429, A2 => n41631, B1 => n48205, B2 => 
                           n41634, ZN => n48180);
   U1834 : AOI22_X1 port map( A1 => n41656, A2 => n49086, B1 => n40979, B2 => 
                           n49089, ZN => n48179);
   U1835 : AOI22_X1 port map( A1 => n40589, A2 => n41629, B1 => n48305, B2 => 
                           n40970, ZN => n48178);
   U1836 : NAND4_X1 port map( A1 => n48181, A2 => n48180, A3 => n48179, A4 => 
                           n48178, ZN => n48187);
   U1837 : AOI22_X1 port map( A1 => n41650, A2 => n40591, B1 => n40950, B2 => 
                           n49093, ZN => n48185);
   U1838 : AOI22_X1 port map( A1 => n40968, A2 => n48273, B1 => n41633, B2 => 
                           n49085, ZN => n48184);
   U1839 : AOI22_X1 port map( A1 => n40951, A2 => n49094, B1 => n41641, B2 => 
                           n49087, ZN => n48183);
   U1840 : AOI22_X1 port map( A1 => n41645, A2 => n48299, B1 => n41642, B2 => 
                           n49091, ZN => n48182);
   U1841 : NAND4_X1 port map( A1 => n48185, A2 => n48184, A3 => n48183, A4 => 
                           n48182, ZN => n48186);
   U1842 : NOR2_X1 port map( A1 => n48187, A2 => n48186, ZN => n48200);
   U1843 : AOI22_X1 port map( A1 => n40876, A2 => n48323, B1 => n40877, B2 => 
                           n48264, ZN => n48191);
   U1844 : AOI22_X1 port map( A1 => n40878, A2 => n49078, B1 => n40894, B2 => 
                           n48314, ZN => n48190);
   U1845 : AOI22_X1 port map( A1 => n40897, A2 => n48313, B1 => n40879, B2 => 
                           n48192, ZN => n48189);
   U1846 : AOI22_X1 port map( A1 => n40889, A2 => n41691, B1 => n40886, B2 => 
                           n48315, ZN => n48188);
   U1847 : NAND4_X1 port map( A1 => n48191, A2 => n48190, A3 => n48189, A4 => 
                           n48188, ZN => n48198);
   U1848 : AOI22_X1 port map( A1 => n41564, A2 => n48314, B1 => n41637, B2 => 
                           n48264, ZN => n48196);
   U1849 : AOI22_X1 port map( A1 => n41592, A2 => n49078, B1 => n41639, B2 => 
                           n49077, ZN => n48195);
   U1850 : AOI22_X1 port map( A1 => n41565, A2 => n48316, B1 => n41593, B2 => 
                           n48285, ZN => n48194);
   U1851 : AOI22_X1 port map( A1 => n41551, A2 => n48313, B1 => n41581, B2 => 
                           n48192, ZN => n48193);
   U1852 : NAND4_X1 port map( A1 => n48196, A2 => n48195, A3 => n48194, A4 => 
                           n48193, ZN => n48197);
   U1853 : AOI22_X1 port map( A1 => n48331, A2 => n48198, B1 => n48329, B2 => 
                           n48197, ZN => n48199);
   U1854 : OAI21_X1 port map( B1 => n48334, B2 => n48200, A => n48199, ZN => 
                           OUT2(5));
   U1855 : AOI22_X1 port map( A1 => n41606, A2 => n48228, B1 => n40964, B2 => 
                           n49092, ZN => n48204);
   U1856 : AOI22_X1 port map( A1 => n48252, A2 => n41622, B1 => n41624, B2 => 
                           n49087, ZN => n48203);
   U1857 : AOI22_X1 port map( A1 => n41623, A2 => n48304, B1 => n40972, B2 => 
                           n49093, ZN => n48202);
   U1858 : AOI22_X1 port map( A1 => n41677, A2 => n49086, B1 => n41602, B2 => 
                           n49085, ZN => n48201);
   U1859 : NAND4_X1 port map( A1 => n48204, A2 => n48203, A3 => n48202, A4 => 
                           n48201, ZN => n48211);
   U1860 : AOI22_X1 port map( A1 => n40967, A2 => n49088, B1 => n41625, B2 => 
                           n49091, ZN => n48209);
   U1861 : AOI22_X1 port map( A1 => n48274, A2 => n41649, B1 => n40952, B2 => 
                           n49094, ZN => n48208);
   U1862 : AOI22_X1 port map( A1 => n41601, A2 => n48205, B1 => n40969, B2 => 
                           n49089, ZN => n48207);
   U1863 : AOI22_X1 port map( A1 => n40973, A2 => n48305, B1 => n41646, B2 => 
                           n48299, ZN => n48206);
   U1864 : NAND4_X1 port map( A1 => n48209, A2 => n48208, A3 => n48207, A4 => 
                           n48206, ZN => n48210);
   U1865 : NOR2_X1 port map( A1 => n48211, A2 => n48210, ZN => n48223);
   U1866 : AOI22_X1 port map( A1 => n40911, A2 => n40565, B1 => n40918, B2 => 
                           n48264, ZN => n48215);
   U1867 : AOI22_X1 port map( A1 => n40912, A2 => n48313, B1 => n40900, B2 => 
                           n48322, ZN => n48214);
   U1868 : AOI22_X1 port map( A1 => n40901, A2 => n49079, B1 => n40905, B2 => 
                           n48314, ZN => n48213);
   U1869 : AOI22_X1 port map( A1 => n40932, A2 => n48312, B1 => n40928, B2 => 
                           n48315, ZN => n48212);
   U1870 : NAND4_X1 port map( A1 => n48215, A2 => n48214, A3 => n48213, A4 => 
                           n48212, ZN => n48221);
   U1871 : AOI22_X1 port map( A1 => n41600, A2 => n48285, B1 => n41560, B2 => 
                           n48314, ZN => n48219);
   U1872 : AOI22_X1 port map( A1 => n41585, A2 => n48312, B1 => n41636, B2 => 
                           n48264, ZN => n48218);
   U1873 : AOI22_X1 port map( A1 => n41590, A2 => n48322, B1 => n41617, B2 => 
                           n48315, ZN => n48217);
   U1874 : AOI22_X1 port map( A1 => n40565, A2 => n41558, B1 => n41549, B2 => 
                           n48259, ZN => n48216);
   U1875 : NAND4_X1 port map( A1 => n48219, A2 => n48218, A3 => n48217, A4 => 
                           n48216, ZN => n48220);
   U1876 : AOI22_X1 port map( A1 => n48331, A2 => n48221, B1 => n48329, B2 => 
                           n48220, ZN => n48222);
   U1877 : OAI21_X1 port map( B1 => n48334, B2 => n48223, A => n48222, ZN => 
                           OUT2(4));
   U1878 : AOI22_X1 port map( A1 => n40953, A2 => n49094, B1 => n40981, B2 => 
                           n48273, ZN => n48227);
   U1879 : AOI22_X1 port map( A1 => n40947, A2 => n40592, B1 => n41675, B2 => 
                           n49086, ZN => n48226);
   U1880 : AOI22_X1 port map( A1 => n41643, A2 => n40591, B1 => n40975, B2 => 
                           n49089, ZN => n48225);
   U1881 : AOI22_X1 port map( A1 => n41621, A2 => n40589, B1 => n41647, B2 => 
                           n49090, ZN => n48224);
   U1882 : NAND4_X1 port map( A1 => n48227, A2 => n48226, A3 => n48225, A4 => 
                           n48224, ZN => n48234);
   U1883 : AOI22_X1 port map( A1 => n48252, A2 => n41620, B1 => n40978, B2 => 
                           n49093, ZN => n48232);
   U1884 : AOI22_X1 port map( A1 => n41613, A2 => n49087, B1 => n41614, B2 => 
                           n49091, ZN => n48231);
   U1885 : AOI22_X1 port map( A1 => n48228, A2 => n41611, B1 => n40588, B2 => 
                           n41608, ZN => n48230);
   U1886 : AOI22_X1 port map( A1 => n41610, A2 => n49085, B1 => n40962, B2 => 
                           n49092, ZN => n48229);
   U1887 : NAND4_X1 port map( A1 => n48232, A2 => n48231, A3 => n48230, A4 => 
                           n48229, ZN => n48233);
   U1888 : NOR2_X1 port map( A1 => n48234, A2 => n48233, ZN => n48247);
   U1889 : AOI22_X1 port map( A1 => n40895, A2 => n48312, B1 => n40908, B2 => 
                           n49078, ZN => n48239);
   U1890 : AOI22_X1 port map( A1 => n40899, A2 => n48313, B1 => n40910, B2 => 
                           n48264, ZN => n48238);
   U1891 : AOI22_X1 port map( A1 => n40896, A2 => n41691, B1 => n40916, B2 => 
                           n48314, ZN => n48237);
   U1892 : AOI22_X1 port map( A1 => n40907, A2 => n48235, B1 => n40909, B2 => 
                           n49079, ZN => n48236);
   U1893 : NAND4_X1 port map( A1 => n48239, A2 => n48238, A3 => n48237, A4 => 
                           n48236, ZN => n48245);
   U1894 : AOI22_X1 port map( A1 => n40565, A2 => n41555, B1 => n41544, B2 => 
                           n48313, ZN => n48243);
   U1895 : AOI22_X1 port map( A1 => n41598, A2 => n48322, B1 => n41548, B2 => 
                           n48314, ZN => n48242);
   U1896 : AOI22_X1 port map( A1 => n41577, A2 => n48312, B1 => n41626, B2 => 
                           n48315, ZN => n48241);
   U1897 : AOI22_X1 port map( A1 => n41596, A2 => n48285, B1 => n41635, B2 => 
                           n48264, ZN => n48240);
   U1898 : NAND4_X1 port map( A1 => n48243, A2 => n48242, A3 => n48241, A4 => 
                           n48240, ZN => n48244);
   U1899 : AOI22_X1 port map( A1 => n48331, A2 => n48245, B1 => n48329, B2 => 
                           n48244, ZN => n48246);
   U1900 : OAI21_X1 port map( B1 => n48334, B2 => n48247, A => n48246, ZN => 
                           OUT2(3));
   U1901 : AOI22_X1 port map( A1 => n40588, A2 => n41612, B1 => n40954, B2 => 
                           n49094, ZN => n48251);
   U1902 : AOI22_X1 port map( A1 => n40971, A2 => n49089, B1 => n41665, B2 => 
                           n49091, ZN => n48250);
   U1903 : AOI22_X1 port map( A1 => n41668, A2 => n40589, B1 => n41657, B2 => 
                           n49087, ZN => n48249);
   U1904 : AOI22_X1 port map( A1 => n40961, A2 => n40592, B1 => n40977, B2 => 
                           n49093, ZN => n48248);
   U1905 : NAND4_X1 port map( A1 => n48251, A2 => n48250, A3 => n48249, A4 => 
                           n48248, ZN => n48258);
   U1906 : AOI22_X1 port map( A1 => n41672, A2 => n48252, B1 => n40959, B2 => 
                           n49092, ZN => n48256);
   U1907 : AOI22_X1 port map( A1 => n41666, A2 => n40591, B1 => n41671, B2 => 
                           n49090, ZN => n48255);
   U1908 : AOI22_X1 port map( A1 => n47429, A2 => n41660, B1 => n41609, B2 => 
                           n49086, ZN => n48254);
   U1909 : AOI22_X1 port map( A1 => n40982, A2 => n48273, B1 => n41659, B2 => 
                           n49085, ZN => n48253);
   U1910 : NAND4_X1 port map( A1 => n48256, A2 => n48255, A3 => n48254, A4 => 
                           n48253, ZN => n48257);
   U1911 : NOR2_X1 port map( A1 => n48258, A2 => n48257, ZN => n48272);
   U1912 : AOI22_X1 port map( A1 => n40924, A2 => n48312, B1 => n40927, B2 => 
                           n49079, ZN => n48263);
   U1913 : AOI22_X1 port map( A1 => n40914, A2 => n41691, B1 => n40906, B2 => 
                           n48259, ZN => n48262);
   U1914 : AOI22_X1 port map( A1 => n40915, A2 => n49076, B1 => n40926, B2 => 
                           n48264, ZN => n48261);
   U1915 : AOI22_X1 port map( A1 => n40902, A2 => n48290, B1 => n40903, B2 => 
                           n48315, ZN => n48260);
   U1916 : NAND4_X1 port map( A1 => n48263, A2 => n48262, A3 => n48261, A4 => 
                           n48260, ZN => n48270);
   U1917 : AOI22_X1 port map( A1 => n41589, A2 => n48285, B1 => n41632, B2 => 
                           n48264, ZN => n48268);
   U1918 : AOI22_X1 port map( A1 => n41579, A2 => n48312, B1 => n41627, B2 => 
                           n48315, ZN => n48267);
   U1919 : AOI22_X1 port map( A1 => n48316, A2 => n41536, B1 => n41537, B2 => 
                           n48313, ZN => n48266);
   U1920 : AOI22_X1 port map( A1 => n41595, A2 => n48290, B1 => n41543, B2 => 
                           n48314, ZN => n48265);
   U1921 : NAND4_X1 port map( A1 => n48268, A2 => n48267, A3 => n48266, A4 => 
                           n48265, ZN => n48269);
   U1922 : AOI22_X1 port map( A1 => n48331, A2 => n48270, B1 => n48329, B2 => 
                           n48269, ZN => n48271);
   U1923 : OAI21_X1 port map( B1 => n48334, B2 => n48272, A => n48271, ZN => 
                           OUT2(2));
   U1924 : AOI22_X1 port map( A1 => n40956, A2 => n49094, B1 => n40963, B2 => 
                           n48273, ZN => n48278);
   U1925 : AOI22_X1 port map( A1 => n40960, A2 => n40592, B1 => n40980, B2 => 
                           n49089, ZN => n48277);
   U1926 : AOI22_X1 port map( A1 => n41604, A2 => n40588, B1 => n40955, B2 => 
                           n49093, ZN => n48276);
   U1927 : AOI22_X1 port map( A1 => n41638, A2 => n48274, B1 => n41603, B2 => 
                           n49086, ZN => n48275);
   U1928 : NAND4_X1 port map( A1 => n48278, A2 => n48277, A3 => n48276, A4 => 
                           n48275, ZN => n48284);
   U1929 : AOI22_X1 port map( A1 => n41670, A2 => n48299, B1 => n40949, B2 => 
                           n49092, ZN => n48282);
   U1930 : AOI22_X1 port map( A1 => n41619, A2 => n40589, B1 => n41605, B2 => 
                           n49085, ZN => n48281);
   U1931 : AOI22_X1 port map( A1 => n47429, A2 => n41607, B1 => n41640, B2 => 
                           n49087, ZN => n48280);
   U1932 : AOI22_X1 port map( A1 => n47428, A2 => n41618, B1 => n41615, B2 => 
                           n49091, ZN => n48279);
   U1933 : NAND4_X1 port map( A1 => n48282, A2 => n48281, A3 => n48280, A4 => 
                           n48279, ZN => n48283);
   U1934 : NOR2_X1 port map( A1 => n48284, A2 => n48283, ZN => n48298);
   U1935 : AOI22_X1 port map( A1 => n40921, A2 => n48312, B1 => n40913, B2 => 
                           n49078, ZN => n48289);
   U1936 : AOI22_X1 port map( A1 => n40936, A2 => n49076, B1 => n40920, B2 => 
                           n49082, ZN => n48288);
   U1937 : AOI22_X1 port map( A1 => n40923, A2 => n48313, B1 => n40917, B2 => 
                           n48285, ZN => n48287);
   U1938 : AOI22_X1 port map( A1 => n40922, A2 => n41691, B1 => n40930, B2 => 
                           n48315, ZN => n48286);
   U1939 : NAND4_X1 port map( A1 => n48289, A2 => n48288, A3 => n48287, A4 => 
                           n48286, ZN => n48296);
   U1940 : AOI22_X1 port map( A1 => n41628, A2 => n49077, B1 => n41599, B2 => 
                           n49079, ZN => n48294);
   U1941 : AOI22_X1 port map( A1 => n48316, A2 => n41563, B1 => n41594, B2 => 
                           n48290, ZN => n48293);
   U1942 : AOI22_X1 port map( A1 => n41586, A2 => n48312, B1 => n41553, B2 => 
                           n48314, ZN => n48292);
   U1943 : AOI22_X1 port map( A1 => n41559, A2 => n48313, B1 => n41630, B2 => 
                           n49082, ZN => n48291);
   U1944 : NAND4_X1 port map( A1 => n48294, A2 => n48293, A3 => n48292, A4 => 
                           n48291, ZN => n48295);
   U1945 : AOI22_X1 port map( A1 => n48331, A2 => n48296, B1 => n48329, B2 => 
                           n48295, ZN => n48297);
   U1946 : OAI21_X1 port map( B1 => n48334, B2 => n48298, A => n48297, ZN => 
                           OUT2(1));
   U1947 : AOI22_X1 port map( A1 => n41570, A2 => n40591, B1 => n41566, B2 => 
                           n49085, ZN => n48303);
   U1948 : AOI22_X1 port map( A1 => n47429, A2 => n41501, B1 => n41571, B2 => 
                           n49086, ZN => n48302);
   U1949 : AOI22_X1 port map( A1 => n40875, A2 => n49088, B1 => n41572, B2 => 
                           n49087, ZN => n48301);
   U1950 : AOI22_X1 port map( A1 => n41567, A2 => n48299, B1 => n40873, B2 => 
                           n49089, ZN => n48300);
   U1951 : NAND4_X1 port map( A1 => n48303, A2 => n48302, A3 => n48301, A4 => 
                           n48300, ZN => n48311);
   U1952 : AOI22_X1 port map( A1 => n47428, A2 => n41575, B1 => n48304, B2 => 
                           n41576, ZN => n48309);
   U1953 : AOI22_X1 port map( A1 => n40872, A2 => n48305, B1 => n41574, B2 => 
                           n49091, ZN => n48308);
   U1954 : AOI22_X1 port map( A1 => n40870, A2 => n49093, B1 => n40871, B2 => 
                           n49092, ZN => n48307);
   U1955 : AOI22_X1 port map( A1 => n40588, A2 => n41487, B1 => n40874, B2 => 
                           n49094, ZN => n48306);
   U1956 : NAND4_X1 port map( A1 => n48309, A2 => n48308, A3 => n48307, A4 => 
                           n48306, ZN => n48310);
   U1957 : NOR2_X1 port map( A1 => n48311, A2 => n48310, ZN => n48333);
   U1958 : AOI22_X1 port map( A1 => n40944, A2 => n48312, B1 => n40945, B2 => 
                           n49082, ZN => n48320);
   U1959 : AOI22_X1 port map( A1 => n40943, A2 => n48313, B1 => n41685, B2 => 
                           n48323, ZN => n48319);
   U1960 : AOI22_X1 port map( A1 => n40941, A2 => n48322, B1 => n40942, B2 => 
                           n48314, ZN => n48318);
   U1961 : AOI22_X1 port map( A1 => n48316, A2 => n40940, B1 => n40946, B2 => 
                           n48315, ZN => n48317);
   U1962 : NAND4_X1 port map( A1 => n48320, A2 => n48319, A3 => n48318, A4 => 
                           n48317, ZN => n48330);
   U1963 : AOI22_X1 port map( A1 => n41440, A2 => n49081, B1 => n41442, B2 => 
                           n48321, ZN => n48327);
   U1964 : AOI22_X1 port map( A1 => n41454, A2 => n49080, B1 => n41492, B2 => 
                           n49077, ZN => n48326);
   U1965 : AOI22_X1 port map( A1 => n40565, A2 => n41441, B1 => n41573, B2 => 
                           n48322, ZN => n48325);
   U1966 : AOI22_X1 port map( A1 => n41568, A2 => n48323, B1 => n41569, B2 => 
                           n49082, ZN => n48324);
   U1967 : NAND4_X1 port map( A1 => n48327, A2 => n48326, A3 => n48325, A4 => 
                           n48324, ZN => n48328);
   U1968 : AOI22_X1 port map( A1 => n48331, A2 => n48330, B1 => n48329, B2 => 
                           n48328, ZN => n48332);
   U1969 : OAI21_X1 port map( B1 => n48334, B2 => n48333, A => n48332, ZN => 
                           OUT2(0));
   U1970 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n48338)
                           ;
   U1971 : NOR2_X1 port map( A1 => n1529, A2 => n48338, ZN => n30068);
   U1972 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n48335);
   U1973 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => n48335, ZN => n47499);
   U1974 : INV_X1 port map( A => ADD_RD1(3), ZN => n48336);
   U1975 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n48336, ZN => n48337);
   U1976 : NOR2_X1 port map( A1 => n48337, A2 => n47499, ZN => n30067);
   U1977 : NOR2_X1 port map( A1 => n1529, A2 => n48337, ZN => n30066);
   U1978 : NOR2_X1 port map( A1 => n48338, A2 => n1532, ZN => n30065);
   U1979 : NOR2_X1 port map( A1 => n48337, A2 => n1530, ZN => n30064);
   U1980 : NOR2_X1 port map( A1 => n48337, A2 => n1531, ZN => n30063);
   U1981 : NOR2_X1 port map( A1 => n48337, A2 => n1528, ZN => n30062);
   U1982 : NOR2_X1 port map( A1 => n48337, A2 => n1532, ZN => n30061);
   U1983 : NOR2_X1 port map( A1 => n48338, A2 => n47499, ZN => n30060);
   U1984 : NOR2_X1 port map( A1 => n48338, A2 => n1531, ZN => n30059);
   U1985 : NOR2_X1 port map( A1 => n48337, A2 => n47501, ZN => n30058);
   U1986 : NOR2_X1 port map( A1 => n48338, A2 => n47501, ZN => n30057);
   U1987 : NOR2_X1 port map( A1 => n48337, A2 => n1527, ZN => n30056);
   U1988 : NOR2_X1 port map( A1 => n48338, A2 => n1528, ZN => n30055);
   U1989 : NOR2_X1 port map( A1 => n48338, A2 => n1530, ZN => n30054);
   U1990 : NOR2_X1 port map( A1 => n48338, A2 => n1527, ZN => n30053);
   U1991 : CLKBUF_X1 port map( A => n40581, Z => n49015);
   U1992 : AOI22_X1 port map( A1 => n41331, A2 => n49015, B1 => n41326, B2 => 
                           n40587, ZN => n48342);
   U1993 : CLKBUF_X1 port map( A => n40582, Z => n49014);
   U1994 : AOI22_X1 port map( A1 => n41327, A2 => n49014, B1 => n41393, B2 => 
                           n40580, ZN => n48341);
   U1995 : AOI22_X1 port map( A1 => n41332, A2 => n49096, B1 => n41329, B2 => 
                           n40583, ZN => n48340);
   U1996 : CLKBUF_X1 port map( A => n40576, Z => n49022);
   U1997 : AOI22_X1 port map( A1 => n40789, A2 => n49022, B1 => n40831, B2 => 
                           n40584, ZN => n48339);
   U1998 : NAND4_X1 port map( A1 => n48342, A2 => n48341, A3 => n48340, A4 => 
                           n48339, ZN => n48348);
   U1999 : CLKBUF_X1 port map( A => n40585, Z => n49023);
   U2000 : AOI22_X1 port map( A1 => n41333, A2 => n49023, B1 => n40803, B2 => 
                           n49095, ZN => n48346);
   U2001 : CLKBUF_X1 port map( A => n40574, Z => n49013);
   U2002 : AOI22_X1 port map( A1 => n41330, A2 => n40586, B1 => n40808, B2 => 
                           n49013, ZN => n48345);
   U2003 : CLKBUF_X1 port map( A => n47431, Z => n48962);
   U2004 : CLKBUF_X1 port map( A => n40577, Z => n48992);
   U2005 : AOI22_X1 port map( A1 => n41325, A2 => n48962, B1 => n41328, B2 => 
                           n48992, ZN => n48344);
   U2006 : AOI22_X1 port map( A1 => n40812, A2 => n49097, B1 => n40823, B2 => 
                           n47430, ZN => n48343);
   U2007 : NAND4_X1 port map( A1 => n48346, A2 => n48345, A3 => n48344, A4 => 
                           n48343, ZN => n48347);
   U2008 : NOR2_X1 port map( A1 => n48348, A2 => n48347, ZN => n48360);
   U2009 : NOR3_X1 port map( A1 => n40656, A2 => n42756, A3 => n49012, ZN => 
                           n48882);
   U2010 : CLKBUF_X1 port map( A => n48882, Z => n48869);
   U2011 : CLKBUF_X1 port map( A => n40655, Z => n48883);
   U2012 : AOI22_X1 port map( A1 => n40663, A2 => n48883, B1 => n40671, B2 => 
                           n40649, ZN => n48352);
   U2013 : INV_X1 port map( A => n47446, ZN => n49063);
   U2014 : AOI22_X1 port map( A1 => n40670, A2 => n41686, B1 => n40672, B2 => 
                           n49063, ZN => n48351);
   U2015 : CLKBUF_X1 port map( A => n40648, Z => n49055);
   U2016 : AOI22_X1 port map( A1 => n40664, A2 => n49083, B1 => n40673, B2 => 
                           n49055, ZN => n48350);
   U2017 : AOI22_X1 port map( A1 => n40676, A2 => n41690, B1 => n40665, B2 => 
                           n40654, ZN => n48349);
   U2018 : NAND4_X1 port map( A1 => n48352, A2 => n48351, A3 => n48350, A4 => 
                           n48349, ZN => n48358);
   U2019 : NOR3_X1 port map( A1 => n42756, A2 => n42722, A3 => n49012, ZN => 
                           n48578);
   U2020 : INV_X1 port map( A => n47447, ZN => n49062);
   U2021 : CLKBUF_X1 port map( A => n49062, Z => n48792);
   U2022 : AOI22_X1 port map( A1 => n41322, A2 => n48792, B1 => n41320, B2 => 
                           n49063, ZN => n48356);
   U2023 : AOI22_X1 port map( A1 => n41321, A2 => n48883, B1 => n41338, B2 => 
                           n41688, ZN => n48355);
   U2024 : CLKBUF_X1 port map( A => n40568, Z => n48979);
   U2025 : AOI22_X1 port map( A1 => n41027, A2 => n48979, B1 => n41123, B2 => 
                           n41689, ZN => n48354);
   U2026 : AOI22_X1 port map( A1 => n41008, A2 => n40649, B1 => n40989, B2 => 
                           n40571, ZN => n48353);
   U2027 : NAND4_X1 port map( A1 => n48356, A2 => n48355, A3 => n48354, A4 => 
                           n48353, ZN => n48357);
   U2028 : AOI22_X1 port map( A1 => n48869, A2 => n48358, B1 => n48578, B2 => 
                           n48357, ZN => n48359);
   U2029 : OAI21_X1 port map( B1 => n49012, B2 => n48360, A => n48359, ZN => 
                           OUT1(31));
   U2030 : CLKBUF_X1 port map( A => n49097, Z => n49017);
   U2031 : AOI22_X1 port map( A1 => n41394, A2 => n40580, B1 => n41062, B2 => 
                           n49017, ZN => n48364);
   U2032 : CLKBUF_X1 port map( A => n49095, Z => n48785);
   U2033 : AOI22_X1 port map( A1 => n41281, A2 => n49096, B1 => n41091, B2 => 
                           n48785, ZN => n48363);
   U2034 : AOI22_X1 port map( A1 => n41279, A2 => n40583, B1 => n41496, B2 => 
                           n40587, ZN => n48362);
   U2035 : CLKBUF_X1 port map( A => n40584, Z => n48968);
   U2036 : AOI22_X1 port map( A1 => n41276, A2 => n40582, B1 => n41493, B2 => 
                           n48968, ZN => n48361);
   U2037 : NAND4_X1 port map( A1 => n48364, A2 => n48363, A3 => n48362, A4 => 
                           n48361, ZN => n48370);
   U2038 : AOI22_X1 port map( A1 => n41278, A2 => n48992, B1 => n41283, B2 => 
                           n47431, ZN => n48368);
   U2039 : AOI22_X1 port map( A1 => n41098, A2 => n40576, B1 => n41103, B2 => 
                           n47430, ZN => n48367);
   U2040 : AOI22_X1 port map( A1 => n41284, A2 => n40585, B1 => n41075, B2 => 
                           n40574, ZN => n48366);
   U2041 : CLKBUF_X1 port map( A => n40586, Z => n48967);
   U2042 : AOI22_X1 port map( A1 => n41280, A2 => n40581, B1 => n41508, B2 => 
                           n48967, ZN => n48365);
   U2043 : NAND4_X1 port map( A1 => n48368, A2 => n48367, A3 => n48366, A4 => 
                           n48365, ZN => n48369);
   U2044 : NOR2_X1 port map( A1 => n48370, A2 => n48369, ZN => n48382);
   U2045 : AOI22_X1 port map( A1 => n41498, A2 => n48792, B1 => n41497, B2 => 
                           n40648, ZN => n48374);
   U2046 : AOI22_X1 port map( A1 => n41503, A2 => n40654, B1 => n41523, B2 => 
                           n41686, ZN => n48373);
   U2047 : AOI22_X1 port map( A1 => n41500, A2 => n49084, B1 => n41087, B2 => 
                           n41687, ZN => n48372);
   U2048 : AOI22_X1 port map( A1 => n41066, A2 => n40571, B1 => n41499, B2 => 
                           n40655, ZN => n48371);
   U2049 : NAND4_X1 port map( A1 => n48374, A2 => n48373, A3 => n48372, A4 => 
                           n48371, ZN => n48380);
   U2050 : CLKBUF_X1 port map( A => n48578, Z => n49070);
   U2051 : CLKBUF_X1 port map( A => n40649, Z => n49057);
   U2052 : AOI22_X1 port map( A1 => n41047, A2 => n49057, B1 => n41275, B2 => 
                           n49083, ZN => n48378);
   U2053 : CLKBUF_X1 port map( A => n40654, Z => n49056);
   U2054 : AOI22_X1 port map( A1 => n41040, A2 => n40571, B1 => n41337, B2 => 
                           n49056, ZN => n48377);
   U2055 : AOI22_X1 port map( A1 => n41104, A2 => n40648, B1 => n41054, B2 => 
                           n48979, ZN => n48376);
   U2056 : AOI22_X1 port map( A1 => n41309, A2 => n49084, B1 => n41513, B2 => 
                           n40655, ZN => n48375);
   U2057 : NAND4_X1 port map( A1 => n48378, A2 => n48377, A3 => n48376, A4 => 
                           n48375, ZN => n48379);
   U2058 : AOI22_X1 port map( A1 => n48869, A2 => n48380, B1 => n49070, B2 => 
                           n48379, ZN => n48381);
   U2059 : OAI21_X1 port map( B1 => n49012, B2 => n48382, A => n48381, ZN => 
                           OUT1(30));
   U2060 : AOI22_X1 port map( A1 => n41302, A2 => n40587, B1 => n40746, B2 => 
                           n49022, ZN => n48386);
   U2061 : AOI22_X1 port map( A1 => n40719, A2 => n49095, B1 => n40814, B2 => 
                           n40584, ZN => n48385);
   U2062 : AOI22_X1 port map( A1 => n41292, A2 => n40581, B1 => n41288, B2 => 
                           n49014, ZN => n48384);
   U2063 : AOI22_X1 port map( A1 => n40759, A2 => n49097, B1 => n41293, B2 => 
                           n49096, ZN => n48383);
   U2064 : NAND4_X1 port map( A1 => n48386, A2 => n48385, A3 => n48384, A4 => 
                           n48383, ZN => n48392);
   U2065 : AOI22_X1 port map( A1 => n41395, A2 => n40580, B1 => n41291, B2 => 
                           n40586, ZN => n48390);
   U2066 : AOI22_X1 port map( A1 => n41301, A2 => n48962, B1 => n41289, B2 => 
                           n48992, ZN => n48389);
   U2067 : AOI22_X1 port map( A1 => n41290, A2 => n40583, B1 => n41295, B2 => 
                           n49023, ZN => n48388);
   U2068 : AOI22_X1 port map( A1 => n40682, A2 => n40574, B1 => n40693, B2 => 
                           n47430, ZN => n48387);
   U2069 : NAND4_X1 port map( A1 => n48390, A2 => n48389, A3 => n48388, A4 => 
                           n48387, ZN => n48391);
   U2070 : NOR2_X1 port map( A1 => n48392, A2 => n48391, ZN => n48404);
   U2071 : AOI22_X1 port map( A1 => n40668, A2 => n40649, B1 => n40669, B2 => 
                           n41690, ZN => n48396);
   U2072 : AOI22_X1 port map( A1 => n40788, A2 => n48883, B1 => n40786, B2 => 
                           n41688, ZN => n48395);
   U2073 : AOI22_X1 port map( A1 => n40787, A2 => n49084, B1 => n40790, B2 => 
                           n49083, ZN => n48394);
   U2074 : AOI22_X1 port map( A1 => n40791, A2 => n49055, B1 => n40792, B2 => 
                           n41686, ZN => n48393);
   U2075 : NAND4_X1 port map( A1 => n48396, A2 => n48395, A3 => n48394, A4 => 
                           n48393, ZN => n48402);
   U2076 : AOI22_X1 port map( A1 => n41310, A2 => n49084, B1 => n41006, B2 => 
                           n49057, ZN => n48400);
   U2077 : AOI22_X1 port map( A1 => n41296, A2 => n40655, B1 => n40996, B2 => 
                           n40568, ZN => n48399);
   U2078 : AOI22_X1 port map( A1 => n41336, A2 => n49056, B1 => n41107, B2 => 
                           n41689, ZN => n48398);
   U2079 : CLKBUF_X1 port map( A => n40571, Z => n49064);
   U2080 : AOI22_X1 port map( A1 => n40995, A2 => n49064, B1 => n41421, B2 => 
                           n49062, ZN => n48397);
   U2081 : NAND4_X1 port map( A1 => n48400, A2 => n48399, A3 => n48398, A4 => 
                           n48397, ZN => n48401);
   U2082 : AOI22_X1 port map( A1 => n48869, A2 => n48402, B1 => n49070, B2 => 
                           n48401, ZN => n48403);
   U2083 : OAI21_X1 port map( B1 => n49012, B2 => n48404, A => n48403, ZN => 
                           OUT1(29));
   U2084 : AOI22_X1 port map( A1 => n41263, A2 => n47431, B1 => n41519, B2 => 
                           n40587, ZN => n48408);
   U2085 : AOI22_X1 port map( A1 => n41094, A2 => n47430, B1 => n41516, B2 => 
                           n40586, ZN => n48407);
   U2086 : AOI22_X1 port map( A1 => n41252, A2 => n40577, B1 => n41518, B2 => 
                           n40584, ZN => n48406);
   U2087 : AOI22_X1 port map( A1 => n41076, A2 => n40574, B1 => n41265, B2 => 
                           n40582, ZN => n48405);
   U2088 : NAND4_X1 port map( A1 => n48408, A2 => n48407, A3 => n48406, A4 => 
                           n48405, ZN => n48414);
   U2089 : AOI22_X1 port map( A1 => n41083, A2 => n49022, B1 => n41253, B2 => 
                           n40583, ZN => n48412);
   U2090 : AOI22_X1 port map( A1 => n41259, A2 => n49096, B1 => n41063, B2 => 
                           n49017, ZN => n48411);
   U2091 : AOI22_X1 port map( A1 => n41258, A2 => n40581, B1 => n41084, B2 => 
                           n48785, ZN => n48410);
   U2092 : AOI22_X1 port map( A1 => n41282, A2 => n40585, B1 => n41402, B2 => 
                           n40580, ZN => n48409);
   U2093 : NAND4_X1 port map( A1 => n48412, A2 => n48411, A3 => n48410, A4 => 
                           n48409, ZN => n48413);
   U2094 : NOR2_X1 port map( A1 => n48414, A2 => n48413, ZN => n48426);
   U2095 : AOI22_X1 port map( A1 => n41506, A2 => n49062, B1 => n41505, B2 => 
                           n41692, ZN => n48418);
   U2096 : CLKBUF_X1 port map( A => n49063, Z => n49003);
   U2097 : AOI22_X1 port map( A1 => n41512, A2 => n41686, B1 => n41504, B2 => 
                           n49003, ZN => n48417);
   U2098 : AOI22_X1 port map( A1 => n41088, A2 => n49057, B1 => n41502, B2 => 
                           n41688, ZN => n48416);
   U2099 : AOI22_X1 port map( A1 => n41511, A2 => n49055, B1 => n41067, B2 => 
                           n40571, ZN => n48415);
   U2100 : NAND4_X1 port map( A1 => n48418, A2 => n48417, A3 => n48416, A4 => 
                           n48415, ZN => n48424);
   U2101 : AOI22_X1 port map( A1 => n41335, A2 => n49056, B1 => n41261, B2 => 
                           n49062, ZN => n48422);
   U2102 : AOI22_X1 port map( A1 => n41048, A2 => n41687, B1 => n41517, B2 => 
                           n40655, ZN => n48421);
   U2103 : AOI22_X1 port map( A1 => n41311, A2 => n49084, B1 => n41070, B2 => 
                           n40571, ZN => n48420);
   U2104 : AOI22_X1 port map( A1 => n41055, A2 => n48979, B1 => n41119, B2 => 
                           n40648, ZN => n48419);
   U2105 : NAND4_X1 port map( A1 => n48422, A2 => n48421, A3 => n48420, A4 => 
                           n48419, ZN => n48423);
   U2106 : AOI22_X1 port map( A1 => n48869, A2 => n48424, B1 => n49070, B2 => 
                           n48423, ZN => n48425);
   U2107 : OAI21_X1 port map( B1 => n49012, B2 => n48426, A => n48425, ZN => 
                           OUT1(28));
   U2108 : AOI22_X1 port map( A1 => n41273, A2 => n40577, B1 => n41079, B2 => 
                           n40576, ZN => n48430);
   U2109 : CLKBUF_X1 port map( A => n40587, Z => n49024);
   U2110 : AOI22_X1 port map( A1 => n41064, A2 => n49097, B1 => n41514, B2 => 
                           n49024, ZN => n48429);
   U2111 : CLKBUF_X1 port map( A => n40580, Z => n49026);
   U2112 : AOI22_X1 port map( A1 => n41271, A2 => n47431, B1 => n41403, B2 => 
                           n49026, ZN => n48428);
   U2113 : AOI22_X1 port map( A1 => n41269, A2 => n40585, B1 => n41515, B2 => 
                           n40584, ZN => n48427);
   U2114 : NAND4_X1 port map( A1 => n48430, A2 => n48429, A3 => n48428, A4 => 
                           n48427, ZN => n48436);
   U2115 : CLKBUF_X1 port map( A => n49096, Z => n48758);
   U2116 : AOI22_X1 port map( A1 => n41266, A2 => n40583, B1 => n41268, B2 => 
                           n48758, ZN => n48434);
   U2117 : CLKBUF_X1 port map( A => n47430, Z => n49016);
   U2118 : AOI22_X1 port map( A1 => n41096, A2 => n49095, B1 => n41085, B2 => 
                           n49016, ZN => n48433);
   U2119 : AOI22_X1 port map( A1 => n41509, A2 => n48967, B1 => n41272, B2 => 
                           n49014, ZN => n48432);
   U2120 : AOI22_X1 port map( A1 => n41077, A2 => n40574, B1 => n41267, B2 => 
                           n49015, ZN => n48431);
   U2121 : NAND4_X1 port map( A1 => n48434, A2 => n48433, A3 => n48432, A4 => 
                           n48431, ZN => n48435);
   U2122 : NOR2_X1 port map( A1 => n48436, A2 => n48435, ZN => n48448);
   U2123 : AOI22_X1 port map( A1 => n41525, A2 => n49062, B1 => n41527, B2 => 
                           n41686, ZN => n48440);
   U2124 : AOI22_X1 port map( A1 => n41071, A2 => n49057, B1 => n41520, B2 => 
                           n41688, ZN => n48439);
   U2125 : AOI22_X1 port map( A1 => n41522, A2 => n49084, B1 => n41535, B2 => 
                           n49055, ZN => n48438);
   U2126 : AOI22_X1 port map( A1 => n41524, A2 => n40655, B1 => n41068, B2 => 
                           n49064, ZN => n48437);
   U2127 : NAND4_X1 port map( A1 => n48440, A2 => n48439, A3 => n48438, A4 => 
                           n48437, ZN => n48446);
   U2128 : AOI22_X1 port map( A1 => n41056, A2 => n48979, B1 => n41521, B2 => 
                           n48883, ZN => n48444);
   U2129 : AOI22_X1 port map( A1 => n41041, A2 => n41690, B1 => n41312, B2 => 
                           n49003, ZN => n48443);
   U2130 : AOI22_X1 port map( A1 => n41270, A2 => n48792, B1 => n41334, B2 => 
                           n40654, ZN => n48442);
   U2131 : AOI22_X1 port map( A1 => n41049, A2 => n49057, B1 => n41105, B2 => 
                           n49055, ZN => n48441);
   U2132 : NAND4_X1 port map( A1 => n48444, A2 => n48443, A3 => n48442, A4 => 
                           n48441, ZN => n48445);
   U2133 : AOI22_X1 port map( A1 => n48869, A2 => n48446, B1 => n48578, B2 => 
                           n48445, ZN => n48447);
   U2134 : OAI21_X1 port map( B1 => n49012, B2 => n48448, A => n48447, ZN => 
                           OUT1(27));
   U2135 : AOI22_X1 port map( A1 => n41238, A2 => n40586, B1 => n41235, B2 => 
                           n40582, ZN => n48452);
   U2136 : AOI22_X1 port map( A1 => n41236, A2 => n40577, B1 => n40681, B2 => 
                           n40574, ZN => n48451);
   U2137 : AOI22_X1 port map( A1 => n40687, A2 => n47430, B1 => n41241, B2 => 
                           n48758, ZN => n48450);
   U2138 : AOI22_X1 port map( A1 => n41233, A2 => n47431, B1 => n40720, B2 => 
                           n48785, ZN => n48449);
   U2139 : NAND4_X1 port map( A1 => n48452, A2 => n48451, A3 => n48450, A4 => 
                           n48449, ZN => n48458);
   U2140 : AOI22_X1 port map( A1 => n40813, A2 => n40584, B1 => n41249, B2 => 
                           n40585, ZN => n48456);
   U2141 : AOI22_X1 port map( A1 => n40758, A2 => n40576, B1 => n41404, B2 => 
                           n49026, ZN => n48455);
   U2142 : AOI22_X1 port map( A1 => n41239, A2 => n49015, B1 => n41234, B2 => 
                           n40587, ZN => n48454);
   U2143 : AOI22_X1 port map( A1 => n40739, A2 => n49097, B1 => n41237, B2 => 
                           n40583, ZN => n48453);
   U2144 : NAND4_X1 port map( A1 => n48456, A2 => n48455, A3 => n48454, A4 => 
                           n48453, ZN => n48457);
   U2145 : NOR2_X1 port map( A1 => n48458, A2 => n48457, ZN => n48470);
   U2146 : AOI22_X1 port map( A1 => n40794, A2 => n40654, B1 => n40805, B2 => 
                           n49055, ZN => n48462);
   U2147 : AOI22_X1 port map( A1 => n40806, A2 => n49062, B1 => n40807, B2 => 
                           n48883, ZN => n48461);
   U2148 : AOI22_X1 port map( A1 => n40667, A2 => n40571, B1 => n40675, B2 => 
                           n40649, ZN => n48460);
   U2149 : AOI22_X1 port map( A1 => n40804, A2 => n40568, B1 => n40793, B2 => 
                           n49003, ZN => n48459);
   U2150 : NAND4_X1 port map( A1 => n48462, A2 => n48461, A3 => n48460, A4 => 
                           n48459, ZN => n48468);
   U2151 : AOI22_X1 port map( A1 => n41230, A2 => n49062, B1 => n41324, B2 => 
                           n40654, ZN => n48466);
   U2152 : AOI22_X1 port map( A1 => n40998, A2 => n49064, B1 => n41021, B2 => 
                           n40649, ZN => n48465);
   U2153 : AOI22_X1 port map( A1 => n41115, A2 => n41689, B1 => n41313, B2 => 
                           n49003, ZN => n48464);
   U2154 : AOI22_X1 port map( A1 => n41020, A2 => n41686, B1 => n41274, B2 => 
                           n41692, ZN => n48463);
   U2155 : NAND4_X1 port map( A1 => n48466, A2 => n48465, A3 => n48464, A4 => 
                           n48463, ZN => n48467);
   U2156 : AOI22_X1 port map( A1 => n48869, A2 => n48468, B1 => n49070, B2 => 
                           n48467, ZN => n48469);
   U2157 : OAI21_X1 port map( B1 => n49012, B2 => n48470, A => n48469, ZN => 
                           OUT1(26));
   U2158 : AOI22_X1 port map( A1 => n41350, A2 => n49023, B1 => n41220, B2 => 
                           n49014, ZN => n48474);
   U2159 : AOI22_X1 port map( A1 => n41351, A2 => n40581, B1 => n41533, B2 => 
                           n40586, ZN => n48473);
   U2160 : CLKBUF_X1 port map( A => n40583, Z => n49025);
   U2161 : AOI22_X1 port map( A1 => n41097, A2 => n49095, B1 => n41222, B2 => 
                           n49025, ZN => n48472);
   U2162 : AOI22_X1 port map( A1 => n41078, A2 => n49013, B1 => n41065, B2 => 
                           n49017, ZN => n48471);
   U2163 : NAND4_X1 port map( A1 => n48474, A2 => n48473, A3 => n48472, A4 => 
                           n48471, ZN => n48480);
   U2164 : AOI22_X1 port map( A1 => n41221, A2 => n48992, B1 => n41219, B2 => 
                           n47431, ZN => n48478);
   U2165 : AOI22_X1 port map( A1 => n41102, A2 => n49016, B1 => n41405, B2 => 
                           n49026, ZN => n48477);
   U2166 : AOI22_X1 port map( A1 => n41349, A2 => n49096, B1 => n41531, B2 => 
                           n48968, ZN => n48476);
   U2167 : AOI22_X1 port map( A1 => n41080, A2 => n49022, B1 => n41532, B2 => 
                           n49024, ZN => n48475);
   U2168 : NAND4_X1 port map( A1 => n48478, A2 => n48477, A3 => n48476, A4 => 
                           n48475, ZN => n48479);
   U2169 : NOR2_X1 port map( A1 => n48480, A2 => n48479, ZN => n48492);
   U2170 : AOI22_X1 port map( A1 => n41479, A2 => n48979, B1 => n41069, B2 => 
                           n40571, ZN => n48484);
   U2171 : AOI22_X1 port map( A1 => n41090, A2 => n40649, B1 => n41534, B2 => 
                           n49063, ZN => n48483);
   U2172 : AOI22_X1 port map( A1 => n41526, A2 => n48792, B1 => n41489, B2 => 
                           n41689, ZN => n48482);
   U2173 : AOI22_X1 port map( A1 => n41528, A2 => n40655, B1 => n41529, B2 => 
                           n41688, ZN => n48481);
   U2174 : NAND4_X1 port map( A1 => n48484, A2 => n48483, A3 => n48482, A4 => 
                           n48481, ZN => n48490);
   U2175 : AOI22_X1 port map( A1 => n41510, A2 => n40655, B1 => n41057, B2 => 
                           n41686, ZN => n48488);
   U2176 : AOI22_X1 port map( A1 => n41108, A2 => n40648, B1 => n41277, B2 => 
                           n48792, ZN => n48487);
   U2177 : AOI22_X1 port map( A1 => n41424, A2 => n49063, B1 => n41372, B2 => 
                           n49056, ZN => n48486);
   U2178 : AOI22_X1 port map( A1 => n41050, A2 => n41687, B1 => n41043, B2 => 
                           n41690, ZN => n48485);
   U2179 : NAND4_X1 port map( A1 => n48488, A2 => n48487, A3 => n48486, A4 => 
                           n48485, ZN => n48489);
   U2180 : AOI22_X1 port map( A1 => n48869, A2 => n48490, B1 => n48578, B2 => 
                           n48489, ZN => n48491);
   U2181 : OAI21_X1 port map( B1 => n49012, B2 => n48492, A => n48491, ZN => 
                           OUT1(25));
   U2182 : AOI22_X1 port map( A1 => n41398, A2 => n48992, B1 => n40751, B2 => 
                           n49097, ZN => n48496);
   U2183 : AOI22_X1 port map( A1 => n40743, A2 => n40576, B1 => n40686, B2 => 
                           n49016, ZN => n48495);
   U2184 : AOI22_X1 port map( A1 => n41148, A2 => n40586, B1 => n40679, B2 => 
                           n40574, ZN => n48494);
   U2185 : AOI22_X1 port map( A1 => n41418, A2 => n40585, B1 => n41399, B2 => 
                           n40582, ZN => n48493);
   U2186 : NAND4_X1 port map( A1 => n48496, A2 => n48495, A3 => n48494, A4 => 
                           n48493, ZN => n48502);
   U2187 : AOI22_X1 port map( A1 => n41401, A2 => n48962, B1 => n41397, B2 => 
                           n40583, ZN => n48500);
   U2188 : AOI22_X1 port map( A1 => n41400, A2 => n49024, B1 => n41426, B2 => 
                           n49026, ZN => n48499);
   U2189 : AOI22_X1 port map( A1 => n41419, A2 => n49096, B1 => n40721, B2 => 
                           n48785, ZN => n48498);
   U2190 : AOI22_X1 port map( A1 => n41396, A2 => n40581, B1 => n40773, B2 => 
                           n48968, ZN => n48497);
   U2191 : NAND4_X1 port map( A1 => n48500, A2 => n48499, A3 => n48498, A4 => 
                           n48497, ZN => n48501);
   U2192 : NOR2_X1 port map( A1 => n48502, A2 => n48501, ZN => n48514);
   U2193 : AOI22_X1 port map( A1 => n40771, A2 => n49063, B1 => n40772, B2 => 
                           n48883, ZN => n48506);
   U2194 : AOI22_X1 port map( A1 => n40776, A2 => n49056, B1 => n40777, B2 => 
                           n48792, ZN => n48505);
   U2195 : AOI22_X1 port map( A1 => n40775, A2 => n40568, B1 => n40774, B2 => 
                           n40648, ZN => n48504);
   U2196 : AOI22_X1 port map( A1 => n40666, A2 => n41687, B1 => n40674, B2 => 
                           n49064, ZN => n48503);
   U2197 : NAND4_X1 port map( A1 => n48506, A2 => n48505, A3 => n48504, A4 => 
                           n48503, ZN => n48512);
   U2198 : AOI22_X1 port map( A1 => n41406, A2 => n48792, B1 => n41010, B2 => 
                           n40571, ZN => n48510);
   U2199 : AOI22_X1 port map( A1 => n41414, A2 => n40655, B1 => n40990, B2 => 
                           n49057, ZN => n48509);
   U2200 : AOI22_X1 port map( A1 => n41415, A2 => n49063, B1 => n41018, B2 => 
                           n48979, ZN => n48508);
   U2201 : AOI22_X1 port map( A1 => n41416, A2 => n40654, B1 => n41114, B2 => 
                           n41689, ZN => n48507);
   U2202 : NAND4_X1 port map( A1 => n48510, A2 => n48509, A3 => n48508, A4 => 
                           n48507, ZN => n48511);
   U2203 : AOI22_X1 port map( A1 => n48869, A2 => n48512, B1 => n48578, B2 => 
                           n48511, ZN => n48513);
   U2204 : OAI21_X1 port map( B1 => n49012, B2 => n48514, A => n48513, ZN => 
                           OUT1(24));
   U2205 : AOI22_X1 port map( A1 => n41154, A2 => n49024, B1 => n41081, B2 => 
                           n40576, ZN => n48518);
   U2206 : AOI22_X1 port map( A1 => n41053, A2 => n40584, B1 => n41134, B2 => 
                           n48967, ZN => n48517);
   U2207 : AOI22_X1 port map( A1 => n41427, A2 => n40580, B1 => n41092, B2 => 
                           n48785, ZN => n48516);
   U2208 : AOI22_X1 port map( A1 => n41135, A2 => n40581, B1 => n41133, B2 => 
                           n49025, ZN => n48515);
   U2209 : NAND4_X1 port map( A1 => n48518, A2 => n48517, A3 => n48516, A4 => 
                           n48515, ZN => n48524);
   U2210 : AOI22_X1 port map( A1 => n41188, A2 => n48992, B1 => n41042, B2 => 
                           n49013, ZN => n48522);
   U2211 : AOI22_X1 port map( A1 => n41147, A2 => n47431, B1 => n41166, B2 => 
                           n40582, ZN => n48521);
   U2212 : AOI22_X1 port map( A1 => n41095, A2 => n49097, B1 => n41093, B2 => 
                           n49016, ZN => n48520);
   U2213 : AOI22_X1 port map( A1 => n41245, A2 => n40585, B1 => n41358, B2 => 
                           n48758, ZN => n48519);
   U2214 : NAND4_X1 port map( A1 => n48522, A2 => n48521, A3 => n48520, A4 => 
                           n48519, ZN => n48523);
   U2215 : NOR2_X1 port map( A1 => n48524, A2 => n48523, ZN => n48536);
   U2216 : AOI22_X1 port map( A1 => n41474, A2 => n49063, B1 => n41507, B2 => 
                           n49055, ZN => n48528);
   U2217 : AOI22_X1 port map( A1 => n41490, A2 => n41690, B1 => n41476, B2 => 
                           n41692, ZN => n48527);
   U2218 : AOI22_X1 port map( A1 => n41495, A2 => n41686, B1 => n41477, B2 => 
                           n48792, ZN => n48526);
   U2219 : AOI22_X1 port map( A1 => n41494, A2 => n41687, B1 => n41471, B2 => 
                           n41688, ZN => n48525);
   U2220 : NAND4_X1 port map( A1 => n48528, A2 => n48527, A3 => n48526, A4 => 
                           n48525, ZN => n48534);
   U2221 : AOI22_X1 port map( A1 => n41481, A2 => n49063, B1 => n41058, B2 => 
                           n48979, ZN => n48532);
   U2222 : AOI22_X1 port map( A1 => n41045, A2 => n41690, B1 => n41323, B2 => 
                           n40654, ZN => n48531);
   U2223 : AOI22_X1 port map( A1 => n41051, A2 => n41687, B1 => n41121, B2 => 
                           n41689, ZN => n48530);
   U2224 : AOI22_X1 port map( A1 => n41472, A2 => n40655, B1 => n41240, B2 => 
                           n49062, ZN => n48529);
   U2225 : NAND4_X1 port map( A1 => n48532, A2 => n48531, A3 => n48530, A4 => 
                           n48529, ZN => n48533);
   U2226 : AOI22_X1 port map( A1 => n48869, A2 => n48534, B1 => n48578, B2 => 
                           n48533, ZN => n48535);
   U2227 : OAI21_X1 port map( B1 => n49075, B2 => n48536, A => n48535, ZN => 
                           OUT1(23));
   U2228 : AOI22_X1 port map( A1 => n41137, A2 => n49015, B1 => n41138, B2 => 
                           n49025, ZN => n48540);
   U2229 : AOI22_X1 port map( A1 => n41165, A2 => n40582, B1 => n41136, B2 => 
                           n40586, ZN => n48539);
   U2230 : AOI22_X1 port map( A1 => n41089, A2 => n49016, B1 => n41073, B2 => 
                           n49097, ZN => n48538);
   U2231 : AOI22_X1 port map( A1 => n41072, A2 => n48968, B1 => n41244, B2 => 
                           n49023, ZN => n48537);
   U2232 : NAND4_X1 port map( A1 => n48540, A2 => n48539, A3 => n48538, A4 => 
                           n48537, ZN => n48546);
   U2233 : AOI22_X1 port map( A1 => n41044, A2 => n49013, B1 => n41359, B2 => 
                           n48758, ZN => n48544);
   U2234 : AOI22_X1 port map( A1 => n41082, A2 => n40576, B1 => n41195, B2 => 
                           n48992, ZN => n48543);
   U2235 : AOI22_X1 port map( A1 => n41428, A2 => n49026, B1 => n41146, B2 => 
                           n48962, ZN => n48542);
   U2236 : AOI22_X1 port map( A1 => n41153, A2 => n40587, B1 => n41060, B2 => 
                           n48785, ZN => n48541);
   U2237 : NAND4_X1 port map( A1 => n48544, A2 => n48543, A3 => n48542, A4 => 
                           n48541, ZN => n48545);
   U2238 : NOR2_X1 port map( A1 => n48546, A2 => n48545, ZN => n48558);
   U2239 : AOI22_X1 port map( A1 => n41484, A2 => n49057, B1 => n41478, B2 => 
                           n48883, ZN => n48550);
   U2240 : AOI22_X1 port map( A1 => n41483, A2 => n41686, B1 => n41482, B2 => 
                           n49055, ZN => n48549);
   U2241 : AOI22_X1 port map( A1 => n41473, A2 => n49056, B1 => n41485, B2 => 
                           n49064, ZN => n48548);
   U2242 : AOI22_X1 port map( A1 => n41480, A2 => n48792, B1 => n41475, B2 => 
                           n49063, ZN => n48547);
   U2243 : NAND4_X1 port map( A1 => n48550, A2 => n48549, A3 => n48548, A4 => 
                           n48547, ZN => n48556);
   U2244 : AOI22_X1 port map( A1 => n41113, A2 => n40648, B1 => n41486, B2 => 
                           n49084, ZN => n48554);
   U2245 : AOI22_X1 port map( A1 => n41488, A2 => n48883, B1 => n41246, B2 => 
                           n48792, ZN => n48553);
   U2246 : AOI22_X1 port map( A1 => n41052, A2 => n41687, B1 => n41059, B2 => 
                           n41686, ZN => n48552);
   U2247 : AOI22_X1 port map( A1 => n41046, A2 => n41690, B1 => n41319, B2 => 
                           n40654, ZN => n48551);
   U2248 : NAND4_X1 port map( A1 => n48554, A2 => n48553, A3 => n48552, A4 => 
                           n48551, ZN => n48555);
   U2249 : AOI22_X1 port map( A1 => n48869, A2 => n48556, B1 => n48578, B2 => 
                           n48555, ZN => n48557);
   U2250 : OAI21_X1 port map( B1 => n49075, B2 => n48558, A => n48557, ZN => 
                           OUT1(22));
   U2251 : AOI22_X1 port map( A1 => n40722, A2 => n49095, B1 => n40685, B2 => 
                           n47430, ZN => n48562);
   U2252 : AOI22_X1 port map( A1 => n41355, A2 => n40582, B1 => n41357, B2 => 
                           n48962, ZN => n48561);
   U2253 : AOI22_X1 port map( A1 => n41367, A2 => n49096, B1 => n41356, B2 => 
                           n40587, ZN => n48560);
   U2254 : AOI22_X1 port map( A1 => n40715, A2 => n49013, B1 => n41429, B2 => 
                           n40580, ZN => n48559);
   U2255 : NAND4_X1 port map( A1 => n48562, A2 => n48561, A3 => n48560, A4 => 
                           n48559, ZN => n48568);
   U2256 : AOI22_X1 port map( A1 => n41352, A2 => n40586, B1 => n40757, B2 => 
                           n49097, ZN => n48566);
   U2257 : AOI22_X1 port map( A1 => n41368, A2 => n49015, B1 => n41353, B2 => 
                           n49025, ZN => n48565);
   U2258 : AOI22_X1 port map( A1 => n41366, A2 => n40585, B1 => n41354, B2 => 
                           n40577, ZN => n48564);
   U2259 : AOI22_X1 port map( A1 => n40737, A2 => n40576, B1 => n40704, B2 => 
                           n40584, ZN => n48563);
   U2260 : NAND4_X1 port map( A1 => n48566, A2 => n48565, A3 => n48564, A4 => 
                           n48563, ZN => n48567);
   U2261 : NOR2_X1 port map( A1 => n48568, A2 => n48567, ZN => n48581);
   U2262 : AOI22_X1 port map( A1 => n40855, A2 => n48883, B1 => n40848, B2 => 
                           n40571, ZN => n48572);
   U2263 : AOI22_X1 port map( A1 => n40850, A2 => n40649, B1 => n40854, B2 => 
                           n48792, ZN => n48571);
   U2264 : AOI22_X1 port map( A1 => n40851, A2 => n48979, B1 => n40856, B2 => 
                           n49084, ZN => n48570);
   U2265 : AOI22_X1 port map( A1 => n40857, A2 => n41688, B1 => n40853, B2 => 
                           n41689, ZN => n48569);
   U2266 : NAND4_X1 port map( A1 => n48572, A2 => n48571, A3 => n48570, A4 => 
                           n48569, ZN => n48579);
   U2267 : AOI22_X1 port map( A1 => n41363, A2 => n48883, B1 => n41004, B2 => 
                           n41690, ZN => n48576);
   U2268 : AOI22_X1 port map( A1 => n41364, A2 => n49063, B1 => n41111, B2 => 
                           n41689, ZN => n48575);
   U2269 : AOI22_X1 port map( A1 => n41362, A2 => n48792, B1 => n41365, B2 => 
                           n41688, ZN => n48574);
   U2270 : AOI22_X1 port map( A1 => n41015, A2 => n41686, B1 => n41031, B2 => 
                           n40649, ZN => n48573);
   U2271 : NAND4_X1 port map( A1 => n48576, A2 => n48575, A3 => n48574, A4 => 
                           n48573, ZN => n48577);
   U2272 : AOI22_X1 port map( A1 => n48869, A2 => n48579, B1 => n48578, B2 => 
                           n48577, ZN => n48580);
   U2273 : OAI21_X1 port map( B1 => n49075, B2 => n48581, A => n48580, ZN => 
                           OUT1(21));
   U2274 : AOI22_X1 port map( A1 => n41152, A2 => n40587, B1 => n41243, B2 => 
                           n40585, ZN => n48585);
   U2275 : AOI22_X1 port map( A1 => n41099, A2 => n47430, B1 => n41074, B2 => 
                           n40584, ZN => n48584);
   U2276 : AOI22_X1 port map( A1 => n41061, A2 => n49095, B1 => n41086, B2 => 
                           n40574, ZN => n48583);
   U2277 : AOI22_X1 port map( A1 => n41127, A2 => n48967, B1 => n41196, B2 => 
                           n40577, ZN => n48582);
   U2278 : NAND4_X1 port map( A1 => n48585, A2 => n48584, A3 => n48583, A4 => 
                           n48582, ZN => n48591);
   U2279 : AOI22_X1 port map( A1 => n41360, A2 => n49096, B1 => n41132, B2 => 
                           n40581, ZN => n48589);
   U2280 : AOI22_X1 port map( A1 => n41126, A2 => n49025, B1 => n41145, B2 => 
                           n48962, ZN => n48588);
   U2281 : AOI22_X1 port map( A1 => n41100, A2 => n40576, B1 => n41164, B2 => 
                           n40582, ZN => n48587);
   U2282 : AOI22_X1 port map( A1 => n41430, A2 => n40580, B1 => n41101, B2 => 
                           n49097, ZN => n48586);
   U2283 : NAND4_X1 port map( A1 => n48589, A2 => n48588, A3 => n48587, A4 => 
                           n48586, ZN => n48590);
   U2284 : NOR2_X1 port map( A1 => n48591, A2 => n48590, ZN => n48603);
   U2285 : AOI22_X1 port map( A1 => n41462, A2 => n40649, B1 => n41459, B2 => 
                           n49083, ZN => n48595);
   U2286 : AOI22_X1 port map( A1 => n41464, A2 => n40655, B1 => n41468, B2 => 
                           n40571, ZN => n48594);
   U2287 : AOI22_X1 port map( A1 => n41470, A2 => n40568, B1 => n41460, B2 => 
                           n49084, ZN => n48593);
   U2288 : AOI22_X1 port map( A1 => n41467, A2 => n40648, B1 => n41461, B2 => 
                           n49056, ZN => n48592);
   U2289 : NAND4_X1 port map( A1 => n48595, A2 => n48594, A3 => n48593, A4 => 
                           n48592, ZN => n48601);
   U2290 : AOI22_X1 port map( A1 => n41247, A2 => n49062, B1 => n41318, B2 => 
                           n40654, ZN => n48599);
   U2291 : AOI22_X1 port map( A1 => n41583, A2 => n49055, B1 => n41491, B2 => 
                           n48883, ZN => n48598);
   U2292 : AOI22_X1 port map( A1 => n41545, A2 => n40571, B1 => n41541, B2 => 
                           n40568, ZN => n48597);
   U2293 : AOI22_X1 port map( A1 => n41538, A2 => n49057, B1 => n41530, B2 => 
                           n49003, ZN => n48596);
   U2294 : NAND4_X1 port map( A1 => n48599, A2 => n48598, A3 => n48597, A4 => 
                           n48596, ZN => n48600);
   U2295 : AOI22_X1 port map( A1 => n48869, A2 => n48601, B1 => n49070, B2 => 
                           n48600, ZN => n48602);
   U2296 : OAI21_X1 port map( B1 => n49075, B2 => n48603, A => n48602, ZN => 
                           OUT1(20));
   U2297 : AOI22_X1 port map( A1 => n40723, A2 => n49095, B1 => n41144, B2 => 
                           n47431, ZN => n48607);
   U2298 : AOI22_X1 port map( A1 => n41129, A2 => n49025, B1 => n40683, B2 => 
                           n47430, ZN => n48606);
   U2299 : AOI22_X1 port map( A1 => n40731, A2 => n49022, B1 => n41130, B2 => 
                           n40586, ZN => n48605);
   U2300 : AOI22_X1 port map( A1 => n41131, A2 => n40581, B1 => n40712, B2 => 
                           n40574, ZN => n48604);
   U2301 : NAND4_X1 port map( A1 => n48607, A2 => n48606, A3 => n48605, A4 => 
                           n48604, ZN => n48613);
   U2302 : AOI22_X1 port map( A1 => n41197, A2 => n40577, B1 => n41163, B2 => 
                           n40582, ZN => n48611);
   U2303 : AOI22_X1 port map( A1 => n40700, A2 => n48968, B1 => n41361, B2 => 
                           n48758, ZN => n48610);
   U2304 : AOI22_X1 port map( A1 => n41242, A2 => n49023, B1 => n41431, B2 => 
                           n40580, ZN => n48609);
   U2305 : AOI22_X1 port map( A1 => n40750, A2 => n49097, B1 => n41151, B2 => 
                           n49024, ZN => n48608);
   U2306 : NAND4_X1 port map( A1 => n48611, A2 => n48610, A3 => n48609, A4 => 
                           n48608, ZN => n48612);
   U2307 : NOR2_X1 port map( A1 => n48613, A2 => n48612, ZN => n48625);
   U2308 : AOI22_X1 port map( A1 => n40866, A2 => n41689, B1 => n40852, B2 => 
                           n48792, ZN => n48617);
   U2309 : AOI22_X1 port map( A1 => n40868, A2 => n40655, B1 => n40869, B2 => 
                           n49084, ZN => n48616);
   U2310 : AOI22_X1 port map( A1 => n40865, A2 => n40568, B1 => n40849, B2 => 
                           n49057, ZN => n48615);
   U2311 : AOI22_X1 port map( A1 => n40837, A2 => n49064, B1 => n40867, B2 => 
                           n40654, ZN => n48614);
   U2312 : NAND4_X1 port map( A1 => n48617, A2 => n48616, A3 => n48615, A4 => 
                           n48614, ZN => n48623);
   U2313 : AOI22_X1 port map( A1 => n41106, A2 => n49055, B1 => n41012, B2 => 
                           n41690, ZN => n48621);
   U2314 : AOI22_X1 port map( A1 => n41014, A2 => n48979, B1 => n41339, B2 => 
                           n49084, ZN => n48620);
   U2315 : AOI22_X1 port map( A1 => n41285, A2 => n40655, B1 => n41017, B2 => 
                           n49057, ZN => n48619);
   U2316 : AOI22_X1 port map( A1 => n41248, A2 => n49062, B1 => n41317, B2 => 
                           n49056, ZN => n48618);
   U2317 : NAND4_X1 port map( A1 => n48621, A2 => n48620, A3 => n48619, A4 => 
                           n48618, ZN => n48622);
   U2318 : AOI22_X1 port map( A1 => n48869, A2 => n48623, B1 => n49070, B2 => 
                           n48622, ZN => n48624);
   U2319 : OAI21_X1 port map( B1 => n49075, B2 => n48625, A => n48624, ZN => 
                           OUT1(19));
   U2320 : AOI22_X1 port map( A1 => n41198, A2 => n40577, B1 => n41143, B2 => 
                           n47431, ZN => n48629);
   U2321 : AOI22_X1 port map( A1 => n41232, A2 => n49023, B1 => n40708, B2 => 
                           n40574, ZN => n48628);
   U2322 : AOI22_X1 port map( A1 => n40699, A2 => n48968, B1 => n41150, B2 => 
                           n40587, ZN => n48627);
   U2323 : AOI22_X1 port map( A1 => n40724, A2 => n49095, B1 => n41432, B2 => 
                           n40580, ZN => n48626);
   U2324 : NAND4_X1 port map( A1 => n48629, A2 => n48628, A3 => n48627, A4 => 
                           n48626, ZN => n48635);
   U2325 : AOI22_X1 port map( A1 => n41139, A2 => n48967, B1 => n40747, B2 => 
                           n49097, ZN => n48633);
   U2326 : AOI22_X1 port map( A1 => n40680, A2 => n47430, B1 => n40729, B2 => 
                           n40576, ZN => n48632);
   U2327 : AOI22_X1 port map( A1 => n41369, A2 => n49096, B1 => n41140, B2 => 
                           n49015, ZN => n48631);
   U2328 : AOI22_X1 port map( A1 => n41141, A2 => n40583, B1 => n41162, B2 => 
                           n49014, ZN => n48630);
   U2329 : NAND4_X1 port map( A1 => n48633, A2 => n48632, A3 => n48631, A4 => 
                           n48630, ZN => n48634);
   U2330 : NOR2_X1 port map( A1 => n48635, A2 => n48634, ZN => n48647);
   U2331 : AOI22_X1 port map( A1 => n40861, A2 => n49083, B1 => n40822, B2 => 
                           n40571, ZN => n48639);
   U2332 : AOI22_X1 port map( A1 => n40864, A2 => n49056, B1 => n40859, B2 => 
                           n48979, ZN => n48638);
   U2333 : AOI22_X1 port map( A1 => n40862, A2 => n41692, B1 => n40858, B2 => 
                           n41687, ZN => n48637);
   U2334 : AOI22_X1 port map( A1 => n40860, A2 => n41689, B1 => n40863, B2 => 
                           n49084, ZN => n48636);
   U2335 : NAND4_X1 port map( A1 => n48639, A2 => n48638, A3 => n48637, A4 => 
                           n48636, ZN => n48645);
   U2336 : AOI22_X1 port map( A1 => n41250, A2 => n49083, B1 => n41286, B2 => 
                           n40655, ZN => n48643);
   U2337 : AOI22_X1 port map( A1 => n41013, A2 => n41686, B1 => n41023, B2 => 
                           n40649, ZN => n48642);
   U2338 : AOI22_X1 port map( A1 => n41118, A2 => n49055, B1 => n41316, B2 => 
                           n41688, ZN => n48641);
   U2339 : AOI22_X1 port map( A1 => n40993, A2 => n49064, B1 => n41340, B2 => 
                           n49063, ZN => n48640);
   U2340 : NAND4_X1 port map( A1 => n48643, A2 => n48642, A3 => n48641, A4 => 
                           n48640, ZN => n48644);
   U2341 : AOI22_X1 port map( A1 => n48869, A2 => n48645, B1 => n49070, B2 => 
                           n48644, ZN => n48646);
   U2342 : OAI21_X1 port map( B1 => n49075, B2 => n48647, A => n48646, ZN => 
                           OUT1(18));
   U2343 : AOI22_X1 port map( A1 => n40695, A2 => n49097, B1 => n40678, B2 => 
                           n47430, ZN => n48651);
   U2344 : AOI22_X1 port map( A1 => n40702, A2 => n40574, B1 => n41384, B2 => 
                           n48962, ZN => n48650);
   U2345 : AOI22_X1 port map( A1 => n41383, A2 => n40587, B1 => n41380, B2 => 
                           n40583, ZN => n48649);
   U2346 : AOI22_X1 port map( A1 => n41391, A2 => n40585, B1 => n41379, B2 => 
                           n40586, ZN => n48648);
   U2347 : NAND4_X1 port map( A1 => n48651, A2 => n48650, A3 => n48649, A4 => 
                           n48648, ZN => n48657);
   U2348 : AOI22_X1 port map( A1 => n41392, A2 => n49096, B1 => n41420, B2 => 
                           n49026, ZN => n48655);
   U2349 : AOI22_X1 port map( A1 => n40698, A2 => n40584, B1 => n40734, B2 => 
                           n48785, ZN => n48654);
   U2350 : AOI22_X1 port map( A1 => n41381, A2 => n48992, B1 => n41377, B2 => 
                           n40581, ZN => n48653);
   U2351 : AOI22_X1 port map( A1 => n41382, A2 => n49014, B1 => n40727, B2 => 
                           n49022, ZN => n48652);
   U2352 : NAND4_X1 port map( A1 => n48655, A2 => n48654, A3 => n48653, A4 => 
                           n48652, ZN => n48656);
   U2353 : NOR2_X1 port map( A1 => n48657, A2 => n48656, ZN => n48669);
   U2354 : AOI22_X1 port map( A1 => n40938, A2 => n48979, B1 => n40933, B2 => 
                           n49084, ZN => n48661);
   U2355 : AOI22_X1 port map( A1 => n40935, A2 => n41688, B1 => n40931, B2 => 
                           n48792, ZN => n48660);
   U2356 : AOI22_X1 port map( A1 => n40830, A2 => n40571, B1 => n40937, B2 => 
                           n41687, ZN => n48659);
   U2357 : AOI22_X1 port map( A1 => n40939, A2 => n40655, B1 => n40929, B2 => 
                           n40648, ZN => n48658);
   U2358 : NAND4_X1 port map( A1 => n48661, A2 => n48660, A3 => n48659, A4 => 
                           n48658, ZN => n48667);
   U2359 : AOI22_X1 port map( A1 => n41557, A2 => n40571, B1 => n41388, B2 => 
                           n41692, ZN => n48665);
   U2360 : AOI22_X1 port map( A1 => n41390, A2 => n40654, B1 => n41584, B2 => 
                           n40648, ZN => n48664);
   U2361 : AOI22_X1 port map( A1 => n41389, A2 => n49063, B1 => n41539, B2 => 
                           n41687, ZN => n48663);
   U2362 : AOI22_X1 port map( A1 => n41387, A2 => n49083, B1 => n41542, B2 => 
                           n41686, ZN => n48662);
   U2363 : NAND4_X1 port map( A1 => n48665, A2 => n48664, A3 => n48663, A4 => 
                           n48662, ZN => n48666);
   U2364 : AOI22_X1 port map( A1 => n48869, A2 => n48667, B1 => n49070, B2 => 
                           n48666, ZN => n48668);
   U2365 : OAI21_X1 port map( B1 => n49075, B2 => n48669, A => n48668, ZN => 
                           OUT1(17));
   U2366 : AOI22_X1 port map( A1 => n41434, A2 => n40580, B1 => n41438, B2 => 
                           n49015, ZN => n48673);
   U2367 : AOI22_X1 port map( A1 => n40694, A2 => n49013, B1 => n41417, B2 => 
                           n40583, ZN => n48672);
   U2368 : AOI22_X1 port map( A1 => n40736, A2 => n49095, B1 => n41412, B2 => 
                           n49023, ZN => n48671);
   U2369 : AOI22_X1 port map( A1 => n40728, A2 => n47430, B1 => n41425, B2 => 
                           n47431, ZN => n48670);
   U2370 : NAND4_X1 port map( A1 => n48673, A2 => n48672, A3 => n48671, A4 => 
                           n48670, ZN => n48679);
   U2371 : AOI22_X1 port map( A1 => n40697, A2 => n40584, B1 => n40754, B2 => 
                           n49097, ZN => n48677);
   U2372 : AOI22_X1 port map( A1 => n41413, A2 => n49096, B1 => n41437, B2 => 
                           n48967, ZN => n48676);
   U2373 : AOI22_X1 port map( A1 => n41423, A2 => n49024, B1 => n41411, B2 => 
                           n40577, ZN => n48675);
   U2374 : AOI22_X1 port map( A1 => n40726, A2 => n40576, B1 => n41422, B2 => 
                           n40582, ZN => n48674);
   U2375 : NAND4_X1 port map( A1 => n48677, A2 => n48676, A3 => n48675, A4 => 
                           n48674, ZN => n48678);
   U2376 : NOR2_X1 port map( A1 => n48679, A2 => n48678, ZN => n48691);
   U2377 : AOI22_X1 port map( A1 => n40934, A2 => n41690, B1 => n40847, B2 => 
                           n40654, ZN => n48683);
   U2378 : AOI22_X1 port map( A1 => n40841, A2 => n41686, B1 => n40840, B2 => 
                           n40649, ZN => n48682);
   U2379 : AOI22_X1 port map( A1 => n40844, A2 => n41692, B1 => n40845, B2 => 
                           n49063, ZN => n48681);
   U2380 : AOI22_X1 port map( A1 => n40843, A2 => n49083, B1 => n40842, B2 => 
                           n41689, ZN => n48680);
   U2381 : NAND4_X1 port map( A1 => n48683, A2 => n48682, A3 => n48681, A4 => 
                           n48680, ZN => n48689);
   U2382 : AOI22_X1 port map( A1 => n41410, A2 => n40654, B1 => n41116, B2 => 
                           n40648, ZN => n48687);
   U2383 : AOI22_X1 port map( A1 => n41005, A2 => n40571, B1 => n41022, B2 => 
                           n41687, ZN => n48686);
   U2384 : AOI22_X1 port map( A1 => n41409, A2 => n49063, B1 => n41407, B2 => 
                           n48792, ZN => n48685);
   U2385 : AOI22_X1 port map( A1 => n41408, A2 => n40655, B1 => n41009, B2 => 
                           n40568, ZN => n48684);
   U2386 : NAND4_X1 port map( A1 => n48687, A2 => n48686, A3 => n48685, A4 => 
                           n48684, ZN => n48688);
   U2387 : AOI22_X1 port map( A1 => n48869, A2 => n48689, B1 => n49070, B2 => 
                           n48688, ZN => n48690);
   U2388 : OAI21_X1 port map( B1 => n49075, B2 => n48691, A => n48690, ZN => 
                           OUT1(16));
   U2389 : AOI22_X1 port map( A1 => n40701, A2 => n40574, B1 => n41176, B2 => 
                           n40587, ZN => n48695);
   U2390 : AOI22_X1 port map( A1 => n41231, A2 => n40585, B1 => n41199, B2 => 
                           n40577, ZN => n48694);
   U2391 : AOI22_X1 port map( A1 => n41177, A2 => n47431, B1 => n41370, B2 => 
                           n48758, ZN => n48693);
   U2392 : AOI22_X1 port map( A1 => n41175, A2 => n40582, B1 => n41178, B2 => 
                           n40583, ZN => n48692);
   U2393 : NAND4_X1 port map( A1 => n48695, A2 => n48694, A3 => n48693, A4 => 
                           n48692, ZN => n48701);
   U2394 : AOI22_X1 port map( A1 => n40725, A2 => n49022, B1 => n41173, B2 => 
                           n40581, ZN => n48699);
   U2395 : AOI22_X1 port map( A1 => n40738, A2 => n49095, B1 => n40677, B2 => 
                           n47430, ZN => n48698);
   U2396 : AOI22_X1 port map( A1 => n40749, A2 => n49097, B1 => n41174, B2 => 
                           n48967, ZN => n48697);
   U2397 : AOI22_X1 port map( A1 => n41433, A2 => n40580, B1 => n40696, B2 => 
                           n40584, ZN => n48696);
   U2398 : NAND4_X1 port map( A1 => n48699, A2 => n48698, A3 => n48697, A4 => 
                           n48696, ZN => n48700);
   U2399 : NOR2_X1 port map( A1 => n48701, A2 => n48700, ZN => n48713);
   U2400 : AOI22_X1 port map( A1 => n40904, A2 => n40649, B1 => n40891, B2 => 
                           n48883, ZN => n48705);
   U2401 : AOI22_X1 port map( A1 => n40882, A2 => n40648, B1 => n40893, B2 => 
                           n48979, ZN => n48704);
   U2402 : AOI22_X1 port map( A1 => n40888, A2 => n49063, B1 => n40887, B2 => 
                           n40654, ZN => n48703);
   U2403 : AOI22_X1 port map( A1 => n40892, A2 => n49083, B1 => n40799, B2 => 
                           n40571, ZN => n48702);
   U2404 : NAND4_X1 port map( A1 => n48705, A2 => n48704, A3 => n48703, A4 => 
                           n48702, ZN => n48711);
   U2405 : AOI22_X1 port map( A1 => n41251, A2 => n49083, B1 => n41341, B2 => 
                           n49063, ZN => n48709);
   U2406 : AOI22_X1 port map( A1 => n41540, A2 => n49057, B1 => n41556, B2 => 
                           n41686, ZN => n48708);
   U2407 : AOI22_X1 port map( A1 => n41580, A2 => n41689, B1 => n41287, B2 => 
                           n48883, ZN => n48707);
   U2408 : AOI22_X1 port map( A1 => n41554, A2 => n49064, B1 => n41315, B2 => 
                           n49056, ZN => n48706);
   U2409 : NAND4_X1 port map( A1 => n48709, A2 => n48708, A3 => n48707, A4 => 
                           n48706, ZN => n48710);
   U2410 : AOI22_X1 port map( A1 => n48869, A2 => n48711, B1 => n49070, B2 => 
                           n48710, ZN => n48712);
   U2411 : OAI21_X1 port map( B1 => n49075, B2 => n48713, A => n48712, ZN => 
                           OUT1(15));
   U2412 : AOI22_X1 port map( A1 => n41179, A2 => n40583, B1 => n41142, B2 => 
                           n47431, ZN => n48717);
   U2413 : AOI22_X1 port map( A1 => n40692, A2 => n48968, B1 => n41200, B2 => 
                           n40577, ZN => n48716);
   U2414 : AOI22_X1 port map( A1 => n41371, A2 => n49096, B1 => n40761, B2 => 
                           n49097, ZN => n48715);
   U2415 : AOI22_X1 port map( A1 => n41229, A2 => n40585, B1 => n41125, B2 => 
                           n48967, ZN => n48714);
   U2416 : NAND4_X1 port map( A1 => n48717, A2 => n48716, A3 => n48715, A4 => 
                           n48714, ZN => n48723);
   U2417 : AOI22_X1 port map( A1 => n40740, A2 => n49095, B1 => n41128, B2 => 
                           n40581, ZN => n48721);
   U2418 : AOI22_X1 port map( A1 => n41149, A2 => n40587, B1 => n40684, B2 => 
                           n47430, ZN => n48720);
   U2419 : AOI22_X1 port map( A1 => n41436, A2 => n49026, B1 => n40717, B2 => 
                           n49022, ZN => n48719);
   U2420 : AOI22_X1 port map( A1 => n41158, A2 => n40582, B1 => n40703, B2 => 
                           n49013, ZN => n48718);
   U2421 : NAND4_X1 port map( A1 => n48721, A2 => n48720, A3 => n48719, A4 => 
                           n48718, ZN => n48722);
   U2422 : NOR2_X1 port map( A1 => n48723, A2 => n48722, ZN => n48735);
   U2423 : AOI22_X1 port map( A1 => n40801, A2 => n49083, B1 => n40795, B2 => 
                           n40568, ZN => n48727);
   U2424 : AOI22_X1 port map( A1 => n40797, A2 => n49056, B1 => n40802, B2 => 
                           n49055, ZN => n48726);
   U2425 : AOI22_X1 port map( A1 => n40925, A2 => n49064, B1 => n40796, B2 => 
                           n49057, ZN => n48725);
   U2426 : AOI22_X1 port map( A1 => n40798, A2 => n49063, B1 => n40800, B2 => 
                           n40655, ZN => n48724);
   U2427 : NAND4_X1 port map( A1 => n48727, A2 => n48726, A3 => n48725, A4 => 
                           n48724, ZN => n48733);
   U2428 : AOI22_X1 port map( A1 => n41342, A2 => n49063, B1 => n41007, B2 => 
                           n40568, ZN => n48731);
   U2429 : AOI22_X1 port map( A1 => n41254, A2 => n49083, B1 => n41294, B2 => 
                           n48883, ZN => n48730);
   U2430 : AOI22_X1 port map( A1 => n41124, A2 => n49055, B1 => n41028, B2 => 
                           n49064, ZN => n48729);
   U2431 : AOI22_X1 port map( A1 => n41030, A2 => n49057, B1 => n41314, B2 => 
                           n40654, ZN => n48728);
   U2432 : NAND4_X1 port map( A1 => n48731, A2 => n48730, A3 => n48729, A4 => 
                           n48728, ZN => n48732);
   U2433 : AOI22_X1 port map( A1 => n48869, A2 => n48733, B1 => n49070, B2 => 
                           n48732, ZN => n48734);
   U2434 : OAI21_X1 port map( B1 => n49075, B2 => n48735, A => n48734, ZN => 
                           OUT1(14));
   U2435 : AOI22_X1 port map( A1 => n41187, A2 => n47431, B1 => n41201, B2 => 
                           n40577, ZN => n48739);
   U2436 : AOI22_X1 port map( A1 => n40745, A2 => n49016, B1 => n41228, B2 => 
                           n49023, ZN => n48738);
   U2437 : AOI22_X1 port map( A1 => n40716, A2 => n40576, B1 => n41435, B2 => 
                           n40580, ZN => n48737);
   U2438 : AOI22_X1 port map( A1 => n40762, A2 => n49097, B1 => n41373, B2 => 
                           n48758, ZN => n48736);
   U2439 : NAND4_X1 port map( A1 => n48739, A2 => n48738, A3 => n48737, A4 => 
                           n48736, ZN => n48745);
   U2440 : AOI22_X1 port map( A1 => n41186, A2 => n40587, B1 => n41182, B2 => 
                           n40581, ZN => n48743);
   U2441 : AOI22_X1 port map( A1 => n41185, A2 => n40582, B1 => n41184, B2 => 
                           n40583, ZN => n48742);
   U2442 : AOI22_X1 port map( A1 => n40742, A2 => n49095, B1 => n40705, B2 => 
                           n49013, ZN => n48741);
   U2443 : AOI22_X1 port map( A1 => n41183, A2 => n40586, B1 => n40691, B2 => 
                           n48968, ZN => n48740);
   U2444 : NAND4_X1 port map( A1 => n48743, A2 => n48742, A3 => n48741, A4 => 
                           n48740, ZN => n48744);
   U2445 : NOR2_X1 port map( A1 => n48745, A2 => n48744, ZN => n48757);
   U2446 : AOI22_X1 port map( A1 => n40815, A2 => n41690, B1 => n40816, B2 => 
                           n40649, ZN => n48749);
   U2447 : AOI22_X1 port map( A1 => n40817, A2 => n41686, B1 => n40810, B2 => 
                           n49063, ZN => n48748);
   U2448 : AOI22_X1 port map( A1 => n40819, A2 => n49083, B1 => n40811, B2 => 
                           n41688, ZN => n48747);
   U2449 : AOI22_X1 port map( A1 => n40809, A2 => n40655, B1 => n40818, B2 => 
                           n49055, ZN => n48746);
   U2450 : NAND4_X1 port map( A1 => n48749, A2 => n48748, A3 => n48747, A4 => 
                           n48746, ZN => n48755);
   U2451 : AOI22_X1 port map( A1 => n41255, A2 => n49083, B1 => n41343, B2 => 
                           n49063, ZN => n48753);
   U2452 : AOI22_X1 port map( A1 => n40994, A2 => n48979, B1 => n41011, B2 => 
                           n40571, ZN => n48752);
   U2453 : AOI22_X1 port map( A1 => n41297, A2 => n41692, B1 => n41001, B2 => 
                           n40649, ZN => n48751);
   U2454 : AOI22_X1 port map( A1 => n41308, A2 => n41688, B1 => n41117, B2 => 
                           n40648, ZN => n48750);
   U2455 : NAND4_X1 port map( A1 => n48753, A2 => n48752, A3 => n48751, A4 => 
                           n48750, ZN => n48754);
   U2456 : AOI22_X1 port map( A1 => n48869, A2 => n48755, B1 => n49070, B2 => 
                           n48754, ZN => n48756);
   U2457 : OAI21_X1 port map( B1 => n49075, B2 => n48757, A => n48756, ZN => 
                           OUT1(13));
   U2458 : AOI22_X1 port map( A1 => n41227, A2 => n49023, B1 => n41374, B2 => 
                           n48758, ZN => n48762);
   U2459 : AOI22_X1 port map( A1 => n40690, A2 => n40584, B1 => n40714, B2 => 
                           n40576, ZN => n48761);
   U2460 : AOI22_X1 port map( A1 => n41193, A2 => n40587, B1 => n41194, B2 => 
                           n47431, ZN => n48760);
   U2461 : AOI22_X1 port map( A1 => n40744, A2 => n49097, B1 => n41192, B2 => 
                           n49014, ZN => n48759);
   U2462 : NAND4_X1 port map( A1 => n48762, A2 => n48761, A3 => n48760, A4 => 
                           n48759, ZN => n48768);
   U2463 : AOI22_X1 port map( A1 => n40706, A2 => n40574, B1 => n41439, B2 => 
                           n40580, ZN => n48766);
   U2464 : AOI22_X1 port map( A1 => n40756, A2 => n49095, B1 => n41202, B2 => 
                           n48992, ZN => n48765);
   U2465 : AOI22_X1 port map( A1 => n41189, A2 => n40581, B1 => n40748, B2 => 
                           n47430, ZN => n48764);
   U2466 : AOI22_X1 port map( A1 => n41190, A2 => n40586, B1 => n41191, B2 => 
                           n49025, ZN => n48763);
   U2467 : NAND4_X1 port map( A1 => n48766, A2 => n48765, A3 => n48764, A4 => 
                           n48763, ZN => n48767);
   U2468 : NOR2_X1 port map( A1 => n48768, A2 => n48767, ZN => n48780);
   U2469 : AOI22_X1 port map( A1 => n40828, A2 => n49083, B1 => n40829, B2 => 
                           n48883, ZN => n48772);
   U2470 : AOI22_X1 port map( A1 => n40827, A2 => n41689, B1 => n40820, B2 => 
                           n49063, ZN => n48771);
   U2471 : AOI22_X1 port map( A1 => n40826, A2 => n40568, B1 => n40825, B2 => 
                           n49057, ZN => n48770);
   U2472 : AOI22_X1 port map( A1 => n40824, A2 => n49064, B1 => n40821, B2 => 
                           n40654, ZN => n48769);
   U2473 : NAND4_X1 port map( A1 => n48772, A2 => n48771, A3 => n48770, A4 => 
                           n48769, ZN => n48778);
   U2474 : AOI22_X1 port map( A1 => n41307, A2 => n41688, B1 => n41256, B2 => 
                           n48792, ZN => n48776);
   U2475 : AOI22_X1 port map( A1 => n41344, A2 => n49063, B1 => n41032, B2 => 
                           n41690, ZN => n48775);
   U2476 : AOI22_X1 port map( A1 => n41109, A2 => n40648, B1 => n41003, B2 => 
                           n40568, ZN => n48774);
   U2477 : AOI22_X1 port map( A1 => n41033, A2 => n40649, B1 => n41298, B2 => 
                           n48883, ZN => n48773);
   U2478 : NAND4_X1 port map( A1 => n48776, A2 => n48775, A3 => n48774, A4 => 
                           n48773, ZN => n48777);
   U2479 : AOI22_X1 port map( A1 => n48869, A2 => n48778, B1 => n49070, B2 => 
                           n48777, ZN => n48779);
   U2480 : OAI21_X1 port map( B1 => n49075, B2 => n48780, A => n48779, ZN => 
                           OUT1(12));
   U2481 : AOI22_X1 port map( A1 => n41207, A2 => n49014, B1 => n41226, B2 => 
                           n40585, ZN => n48784);
   U2482 : AOI22_X1 port map( A1 => n40707, A2 => n40574, B1 => n41378, B2 => 
                           n49026, ZN => n48783);
   U2483 : AOI22_X1 port map( A1 => n41375, A2 => n49096, B1 => n40760, B2 => 
                           n49097, ZN => n48782);
   U2484 : AOI22_X1 port map( A1 => n41203, A2 => n40581, B1 => n40752, B2 => 
                           n49016, ZN => n48781);
   U2485 : NAND4_X1 port map( A1 => n48784, A2 => n48783, A3 => n48782, A4 => 
                           n48781, ZN => n48791);
   U2486 : AOI22_X1 port map( A1 => n40713, A2 => n49022, B1 => n41209, B2 => 
                           n48962, ZN => n48789);
   U2487 : AOI22_X1 port map( A1 => n41205, A2 => n40583, B1 => n41206, B2 => 
                           n48992, ZN => n48788);
   U2488 : AOI22_X1 port map( A1 => n41204, A2 => n40586, B1 => n41693, B2 => 
                           n40584, ZN => n48787);
   U2489 : AOI22_X1 port map( A1 => n41208, A2 => n49024, B1 => n40732, B2 => 
                           n48785, ZN => n48786);
   U2490 : NAND4_X1 port map( A1 => n48789, A2 => n48788, A3 => n48787, A4 => 
                           n48786, ZN => n48790);
   U2491 : NOR2_X1 port map( A1 => n48791, A2 => n48790, ZN => n48804);
   U2492 : AOI22_X1 port map( A1 => n40836, A2 => n49055, B1 => n40838, B2 => 
                           n48792, ZN => n48796);
   U2493 : AOI22_X1 port map( A1 => n40846, A2 => n49084, B1 => n40835, B2 => 
                           n48979, ZN => n48795);
   U2494 : AOI22_X1 port map( A1 => n40832, A2 => n49056, B1 => n40834, B2 => 
                           n41687, ZN => n48794);
   U2495 : AOI22_X1 port map( A1 => n40839, A2 => n48883, B1 => n40833, B2 => 
                           n49064, ZN => n48793);
   U2496 : NAND4_X1 port map( A1 => n48796, A2 => n48795, A3 => n48794, A4 => 
                           n48793, ZN => n48802);
   U2497 : AOI22_X1 port map( A1 => n41110, A2 => n41689, B1 => n41345, B2 => 
                           n49063, ZN => n48800);
   U2498 : AOI22_X1 port map( A1 => n41257, A2 => n49083, B1 => n41303, B2 => 
                           n41692, ZN => n48799);
   U2499 : AOI22_X1 port map( A1 => n41019, A2 => n40571, B1 => n40999, B2 => 
                           n41687, ZN => n48798);
   U2500 : AOI22_X1 port map( A1 => n41002, A2 => n48979, B1 => n41306, B2 => 
                           n49056, ZN => n48797);
   U2501 : NAND4_X1 port map( A1 => n48800, A2 => n48799, A3 => n48798, A4 => 
                           n48797, ZN => n48801);
   U2502 : AOI22_X1 port map( A1 => n48869, A2 => n48802, B1 => n49070, B2 => 
                           n48801, ZN => n48803);
   U2503 : OAI21_X1 port map( B1 => n49075, B2 => n48804, A => n48803, ZN => 
                           OUT1(11));
   U2504 : AOI22_X1 port map( A1 => n41217, A2 => n48962, B1 => n40988, B2 => 
                           n49095, ZN => n48808);
   U2505 : AOI22_X1 port map( A1 => n40986, A2 => n40574, B1 => n41216, B2 => 
                           n40587, ZN => n48807);
   U2506 : AOI22_X1 port map( A1 => n41213, A2 => n49025, B1 => n40983, B2 => 
                           n40584, ZN => n48806);
   U2507 : AOI22_X1 port map( A1 => n40985, A2 => n49016, B1 => n41376, B2 => 
                           n49096, ZN => n48805);
   U2508 : NAND4_X1 port map( A1 => n48808, A2 => n48807, A3 => n48806, A4 => 
                           n48805, ZN => n48814);
   U2509 : AOI22_X1 port map( A1 => n41451, A2 => n48967, B1 => n41212, B2 => 
                           n40581, ZN => n48812);
   U2510 : AOI22_X1 port map( A1 => n41172, A2 => n49026, B1 => n41214, B2 => 
                           n48992, ZN => n48811);
   U2511 : AOI22_X1 port map( A1 => n40984, A2 => n40576, B1 => n41215, B2 => 
                           n49014, ZN => n48810);
   U2512 : AOI22_X1 port map( A1 => n41225, A2 => n40585, B1 => n40987, B2 => 
                           n49097, ZN => n48809);
   U2513 : NAND4_X1 port map( A1 => n48812, A2 => n48811, A3 => n48810, A4 => 
                           n48809, ZN => n48813);
   U2514 : NOR2_X1 port map( A1 => n48814, A2 => n48813, ZN => n48826);
   U2515 : AOI22_X1 port map( A1 => n41453, A2 => n40649, B1 => n41443, B2 => 
                           n41692, ZN => n48818);
   U2516 : AOI22_X1 port map( A1 => n41449, A2 => n49083, B1 => n41448, B2 => 
                           n49003, ZN => n48817);
   U2517 : AOI22_X1 port map( A1 => n41450, A2 => n40568, B1 => n41452, B2 => 
                           n40571, ZN => n48816);
   U2518 : AOI22_X1 port map( A1 => n41446, A2 => n40648, B1 => n41445, B2 => 
                           n40654, ZN => n48815);
   U2519 : NAND4_X1 port map( A1 => n48818, A2 => n48817, A3 => n48816, A4 => 
                           n48815, ZN => n48824);
   U2520 : AOI22_X1 port map( A1 => n41260, A2 => n49083, B1 => n41026, B2 => 
                           n49057, ZN => n48822);
   U2521 : AOI22_X1 port map( A1 => n41348, A2 => n49084, B1 => n41447, B2 => 
                           n40654, ZN => n48821);
   U2522 : AOI22_X1 port map( A1 => n41016, A2 => n49064, B1 => n41112, B2 => 
                           n40648, ZN => n48820);
   U2523 : AOI22_X1 port map( A1 => n41444, A2 => n48883, B1 => n40992, B2 => 
                           n48979, ZN => n48819);
   U2524 : NAND4_X1 port map( A1 => n48822, A2 => n48821, A3 => n48820, A4 => 
                           n48819, ZN => n48823);
   U2525 : AOI22_X1 port map( A1 => n48869, A2 => n48824, B1 => n49070, B2 => 
                           n48823, ZN => n48825);
   U2526 : OAI21_X1 port map( B1 => n49012, B2 => n48826, A => n48825, ZN => 
                           OUT1(10));
   U2527 : AOI22_X1 port map( A1 => n40689, A2 => n40584, B1 => n40753, B2 => 
                           n49016, ZN => n48830);
   U2528 : AOI22_X1 port map( A1 => n40741, A2 => n49097, B1 => n41171, B2 => 
                           n48967, ZN => n48829);
   U2529 : AOI22_X1 port map( A1 => n41210, A2 => n40577, B1 => n41218, B2 => 
                           n48962, ZN => n48828);
   U2530 : AOI22_X1 port map( A1 => n41224, A2 => n40585, B1 => n41167, B2 => 
                           n49015, ZN => n48827);
   U2531 : NAND4_X1 port map( A1 => n48830, A2 => n48829, A3 => n48828, A4 => 
                           n48827, ZN => n48836);
   U2532 : AOI22_X1 port map( A1 => n41168, A2 => n40580, B1 => n41170, B2 => 
                           n49014, ZN => n48834);
   U2533 : AOI22_X1 port map( A1 => n41169, A2 => n49024, B1 => n40733, B2 => 
                           n49095, ZN => n48833);
   U2534 : AOI22_X1 port map( A1 => n41385, A2 => n49096, B1 => n41180, B2 => 
                           n40583, ZN => n48832);
   U2535 : AOI22_X1 port map( A1 => n40709, A2 => n49013, B1 => n40711, B2 => 
                           n40576, ZN => n48831);
   U2536 : NAND4_X1 port map( A1 => n48834, A2 => n48833, A3 => n48832, A4 => 
                           n48831, ZN => n48835);
   U2537 : NOR2_X1 port map( A1 => n48836, A2 => n48835, ZN => n48848);
   U2538 : AOI22_X1 port map( A1 => n40766, A2 => n49062, B1 => n40767, B2 => 
                           n41687, ZN => n48840);
   U2539 : AOI22_X1 port map( A1 => n40769, A2 => n49056, B1 => n40768, B2 => 
                           n48883, ZN => n48839);
   U2540 : AOI22_X1 port map( A1 => n40764, A2 => n41689, B1 => n40765, B2 => 
                           n40568, ZN => n48838);
   U2541 : AOI22_X1 port map( A1 => n40770, A2 => n49084, B1 => n40763, B2 => 
                           n49064, ZN => n48837);
   U2542 : NAND4_X1 port map( A1 => n48840, A2 => n48839, A3 => n48838, A4 => 
                           n48837, ZN => n48846);
   U2543 : AOI22_X1 port map( A1 => n41262, A2 => n49083, B1 => n41304, B2 => 
                           n40655, ZN => n48844);
   U2544 : AOI22_X1 port map( A1 => n41347, A2 => n49084, B1 => n41122, B2 => 
                           n40648, ZN => n48843);
   U2545 : AOI22_X1 port map( A1 => n41300, A2 => n41688, B1 => n40991, B2 => 
                           n40571, ZN => n48842);
   U2546 : AOI22_X1 port map( A1 => n41000, A2 => n40568, B1 => n41025, B2 => 
                           n40649, ZN => n48841);
   U2547 : NAND4_X1 port map( A1 => n48844, A2 => n48843, A3 => n48842, A4 => 
                           n48841, ZN => n48845);
   U2548 : AOI22_X1 port map( A1 => n48869, A2 => n48846, B1 => n49070, B2 => 
                           n48845, ZN => n48847);
   U2549 : OAI21_X1 port map( B1 => n49075, B2 => n48848, A => n48847, ZN => 
                           OUT1(9));
   U2550 : AOI22_X1 port map( A1 => n41181, A2 => n40583, B1 => n40735, B2 => 
                           n49095, ZN => n48852);
   U2551 : AOI22_X1 port map( A1 => n41155, A2 => n40586, B1 => n41157, B2 => 
                           n49026, ZN => n48851);
   U2552 : AOI22_X1 port map( A1 => n41223, A2 => n40585, B1 => n40718, B2 => 
                           n40574, ZN => n48850);
   U2553 : AOI22_X1 port map( A1 => n41156, A2 => n49015, B1 => n41386, B2 => 
                           n49096, ZN => n48849);
   U2554 : NAND4_X1 port map( A1 => n48852, A2 => n48851, A3 => n48850, A4 => 
                           n48849, ZN => n48858);
   U2555 : AOI22_X1 port map( A1 => n40688, A2 => n40584, B1 => n41211, B2 => 
                           n40577, ZN => n48856);
   U2556 : AOI22_X1 port map( A1 => n40755, A2 => n47430, B1 => n41160, B2 => 
                           n49024, ZN => n48855);
   U2557 : AOI22_X1 port map( A1 => n40730, A2 => n49097, B1 => n40710, B2 => 
                           n49022, ZN => n48854);
   U2558 : AOI22_X1 port map( A1 => n41161, A2 => n49014, B1 => n41159, B2 => 
                           n47431, ZN => n48853);
   U2559 : NAND4_X1 port map( A1 => n48856, A2 => n48855, A3 => n48854, A4 => 
                           n48853, ZN => n48857);
   U2560 : NOR2_X1 port map( A1 => n48858, A2 => n48857, ZN => n48871);
   U2561 : AOI22_X1 port map( A1 => n40785, A2 => n49084, B1 => n40782, B2 => 
                           n41687, ZN => n48862);
   U2562 : AOI22_X1 port map( A1 => n40778, A2 => n49056, B1 => n40783, B2 => 
                           n49055, ZN => n48861);
   U2563 : AOI22_X1 port map( A1 => n40779, A2 => n49062, B1 => n40781, B2 => 
                           n40571, ZN => n48860);
   U2564 : AOI22_X1 port map( A1 => n40780, A2 => n40568, B1 => n40784, B2 => 
                           n40655, ZN => n48859);
   U2565 : NAND4_X1 port map( A1 => n48862, A2 => n48861, A3 => n48860, A4 => 
                           n48859, ZN => n48868);
   U2566 : AOI22_X1 port map( A1 => n41264, A2 => n49062, B1 => n41024, B2 => 
                           n49064, ZN => n48866);
   U2567 : AOI22_X1 port map( A1 => n41299, A2 => n40654, B1 => n41029, B2 => 
                           n49057, ZN => n48865);
   U2568 : AOI22_X1 port map( A1 => n41120, A2 => n40648, B1 => n41346, B2 => 
                           n49003, ZN => n48864);
   U2569 : AOI22_X1 port map( A1 => n40997, A2 => n40568, B1 => n41305, B2 => 
                           n41692, ZN => n48863);
   U2570 : NAND4_X1 port map( A1 => n48866, A2 => n48865, A3 => n48864, A4 => 
                           n48863, ZN => n48867);
   U2571 : AOI22_X1 port map( A1 => n48869, A2 => n48868, B1 => n49070, B2 => 
                           n48867, ZN => n48870);
   U2572 : OAI21_X1 port map( B1 => n49075, B2 => n48871, A => n48870, ZN => 
                           OUT1(8));
   U2573 : AOI22_X1 port map( A1 => n41679, A2 => n48962, B1 => n41034, B2 => 
                           n49095, ZN => n48875);
   U2574 : AOI22_X1 port map( A1 => n41664, A2 => n49096, B1 => n41655, B2 => 
                           n40585, ZN => n48874);
   U2575 : AOI22_X1 port map( A1 => n41674, A2 => n40581, B1 => n41039, B2 => 
                           n40574, ZN => n48873);
   U2576 : AOI22_X1 port map( A1 => n41669, A2 => n40582, B1 => n41038, B2 => 
                           n49017, ZN => n48872);
   U2577 : NAND4_X1 port map( A1 => n48875, A2 => n48874, A3 => n48873, A4 => 
                           n48872, ZN => n48881);
   U2578 : AOI22_X1 port map( A1 => n41683, A2 => n40583, B1 => n41684, B2 => 
                           n40586, ZN => n48879);
   U2579 : AOI22_X1 port map( A1 => n41678, A2 => n40587, B1 => n41036, B2 => 
                           n49022, ZN => n48878);
   U2580 : AOI22_X1 port map( A1 => n41035, A2 => n48968, B1 => n41667, B2 => 
                           n40577, ZN => n48877);
   U2581 : AOI22_X1 port map( A1 => n41037, A2 => n47430, B1 => n41682, B2 => 
                           n49026, ZN => n48876);
   U2582 : NAND4_X1 port map( A1 => n48879, A2 => n48878, A3 => n48877, A4 => 
                           n48876, ZN => n48880);
   U2583 : NOR2_X1 port map( A1 => n48881, A2 => n48880, ZN => n48895);
   U2584 : CLKBUF_X1 port map( A => n48882, Z => n49072);
   U2585 : AOI22_X1 port map( A1 => n41463, A2 => n48883, B1 => n41455, B2 => 
                           n49062, ZN => n48887);
   U2586 : AOI22_X1 port map( A1 => n41456, A2 => n49084, B1 => n41458, B2 => 
                           n40649, ZN => n48886);
   U2587 : AOI22_X1 port map( A1 => n41466, A2 => n41689, B1 => n41457, B2 => 
                           n41688, ZN => n48885);
   U2588 : AOI22_X1 port map( A1 => n41465, A2 => n48979, B1 => n41469, B2 => 
                           n40571, ZN => n48884);
   U2589 : NAND4_X1 port map( A1 => n48887, A2 => n48886, A3 => n48885, A4 => 
                           n48884, ZN => n48893);
   U2590 : AOI22_X1 port map( A1 => n41547, A2 => n49064, B1 => n41616, B2 => 
                           n41688, ZN => n48891);
   U2591 : AOI22_X1 port map( A1 => n41578, A2 => n49055, B1 => n41550, B2 => 
                           n41687, ZN => n48890);
   U2592 : AOI22_X1 port map( A1 => n41591, A2 => n41692, B1 => n41681, B2 => 
                           n49062, ZN => n48889);
   U2593 : AOI22_X1 port map( A1 => n41552, A2 => n48979, B1 => n41588, B2 => 
                           n49003, ZN => n48888);
   U2594 : NAND4_X1 port map( A1 => n48891, A2 => n48890, A3 => n48889, A4 => 
                           n48888, ZN => n48892);
   U2595 : AOI22_X1 port map( A1 => n49072, A2 => n48893, B1 => n49070, B2 => 
                           n48892, ZN => n48894);
   U2596 : OAI21_X1 port map( B1 => n49075, B2 => n48895, A => n48894, ZN => 
                           OUT1(7));
   U2597 : AOI22_X1 port map( A1 => n41654, A2 => n40581, B1 => n41652, B2 => 
                           n49024, ZN => n48899);
   U2598 : AOI22_X1 port map( A1 => n41676, A2 => n40582, B1 => n41658, B2 => 
                           n49096, ZN => n48898);
   U2599 : AOI22_X1 port map( A1 => n40976, A2 => n40574, B1 => n41648, B2 => 
                           n40577, ZN => n48897);
   U2600 : AOI22_X1 port map( A1 => n41653, A2 => n40586, B1 => n40957, B2 => 
                           n49017, ZN => n48896);
   U2601 : NAND4_X1 port map( A1 => n48899, A2 => n48898, A3 => n48897, A4 => 
                           n48896, ZN => n48905);
   U2602 : AOI22_X1 port map( A1 => n41651, A2 => n40583, B1 => n40966, B2 => 
                           n40576, ZN => n48903);
   U2603 : AOI22_X1 port map( A1 => n41680, A2 => n40580, B1 => n40948, B2 => 
                           n49016, ZN => n48902);
   U2604 : AOI22_X1 port map( A1 => n41661, A2 => n49023, B1 => n40974, B2 => 
                           n40584, ZN => n48901);
   U2605 : AOI22_X1 port map( A1 => n41673, A2 => n47431, B1 => n40958, B2 => 
                           n49095, ZN => n48900);
   U2606 : NAND4_X1 port map( A1 => n48903, A2 => n48902, A3 => n48901, A4 => 
                           n48900, ZN => n48904);
   U2607 : NOR2_X1 port map( A1 => n48905, A2 => n48904, ZN => n48917);
   U2608 : AOI22_X1 port map( A1 => n40884, A2 => n49084, B1 => n40890, B2 => 
                           n41686, ZN => n48909);
   U2609 : AOI22_X1 port map( A1 => n40883, A2 => n41692, B1 => n40881, B2 => 
                           n49062, ZN => n48908);
   U2610 : AOI22_X1 port map( A1 => n40885, A2 => n40654, B1 => n40919, B2 => 
                           n49064, ZN => n48907);
   U2611 : AOI22_X1 port map( A1 => n40898, A2 => n49057, B1 => n40880, B2 => 
                           n40648, ZN => n48906);
   U2612 : NAND4_X1 port map( A1 => n48909, A2 => n48908, A3 => n48907, A4 => 
                           n48906, ZN => n48915);
   U2613 : AOI22_X1 port map( A1 => n41561, A2 => n40649, B1 => n41587, B2 => 
                           n49003, ZN => n48913);
   U2614 : AOI22_X1 port map( A1 => n41562, A2 => n48979, B1 => n41546, B2 => 
                           n40571, ZN => n48912);
   U2615 : AOI22_X1 port map( A1 => n41662, A2 => n49056, B1 => n41582, B2 => 
                           n40648, ZN => n48911);
   U2616 : AOI22_X1 port map( A1 => n41597, A2 => n40655, B1 => n41663, B2 => 
                           n49062, ZN => n48910);
   U2617 : NAND4_X1 port map( A1 => n48913, A2 => n48912, A3 => n48911, A4 => 
                           n48910, ZN => n48914);
   U2618 : AOI22_X1 port map( A1 => n49072, A2 => n48915, B1 => n49070, B2 => 
                           n48914, ZN => n48916);
   U2619 : OAI21_X1 port map( B1 => n49075, B2 => n48917, A => n48916, ZN => 
                           OUT1(6));
   U2620 : AOI22_X1 port map( A1 => n40950, A2 => n48968, B1 => n41656, B2 => 
                           n40585, ZN => n48921);
   U2621 : AOI22_X1 port map( A1 => n40970, A2 => n49097, B1 => n40979, B2 => 
                           n40574, ZN => n48920);
   U2622 : AOI22_X1 port map( A1 => n40965, A2 => n40576, B1 => n41629, B2 => 
                           n40577, ZN => n48919);
   U2623 : AOI22_X1 port map( A1 => n40951, A2 => n47430, B1 => n41641, B2 => 
                           n40580, ZN => n48918);
   U2624 : NAND4_X1 port map( A1 => n48921, A2 => n48920, A3 => n48919, A4 => 
                           n48918, ZN => n48927);
   U2625 : AOI22_X1 port map( A1 => n41642, A2 => n47431, B1 => n41645, B2 => 
                           n40582, ZN => n48925);
   U2626 : AOI22_X1 port map( A1 => n40968, A2 => n49095, B1 => n41631, B2 => 
                           n48967, ZN => n48924);
   U2627 : AOI22_X1 port map( A1 => n41633, A2 => n40581, B1 => n41650, B2 => 
                           n49025, ZN => n48923);
   U2628 : AOI22_X1 port map( A1 => n41634, A2 => n49096, B1 => n41644, B2 => 
                           n40587, ZN => n48922);
   U2629 : NAND4_X1 port map( A1 => n48925, A2 => n48924, A3 => n48923, A4 => 
                           n48922, ZN => n48926);
   U2630 : NOR2_X1 port map( A1 => n48927, A2 => n48926, ZN => n48939);
   U2631 : AOI22_X1 port map( A1 => n40894, A2 => n40571, B1 => n40886, B2 => 
                           n41688, ZN => n48931);
   U2632 : AOI22_X1 port map( A1 => n40897, A2 => n41687, B1 => n40889, B2 => 
                           n40568, ZN => n48930);
   U2633 : AOI22_X1 port map( A1 => n40877, A2 => n49083, B1 => n40879, B2 => 
                           n40648, ZN => n48929);
   U2634 : AOI22_X1 port map( A1 => n40876, A2 => n40655, B1 => n40878, B2 => 
                           n49003, ZN => n48928);
   U2635 : NAND4_X1 port map( A1 => n48931, A2 => n48930, A3 => n48929, A4 => 
                           n48928, ZN => n48937);
   U2636 : AOI22_X1 port map( A1 => n41639, A2 => n40654, B1 => n41581, B2 => 
                           n49055, ZN => n48935);
   U2637 : AOI22_X1 port map( A1 => n41564, A2 => n41690, B1 => n41637, B2 => 
                           n49062, ZN => n48934);
   U2638 : AOI22_X1 port map( A1 => n41592, A2 => n49084, B1 => n41565, B2 => 
                           n40568, ZN => n48933);
   U2639 : AOI22_X1 port map( A1 => n41593, A2 => n41692, B1 => n41551, B2 => 
                           n40649, ZN => n48932);
   U2640 : NAND4_X1 port map( A1 => n48935, A2 => n48934, A3 => n48933, A4 => 
                           n48932, ZN => n48936);
   U2641 : AOI22_X1 port map( A1 => n49072, A2 => n48937, B1 => n49070, B2 => 
                           n48936, ZN => n48938);
   U2642 : OAI21_X1 port map( B1 => n49012, B2 => n48939, A => n48938, ZN => 
                           OUT1(5));
   U2643 : AOI22_X1 port map( A1 => n40973, A2 => n49097, B1 => n40964, B2 => 
                           n40576, ZN => n48943);
   U2644 : AOI22_X1 port map( A1 => n40969, A2 => n49013, B1 => n40972, B2 => 
                           n48968, ZN => n48942);
   U2645 : AOI22_X1 port map( A1 => n41601, A2 => n49096, B1 => n41624, B2 => 
                           n40580, ZN => n48941);
   U2646 : AOI22_X1 port map( A1 => n41649, A2 => n49025, B1 => n41622, B2 => 
                           n49024, ZN => n48940);
   U2647 : NAND4_X1 port map( A1 => n48943, A2 => n48942, A3 => n48941, A4 => 
                           n48940, ZN => n48949);
   U2648 : AOI22_X1 port map( A1 => n41606, A2 => n40586, B1 => n41602, B2 => 
                           n40581, ZN => n48947);
   U2649 : AOI22_X1 port map( A1 => n41677, A2 => n49023, B1 => n41623, B2 => 
                           n40577, ZN => n48946);
   U2650 : AOI22_X1 port map( A1 => n41625, A2 => n47431, B1 => n40967, B2 => 
                           n49095, ZN => n48945);
   U2651 : AOI22_X1 port map( A1 => n40952, A2 => n49016, B1 => n41646, B2 => 
                           n40582, ZN => n48944);
   U2652 : NAND4_X1 port map( A1 => n48947, A2 => n48946, A3 => n48945, A4 => 
                           n48944, ZN => n48948);
   U2653 : NOR2_X1 port map( A1 => n48949, A2 => n48948, ZN => n48961);
   U2654 : AOI22_X1 port map( A1 => n40911, A2 => n40568, B1 => n40912, B2 => 
                           n49057, ZN => n48953);
   U2655 : AOI22_X1 port map( A1 => n40905, A2 => n41690, B1 => n40932, B2 => 
                           n49055, ZN => n48952);
   U2656 : AOI22_X1 port map( A1 => n40918, A2 => n49083, B1 => n40900, B2 => 
                           n49003, ZN => n48951);
   U2657 : AOI22_X1 port map( A1 => n40901, A2 => n40655, B1 => n40928, B2 => 
                           n49056, ZN => n48950);
   U2658 : NAND4_X1 port map( A1 => n48953, A2 => n48952, A3 => n48951, A4 => 
                           n48950, ZN => n48959);
   U2659 : AOI22_X1 port map( A1 => n41600, A2 => n41692, B1 => n41560, B2 => 
                           n41690, ZN => n48957);
   U2660 : AOI22_X1 port map( A1 => n41617, A2 => n41688, B1 => n41549, B2 => 
                           n41687, ZN => n48956);
   U2661 : AOI22_X1 port map( A1 => n41636, A2 => n49083, B1 => n41590, B2 => 
                           n49003, ZN => n48955);
   U2662 : AOI22_X1 port map( A1 => n41585, A2 => n40648, B1 => n41558, B2 => 
                           n48979, ZN => n48954);
   U2663 : NAND4_X1 port map( A1 => n48957, A2 => n48956, A3 => n48955, A4 => 
                           n48954, ZN => n48958);
   U2664 : AOI22_X1 port map( A1 => n49072, A2 => n48959, B1 => n49070, B2 => 
                           n48958, ZN => n48960);
   U2665 : OAI21_X1 port map( B1 => n49075, B2 => n48961, A => n48960, ZN => 
                           OUT1(4));
   U2666 : AOI22_X1 port map( A1 => n41614, A2 => n48962, B1 => n41608, B2 => 
                           n49096, ZN => n48966);
   U2667 : AOI22_X1 port map( A1 => n41620, A2 => n40587, B1 => n40953, B2 => 
                           n47430, ZN => n48965);
   U2668 : AOI22_X1 port map( A1 => n41675, A2 => n40585, B1 => n40947, B2 => 
                           n49017, ZN => n48964);
   U2669 : AOI22_X1 port map( A1 => n41610, A2 => n49015, B1 => n41621, B2 => 
                           n40577, ZN => n48963);
   U2670 : NAND4_X1 port map( A1 => n48966, A2 => n48965, A3 => n48964, A4 => 
                           n48963, ZN => n48974);
   U2671 : AOI22_X1 port map( A1 => n40962, A2 => n40576, B1 => n41643, B2 => 
                           n40583, ZN => n48972);
   U2672 : AOI22_X1 port map( A1 => n41611, A2 => n48967, B1 => n41647, B2 => 
                           n40582, ZN => n48971);
   U2673 : AOI22_X1 port map( A1 => n40981, A2 => n49095, B1 => n40975, B2 => 
                           n49013, ZN => n48970);
   U2674 : AOI22_X1 port map( A1 => n41613, A2 => n40580, B1 => n40978, B2 => 
                           n48968, ZN => n48969);
   U2675 : NAND4_X1 port map( A1 => n48972, A2 => n48971, A3 => n48970, A4 => 
                           n48969, ZN => n48973);
   U2676 : NOR2_X1 port map( A1 => n48974, A2 => n48973, ZN => n48987);
   U2677 : AOI22_X1 port map( A1 => n40907, A2 => n40654, B1 => n40909, B2 => 
                           n41692, ZN => n48978);
   U2678 : AOI22_X1 port map( A1 => n40896, A2 => n41686, B1 => n40916, B2 => 
                           n41690, ZN => n48977);
   U2679 : AOI22_X1 port map( A1 => n40899, A2 => n40649, B1 => n40910, B2 => 
                           n49062, ZN => n48976);
   U2680 : AOI22_X1 port map( A1 => n40908, A2 => n49084, B1 => n40895, B2 => 
                           n41689, ZN => n48975);
   U2681 : NAND4_X1 port map( A1 => n48978, A2 => n48977, A3 => n48976, A4 => 
                           n48975, ZN => n48985);
   U2682 : AOI22_X1 port map( A1 => n41555, A2 => n48979, B1 => n41596, B2 => 
                           n40655, ZN => n48983);
   U2683 : AOI22_X1 port map( A1 => n41544, A2 => n49057, B1 => n41635, B2 => 
                           n49062, ZN => n48982);
   U2684 : AOI22_X1 port map( A1 => n41548, A2 => n41690, B1 => n41577, B2 => 
                           n40648, ZN => n48981);
   U2685 : AOI22_X1 port map( A1 => n41598, A2 => n49084, B1 => n41626, B2 => 
                           n40654, ZN => n48980);
   U2686 : NAND4_X1 port map( A1 => n48983, A2 => n48982, A3 => n48981, A4 => 
                           n48980, ZN => n48984);
   U2687 : AOI22_X1 port map( A1 => n49072, A2 => n48985, B1 => n49070, B2 => 
                           n48984, ZN => n48986);
   U2688 : OAI21_X1 port map( B1 => n49075, B2 => n48987, A => n48986, ZN => 
                           OUT1(3));
   U2689 : AOI22_X1 port map( A1 => n40959, A2 => n40576, B1 => n40961, B2 => 
                           n49017, ZN => n48991);
   U2690 : AOI22_X1 port map( A1 => n40982, A2 => n49095, B1 => n41660, B2 => 
                           n40586, ZN => n48990);
   U2691 : AOI22_X1 port map( A1 => n41659, A2 => n49015, B1 => n41612, B2 => 
                           n49096, ZN => n48989);
   U2692 : AOI22_X1 port map( A1 => n41609, A2 => n40585, B1 => n40954, B2 => 
                           n47430, ZN => n48988);
   U2693 : NAND4_X1 port map( A1 => n48991, A2 => n48990, A3 => n48989, A4 => 
                           n48988, ZN => n48998);
   U2694 : AOI22_X1 port map( A1 => n41672, A2 => n40587, B1 => n40977, B2 => 
                           n40584, ZN => n48996);
   U2695 : AOI22_X1 port map( A1 => n41665, A2 => n47431, B1 => n41668, B2 => 
                           n48992, ZN => n48995);
   U2696 : AOI22_X1 port map( A1 => n41666, A2 => n49025, B1 => n41671, B2 => 
                           n40582, ZN => n48994);
   U2697 : AOI22_X1 port map( A1 => n40971, A2 => n40574, B1 => n41657, B2 => 
                           n40580, ZN => n48993);
   U2698 : NAND4_X1 port map( A1 => n48996, A2 => n48995, A3 => n48994, A4 => 
                           n48993, ZN => n48997);
   U2699 : NOR2_X1 port map( A1 => n48998, A2 => n48997, ZN => n49011);
   U2700 : AOI22_X1 port map( A1 => n40906, A2 => n40649, B1 => n40902, B2 => 
                           n49003, ZN => n49002);
   U2701 : AOI22_X1 port map( A1 => n40914, A2 => n40568, B1 => n40926, B2 => 
                           n49062, ZN => n49001);
   U2702 : AOI22_X1 port map( A1 => n40927, A2 => n40655, B1 => n40915, B2 => 
                           n49064, ZN => n49000);
   U2703 : AOI22_X1 port map( A1 => n40924, A2 => n49055, B1 => n40903, B2 => 
                           n49056, ZN => n48999);
   U2704 : NAND4_X1 port map( A1 => n49002, A2 => n49001, A3 => n49000, A4 => 
                           n48999, ZN => n49009);
   U2705 : AOI22_X1 port map( A1 => n41632, A2 => n49083, B1 => n41543, B2 => 
                           n41690, ZN => n49007);
   U2706 : AOI22_X1 port map( A1 => n41537, A2 => n40649, B1 => n41595, B2 => 
                           n49003, ZN => n49006);
   U2707 : AOI22_X1 port map( A1 => n41579, A2 => n40648, B1 => n41627, B2 => 
                           n49056, ZN => n49005);
   U2708 : AOI22_X1 port map( A1 => n41589, A2 => n41692, B1 => n41536, B2 => 
                           n40568, ZN => n49004);
   U2709 : NAND4_X1 port map( A1 => n49007, A2 => n49006, A3 => n49005, A4 => 
                           n49004, ZN => n49008);
   U2710 : AOI22_X1 port map( A1 => n49072, A2 => n49009, B1 => n49070, B2 => 
                           n49008, ZN => n49010);
   U2711 : OAI21_X1 port map( B1 => n49012, B2 => n49011, A => n49010, ZN => 
                           OUT1(2));
   U2712 : AOI22_X1 port map( A1 => n40980, A2 => n49013, B1 => n41604, B2 => 
                           n49096, ZN => n49021);
   U2713 : AOI22_X1 port map( A1 => n41605, A2 => n49015, B1 => n41670, B2 => 
                           n49014, ZN => n49020);
   U2714 : AOI22_X1 port map( A1 => n40963, A2 => n49095, B1 => n40956, B2 => 
                           n49016, ZN => n49019);
   U2715 : AOI22_X1 port map( A1 => n41619, A2 => n40577, B1 => n40960, B2 => 
                           n49017, ZN => n49018);
   U2716 : NAND4_X1 port map( A1 => n49021, A2 => n49020, A3 => n49019, A4 => 
                           n49018, ZN => n49032);
   U2717 : AOI22_X1 port map( A1 => n40949, A2 => n49022, B1 => n40955, B2 => 
                           n40584, ZN => n49030);
   U2718 : AOI22_X1 port map( A1 => n41618, A2 => n49024, B1 => n41603, B2 => 
                           n49023, ZN => n49029);
   U2719 : AOI22_X1 port map( A1 => n41615, A2 => n47431, B1 => n41607, B2 => 
                           n40586, ZN => n49028);
   U2720 : AOI22_X1 port map( A1 => n41640, A2 => n49026, B1 => n41638, B2 => 
                           n49025, ZN => n49027);
   U2721 : NAND4_X1 port map( A1 => n49030, A2 => n49029, A3 => n49028, A4 => 
                           n49027, ZN => n49031);
   U2722 : NOR2_X1 port map( A1 => n49032, A2 => n49031, ZN => n49044);
   U2723 : AOI22_X1 port map( A1 => n40913, A2 => n49084, B1 => n40923, B2 => 
                           n49057, ZN => n49036);
   U2724 : AOI22_X1 port map( A1 => n40917, A2 => n41692, B1 => n40930, B2 => 
                           n40654, ZN => n49035);
   U2725 : AOI22_X1 port map( A1 => n40920, A2 => n49083, B1 => n40922, B2 => 
                           n41686, ZN => n49034);
   U2726 : AOI22_X1 port map( A1 => n40921, A2 => n41689, B1 => n40936, B2 => 
                           n40571, ZN => n49033);
   U2727 : NAND4_X1 port map( A1 => n49036, A2 => n49035, A3 => n49034, A4 => 
                           n49033, ZN => n49042);
   U2728 : AOI22_X1 port map( A1 => n41563, A2 => n40568, B1 => n41559, B2 => 
                           n41687, ZN => n49040);
   U2729 : AOI22_X1 port map( A1 => n41594, A2 => n49084, B1 => n41630, B2 => 
                           n49083, ZN => n49039);
   U2730 : AOI22_X1 port map( A1 => n41628, A2 => n49056, B1 => n41586, B2 => 
                           n40648, ZN => n49038);
   U2731 : AOI22_X1 port map( A1 => n41599, A2 => n41692, B1 => n41553, B2 => 
                           n49064, ZN => n49037);
   U2732 : NAND4_X1 port map( A1 => n49040, A2 => n49039, A3 => n49038, A4 => 
                           n49037, ZN => n49041);
   U2733 : AOI22_X1 port map( A1 => n49072, A2 => n49042, B1 => n49070, B2 => 
                           n49041, ZN => n49043);
   U2734 : OAI21_X1 port map( B1 => n49075, B2 => n49044, A => n49043, ZN => 
                           OUT1(1));
   U2735 : AOI22_X1 port map( A1 => n41566, A2 => n40581, B1 => n40875, B2 => 
                           n49095, ZN => n49048);
   U2736 : AOI22_X1 port map( A1 => n41576, A2 => n40577, B1 => n40874, B2 => 
                           n47430, ZN => n49047);
   U2737 : AOI22_X1 port map( A1 => n41575, A2 => n40587, B1 => n41487, B2 => 
                           n49096, ZN => n49046);
   U2738 : AOI22_X1 port map( A1 => n40871, A2 => n40576, B1 => n41501, B2 => 
                           n40586, ZN => n49045);
   U2739 : NAND4_X1 port map( A1 => n49048, A2 => n49047, A3 => n49046, A4 => 
                           n49045, ZN => n49054);
   U2740 : AOI22_X1 port map( A1 => n41570, A2 => n40583, B1 => n41567, B2 => 
                           n40582, ZN => n49052);
   U2741 : AOI22_X1 port map( A1 => n41574, A2 => n47431, B1 => n41572, B2 => 
                           n40580, ZN => n49051);
   U2742 : AOI22_X1 port map( A1 => n40872, A2 => n49097, B1 => n40873, B2 => 
                           n40574, ZN => n49050);
   U2743 : AOI22_X1 port map( A1 => n40870, A2 => n40584, B1 => n41571, B2 => 
                           n40585, ZN => n49049);
   U2744 : NAND4_X1 port map( A1 => n49052, A2 => n49051, A3 => n49050, A4 => 
                           n49049, ZN => n49053);
   U2745 : NOR2_X1 port map( A1 => n49054, A2 => n49053, ZN => n49074);
   U2746 : AOI22_X1 port map( A1 => n40945, A2 => n49062, B1 => n40941, B2 => 
                           n49063, ZN => n49061);
   U2747 : AOI22_X1 port map( A1 => n40944, A2 => n49055, B1 => n41685, B2 => 
                           n41692, ZN => n49060);
   U2748 : AOI22_X1 port map( A1 => n40946, A2 => n49056, B1 => n40940, B2 => 
                           n40568, ZN => n49059);
   U2749 : AOI22_X1 port map( A1 => n40943, A2 => n49057, B1 => n40942, B2 => 
                           n41690, ZN => n49058);
   U2750 : NAND4_X1 port map( A1 => n49061, A2 => n49060, A3 => n49059, A4 => 
                           n49058, ZN => n49071);
   U2751 : AOI22_X1 port map( A1 => n41440, A2 => n40649, B1 => n41569, B2 => 
                           n49062, ZN => n49068);
   U2752 : AOI22_X1 port map( A1 => n41454, A2 => n41689, B1 => n41573, B2 => 
                           n49063, ZN => n49067);
   U2753 : AOI22_X1 port map( A1 => n41441, A2 => n40568, B1 => n41568, B2 => 
                           n41692, ZN => n49066);
   U2754 : AOI22_X1 port map( A1 => n41442, A2 => n49064, B1 => n41492, B2 => 
                           n41688, ZN => n49065);
   U2755 : NAND4_X1 port map( A1 => n49068, A2 => n49067, A3 => n49066, A4 => 
                           n49065, ZN => n49069);
   U2756 : AOI22_X1 port map( A1 => n49072, A2 => n49071, B1 => n49070, B2 => 
                           n49069, ZN => n49073);
   U2757 : OAI21_X1 port map( B1 => n49075, B2 => n49074, A => n49073, ZN => 
                           OUT1(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_17_port, curr_instruction_to_cu_i_16_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n151, cu_i_n135, 
      cu_i_N279, cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, 
      cu_i_N273, cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, 
      cu_i_cmd_alu_op_type_0_port, cu_i_cmd_alu_op_type_1_port, 
      cu_i_cmd_alu_op_type_2_port, cu_i_cmd_alu_op_type_3_port, 
      cu_i_cmd_word_3_port, cu_i_cmd_word_6_port, cu_i_cmd_word_8_port, 
      datapath_i_alu_output_val_i_0_port, datapath_i_alu_output_val_i_1_port, 
      datapath_i_alu_output_val_i_2_port, datapath_i_alu_output_val_i_3_port, 
      datapath_i_alu_output_val_i_4_port, datapath_i_alu_output_val_i_5_port, 
      datapath_i_alu_output_val_i_6_port, datapath_i_alu_output_val_i_7_port, 
      datapath_i_alu_output_val_i_8_port, datapath_i_alu_output_val_i_9_port, 
      datapath_i_alu_output_val_i_10_port, datapath_i_alu_output_val_i_11_port,
      datapath_i_alu_output_val_i_12_port, datapath_i_alu_output_val_i_13_port,
      datapath_i_alu_output_val_i_14_port, datapath_i_alu_output_val_i_15_port,
      datapath_i_alu_output_val_i_16_port, datapath_i_alu_output_val_i_17_port,
      datapath_i_alu_output_val_i_18_port, datapath_i_alu_output_val_i_19_port,
      datapath_i_alu_output_val_i_20_port, datapath_i_alu_output_val_i_21_port,
      datapath_i_alu_output_val_i_22_port, datapath_i_alu_output_val_i_23_port,
      datapath_i_alu_output_val_i_24_port, datapath_i_alu_output_val_i_25_port,
      datapath_i_alu_output_val_i_26_port, datapath_i_alu_output_val_i_27_port,
      datapath_i_alu_output_val_i_28_port, datapath_i_alu_output_val_i_29_port,
      datapath_i_alu_output_val_i_30_port, datapath_i_alu_output_val_i_31_port,
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_decode_stage_dp_n44, datapath_i_decode_stage_dp_n43, 
      datapath_i_decode_stage_dp_n42, datapath_i_decode_stage_dp_n41, 
      datapath_i_decode_stage_dp_n40, datapath_i_decode_stage_dp_n39, 
      datapath_i_decode_stage_dp_n38, datapath_i_decode_stage_dp_n37, 
      datapath_i_decode_stage_dp_n36, datapath_i_decode_stage_dp_n35, 
      datapath_i_decode_stage_dp_n34, datapath_i_decode_stage_dp_n33, 
      datapath_i_decode_stage_dp_n32, datapath_i_decode_stage_dp_n31, 
      datapath_i_decode_stage_dp_n30, datapath_i_decode_stage_dp_n29, 
      datapath_i_decode_stage_dp_n28, datapath_i_decode_stage_dp_n27, 
      datapath_i_decode_stage_dp_n26, datapath_i_decode_stage_dp_n25, 
      datapath_i_decode_stage_dp_n24, datapath_i_decode_stage_dp_n23, 
      datapath_i_decode_stage_dp_n22, datapath_i_decode_stage_dp_n21, 
      datapath_i_decode_stage_dp_n20, datapath_i_decode_stage_dp_n19, 
      datapath_i_decode_stage_dp_n18, datapath_i_decode_stage_dp_n17, 
      datapath_i_decode_stage_dp_n16, datapath_i_decode_stage_dp_n15, 
      datapath_i_decode_stage_dp_n14, datapath_i_decode_stage_dp_n13, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, n302, n474, n477, n492, n1443, 
      n1445, n1447, n1449, n1453, n1613, n1614, n1615, n1617, n1619, n1621, 
      n1623, n1625, n1627, n1629, n1631, n1633, n1635, n1637, n1639, n1641, 
      n1643, n1645, n1647, n1649, n1651, n1653, n1655, n1657, n1659, n1661, 
      n1663, n1665, n1667, n1669, n1671, n1673, n2299, n5478, n5479, n3284, 
      n3596, n4052, n4060, n4128, n4231, n4337, n4341, n4417, n5542, n4953, 
      n4954, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, 
      n4965, n4966, n4968, n4969, n4970, n4971, n4972, n4974, n4975, n4976, 
      n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, 
      n4987, n4989, n5006, n5009, n5010, n5011, n5012, n5013, n5014, n5015, 
      n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, 
      n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, 
      n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, 
      n5046, n5047, n5048, n5049, n5051, n5052, n5053, n5065, n5067, n5069, 
      n5071, n5073, n5075, n5076, n5077, n5079, n5084, n5085, n5089, n5092, 
      n5097, n5098, n5117, n5120, n5122, n5131, n5136, n5139, n5142, n5145, 
      n5148, n5151, n5154, n5157, n5160, n5163, n5166, n5169, n5172, n5175, 
      n5178, n5181, n5184, n5187, n5190, n5193, n5196, n5199, n5202, n5205, 
      n5208, n5211, n5214, n5217, n5220, n5223, n5226, n5229, n5285, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5358, n5388, n5405, 
      n5506, n5507, n5880, n6081, n6082, n6096, n6113, n6157, n6159, n6178, 
      n6207, n6209, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6783, n6784, 
      n6785, IRAM_ADDRESS_10_port, IRAM_ADDRESS_8_port, n6788, n6789, n6790, 
      n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, 
      n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, 
      n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, 
      n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6831, 
      n6832, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, 
      n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, 
      n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, 
      n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, 
      n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, 
      n6883, IRAM_ADDRESS_6_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, 
      n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6907, n6908, 
      n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, 
      n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, 
      n6929, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
      n6940, n6941, n6942, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
      n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
      n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, 
      n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, 
      n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, 
      n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, 
      n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, 
      n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, 
      n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, 
      n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7103, 
      n7104, n7106, n7107, n7109, n7110, n7112, n7113, n7114, n7115, n7117, 
      n7118, n7120, n7121, n7123, n7124, n7126, n7127, n7129, n7130, n7132, 
      n7133, n7135, n7136, n7138, n7139, n7141, n7142, n7144, n7145, n7147, 
      n7148, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, 
      n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7168, n7169, 
      n7170, n7171, n7172, IRAM_ADDRESS_2_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_9_port, IRAM_ADDRESS_7_port, n7179, n7180, n7181, n7182, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_19_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_29_port, n7193, n7194, n7195, n7196, n7197, n7198, n7199, 
      n7200, n7201, n7202, n7203, n7204, n7205, n7215, n7216, n7217, n7218, 
      n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, 
      n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, 
      n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, 
      n7249, n7250, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, 
      n7260, n7261, n7262, n7264, n7265, n7266, n7267, n7268, n7269, n7270, 
      IRAM_ADDRESS_31_port, n7274, n7275, n7277, n7307, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7333, n7334, 
      n7335, n7336, n7337, n7338, n7339, n7341, n7342, n7343, n7344, n7345, 
      n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, 
      n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, 
      n7366, n7367, n7369, n7525, n7526, n7527, n7528, n7529, n7530, n7531, 
      n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, 
      n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, 
      n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7694, n7695, n7696, 
      n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, 
      n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, 
      n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, 
      n7727, n7728, n7729, n7730, n7731, n7732, IRAM_ADDRESS_1_port, 
      IRAM_ADDRESS_0_port, n7735, n7736, n7737, n7738, n7739, n7740, n7741, 
      n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, 
      n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, 
      n7762, n7763, n7764, IRAM_ADDRESS_14_port, IRAM_ADDRESS_16_port, 
      IRAM_ADDRESS_18_port, IRAM_ADDRESS_20_port, IRAM_ADDRESS_22_port, 
      IRAM_ADDRESS_24_port, IRAM_ADDRESS_26_port, IRAM_ADDRESS_28_port, 
      IRAM_ADDRESS_30_port, n7774, n7775, n7776, n7777, n7778, n7779, n7780, 
      n7781, n7782, n7783, n7784, n7785, n7786, IRAM_ADDRESS_12_port, n7789, 
      n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, 
      n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, 
      n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, 
      n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, 
      n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, 
      n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, 
      n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, 
      n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, 
      n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, 
      n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, 
      n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, 
      n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, 
      n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, 
      n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, 
      n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, 
      n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, 
      n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, 
      n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, 
      n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, 
      n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, 
      n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, 
      n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, 
      n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, 
      n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, 
      n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, 
      n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, 
      n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, 
      n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, 
      n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, 
      n8080, n8081, n8082, n8083, n8084, n_3782, n_3783, n_3784, n_3785, n_3786
      , n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795,
      n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, 
      n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, 
      n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, 
      n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, 
      n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, 
      n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, 
      n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, 
      n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, 
      n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, 
      n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, 
      n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, 
      n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, 
      n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, 
      n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, 
      n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, 
      n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, 
      n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, 
      n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, 
      n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, 
      n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, 
      n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, 
      n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, 
      n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, 
      n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, 
      n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, 
      n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, 
      n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, 
      n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, 
      n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, 
      n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, 
      n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, 
      n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, 
      n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, 
      n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, 
      n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, 
      n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, 
      n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, 
      n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, 
      n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, 
      n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, 
      n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, 
      n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, 
      n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, 
      n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, 
      n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, 
      n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, 
      n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, 
      n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, 
      n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, 
      n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, 
      n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, 
      n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, 
      n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, 
      n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, 
      n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290 : 
      std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => n4417);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_n151);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => n5131);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n8076, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n8079, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n8079, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n8079, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n8079, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n8079, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n8079, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n8079, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n8079, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n8079, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n8079, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n8079, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n7193, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n7193, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n7193, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n7193, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n7193, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n8079, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n8076, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n8076, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n8076, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n8076, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n8076, Z 
                           => DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n8076, Z 
                           => DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n8076, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n8076, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n8076, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n8076, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n8076, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n8076, Z 
                           => DRAM_ADDRESS_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n7737, D => n7363, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n8082, D => n6897, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n8082, D => n6899, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n8082, D => n6898, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n7737, D => n6900, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n7737, D => n7257, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n7737, D => n6869, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n7737, D => n6870, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n7737, D => n6871, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n7737, D => n6872, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n7737, D => n6873, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n7737, D => n6889, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n7737, D => n6892, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n8082, D => n7268, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n8082, D => n6890, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n7737, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n7737, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n7737, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n7737, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n8082, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n7742, D => n7363, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n7742, D => n6897, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n8081, D => n6899, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n7742, D => n6898, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n8081, D => n6900, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n7742, D => n7257, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n8081, D => n6869, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n8081, D => n6870, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n7742, D => n6871, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n8081, D => n6872, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n7742, D => n6873, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n8081, D => n6889, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n7742, D => n6892, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n7742, D => n7268, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n7742, D => n6890, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n7742, D => n6887, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n8081, D => n6895, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n7742, D => n6893, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n7742, D => n7254, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n8081, D => n6891, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n7742, D => n6888, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n7742, D => n6874, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n7742, D => n6902, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n8081, D => n6881, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n7742, D => n6875, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n7742, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n7742, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n7742, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n7742, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n8081, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n7742, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n8081, D => n6876, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   clk_r_REG13304_S5 : DFFS_X1 port map( D => n7275, CK => CLK, SN => RST, Q =>
                           n7274, QN => n_3782);
   clk_r_REG11939_S5 : DFFR_X1 port map( D => n5478, CK => CLK, RN => RST, Q =>
                           n_3783, QN => n7311);
   clk_r_REG13281_S8 : DFFR_X1 port map( D => n5479, CK => CLK, RN => RST, Q =>
                           n_3784, QN => n7319);
   clk_r_REG11071_S15 : DFFR_X1 port map( D => n5542, CK => CLK, RN => RST, Q 
                           => IRAM_ADDRESS_31_port, QN => n_3785);
   clk_r_REG13440_S4 : DFFS_X1 port map( D => n7343, CK => CLK, SN => RST, Q =>
                           n7270, QN => n_3786);
   clk_r_REG13477_S6 : DFFR_X1 port map( D => n5388, CK => CLK, RN => RST, Q =>
                           n8066, QN => n7269);
   clk_r_REG13574_S7 : DFFR_X1 port map( D => n7752, CK => CLK, RN => RST, Q =>
                           n7268, QN => n_3787);
   clk_r_REG13534_S7 : DFFR_X1 port map( D => n7747, CK => CLK, RN => RST, Q =>
                           n7267, QN => n_3788);
   clk_r_REG13558_S7 : DFFR_X1 port map( D => n7746, CK => CLK, RN => RST, Q =>
                           n7266, QN => n_3789);
   clk_r_REG13557_S1 : DFFR_X1 port map( D => n7745, CK => CLK, RN => RST, Q =>
                           n7265, QN => n_3790);
   clk_r_REG13560_S7 : DFFR_X1 port map( D => n7741, CK => CLK, RN => RST, Q =>
                           n7264, QN => n_3791);
   clk_r_REG13428_S2 : DFFR_X1 port map( D => n7707, CK => CLK, RN => RST, Q =>
                           DRAM_READNOTWRITE, QN => n_3792);
   clk_r_REG11006_S15 : DFFS_X1 port map( D => n7785, CK => CLK, SN => RST, Q 
                           => n7262, QN => n_3793);
   clk_r_REG11119_S16 : DFFS_X1 port map( D => n7262, CK => CLK, SN => RST, Q 
                           => n7261, QN => n_3794);
   clk_r_REG11016_S15 : DFFS_X1 port map( D => n7784, CK => CLK, SN => RST, Q 
                           => n7260, QN => n_3795);
   clk_r_REG11112_S16 : DFFS_X1 port map( D => n7260, CK => CLK, SN => RST, Q 
                           => n7259, QN => n_3796);
   clk_r_REG13366_S1 : DFFR_X1 port map( D => n7744, CK => CLK, RN => RST, Q =>
                           n7258, QN => n_3797);
   clk_r_REG13565_S7 : DFFR_X1 port map( D => n7735, CK => CLK, RN => RST, Q =>
                           n7257, QN => n_3798);
   clk_r_REG11023_S15 : DFFS_X1 port map( D => n7783, CK => CLK, SN => RST, Q 
                           => n7256, QN => n_3799);
   clk_r_REG11106_S16 : DFFS_X1 port map( D => n7256, CK => CLK, SN => RST, Q 
                           => n7255, QN => n_3800);
   clk_r_REG13575_S7 : DFFR_X1 port map( D => n7756, CK => CLK, RN => RST, Q =>
                           n7254, QN => n_3801);
   clk_r_REG11034_S15 : DFFS_X1 port map( D => n7782, CK => CLK, SN => RST, Q 
                           => n7253, QN => n_3802);
   clk_r_REG11099_S16 : DFFS_X1 port map( D => n7253, CK => CLK, SN => RST, Q 
                           => n7252, QN => n_3803);
   clk_r_REG13631_S4 : DFFS_X1 port map( D => n7699, CK => CLK, SN => RST, Q =>
                           n_3804, QN => n7366);
   clk_r_REG13537_S3 : DFFR_X1 port map( D => n8080, CK => CLK, RN => RST, Q =>
                           n7249, QN => n_3805);
   clk_r_REG13533_S2 : DFFR_X1 port map( D => n8082, CK => CLK, RN => RST, Q =>
                           n7248, QN => n_3806);
   clk_r_REG11043_S15 : DFFS_X1 port map( D => n7781, CK => CLK, SN => RST, Q 
                           => n7247, QN => n_3807);
   clk_r_REG11093_S16 : DFFS_X1 port map( D => n7247, CK => CLK, SN => RST, Q 
                           => n7246, QN => n_3808);
   clk_r_REG11051_S15 : DFFS_X1 port map( D => n7780, CK => CLK, SN => RST, Q 
                           => n7245, QN => n_3809);
   clk_r_REG11087_S16 : DFFS_X1 port map( D => n7245, CK => CLK, SN => RST, Q 
                           => n7244, QN => n_3810);
   clk_r_REG11058_S15 : DFFS_X1 port map( D => n7779, CK => CLK, SN => RST, Q 
                           => n7243, QN => n_3811);
   clk_r_REG11081_S16 : DFFS_X1 port map( D => n7243, CK => CLK, SN => RST, Q 
                           => n7242, QN => n_3812);
   clk_r_REG11069_S15 : DFFS_X1 port map( D => n7732, CK => CLK, SN => RST, Q 
                           => n7241, QN => n_3813);
   clk_r_REG11073_S16 : DFFS_X1 port map( D => n7241, CK => CLK, SN => RST, Q 
                           => n7240, QN => n_3814);
   clk_r_REG11065_S15 : DFFS_X1 port map( D => n7778, CK => CLK, SN => RST, Q 
                           => n7239, QN => n_3815);
   clk_r_REG11074_S16 : DFFS_X1 port map( D => n7239, CK => CLK, SN => RST, Q 
                           => n7238, QN => n_3816);
   clk_r_REG11791_S6 : DFFR_X1 port map( D => n6207, CK => CLK, RN => RST, Q =>
                           n_3817, QN => n7237);
   clk_r_REG11793_S7 : DFFS_X1 port map( D => n7237, CK => CLK, SN => RST, Q =>
                           n7236, QN => n_3818);
   clk_r_REG11794_S8 : DFFS_X1 port map( D => n7236, CK => CLK, SN => RST, Q =>
                           n7235, QN => n_3819);
   clk_r_REG11650_S6 : DFFR_X1 port map( D => n6209, CK => CLK, RN => RST, Q =>
                           n_3820, QN => n7234);
   clk_r_REG11652_S7 : DFFS_X1 port map( D => n7234, CK => CLK, SN => RST, Q =>
                           n7233, QN => n_3821);
   clk_r_REG11653_S8 : DFFS_X1 port map( D => n7233, CK => CLK, SN => RST, Q =>
                           n7232, QN => n_3822);
   clk_r_REG11353_S6 : DFFR_X1 port map( D => n6113, CK => CLK, RN => RST, Q =>
                           n_3823, QN => n7231);
   clk_r_REG11355_S7 : DFFS_X1 port map( D => n7231, CK => CLK, SN => RST, Q =>
                           n7230, QN => n_3824);
   clk_r_REG11356_S8 : DFFS_X1 port map( D => n7230, CK => CLK, SN => RST, Q =>
                           n7229, QN => n_3825);
   clk_r_REG11367_S6 : DFFR_X1 port map( D => n6096, CK => CLK, RN => RST, Q =>
                           n_3826, QN => n7228);
   clk_r_REG11370_S7 : DFFS_X1 port map( D => n7228, CK => CLK, SN => RST, Q =>
                           n7227, QN => n_3827);
   clk_r_REG11371_S8 : DFFS_X1 port map( D => n7227, CK => CLK, SN => RST, Q =>
                           n7226, QN => n_3828);
   clk_r_REG10955_S13 : DFFS_X1 port map( D => n7762, CK => CLK, SN => RST, Q 
                           => n7225, QN => n_3829);
   clk_r_REG10956_S14 : DFFS_X1 port map( D => n7225, CK => CLK, SN => RST, Q 
                           => n7224, QN => n_3830);
   clk_r_REG10957_S15 : DFFS_X1 port map( D => n7224, CK => CLK, SN => RST, Q 
                           => n7223, QN => n_3831);
   clk_r_REG10966_S13 : DFFS_X1 port map( D => n7341, CK => CLK, SN => RST, Q 
                           => n7222, QN => n_3832);
   clk_r_REG10967_S14 : DFFS_X1 port map( D => n7222, CK => CLK, SN => RST, Q 
                           => n7221, QN => n_3833);
   clk_r_REG11153_S15 : DFFS_X1 port map( D => n7221, CK => CLK, SN => RST, Q 
                           => n7220, QN => n_3834);
   clk_r_REG10974_S14 : DFFS_X1 port map( D => n7777, CK => CLK, SN => RST, Q 
                           => n7219, QN => n_3835);
   clk_r_REG11126_S15 : DFFS_X1 port map( D => n7219, CK => CLK, SN => RST, Q 
                           => n7218, QN => n_3836);
   clk_r_REG11140_S14 : DFFS_X1 port map( D => n7776, CK => CLK, SN => RST, Q 
                           => n7217, QN => n_3837);
   clk_r_REG11143_S15 : DFFS_X1 port map( D => n7217, CK => CLK, SN => RST, Q 
                           => n7216, QN => n_3838);
   clk_r_REG10976_S14 : DFFR_X1 port map( D => n1443, CK => CLK, RN => RST, Q 
                           => n_3839, QN => n7313);
   clk_r_REG11008_S15 : DFFR_X1 port map( D => n5342, CK => CLK, RN => RST, Q 
                           => n_3840, QN => n7314);
   clk_r_REG11018_S15 : DFFR_X1 port map( D => n5343, CK => CLK, RN => RST, Q 
                           => n_3841, QN => n7315);
   clk_r_REG11025_S15 : DFFR_X1 port map( D => n5344, CK => CLK, RN => RST, Q 
                           => n_3842, QN => n7316);
   clk_r_REG11036_S15 : DFFR_X1 port map( D => n5345, CK => CLK, RN => RST, Q 
                           => n_3843, QN => n7317);
   clk_r_REG11045_S15 : DFFR_X1 port map( D => n5346, CK => CLK, RN => RST, Q 
                           => n_3844, QN => n7309);
   clk_r_REG11053_S15 : DFFR_X1 port map( D => n5347, CK => CLK, RN => RST, Q 
                           => n_3845, QN => n7307);
   clk_r_REG11060_S15 : DFFR_X1 port map( D => n5348, CK => CLK, RN => RST, Q 
                           => n_3846, QN => n7310);
   clk_r_REG11067_S15 : DFFR_X1 port map( D => n5349, CK => CLK, RN => RST, Q 
                           => n_3847, QN => n7318);
   clk_r_REG13297_S4 : DFFR_X1 port map( D => n7346, CK => CLK, RN => RST, Q =>
                           n7205, QN => n_3848);
   clk_r_REG13290_S4 : DFFS_X1 port map( D => n7345, CK => CLK, SN => RST, Q =>
                           n7204, QN => n8071);
   clk_r_REG13294_S4 : DFFR_X1 port map( D => n7359, CK => CLK, RN => RST, Q =>
                           n7203, QN => n_3849);
   clk_r_REG13303_S5 : DFFR_X1 port map( D => n7202, CK => CLK, RN => RST, Q =>
                           n7201, QN => n_3850);
   clk_r_REG13439_S4 : DFFS_X1 port map( D => n7343, CK => CLK, SN => RST, Q =>
                           n7199, QN => n_3851);
   clk_r_REG13423_S2 : DFFS_X1 port map( D => n5405, CK => CLK, SN => RST, Q =>
                           n7198, QN => n_3852);
   clk_r_REG13301_S4 : DFFR_X1 port map( D => n7704, CK => CLK, RN => RST, Q =>
                           n7197, QN => n_3853);
   clk_r_REG11375_S7 : DFFS_X1 port map( D => n7344, CK => CLK, SN => RST, Q =>
                           n7196, QN => n_3854);
   clk_r_REG11792_S6 : DFFR_X1 port map( D => n6207, CK => CLK, RN => RST, Q =>
                           n7195, QN => n_3855);
   clk_r_REG11361_S6 : DFFR_X1 port map( D => n7710, CK => CLK, RN => RST, Q =>
                           n7194, QN => n_3856);
   clk_r_REG13425_S2 : DFFS_X1 port map( D => n5358, CK => CLK, SN => RST, Q =>
                           n7193, QN => n_3857);
   clk_r_REG11064_S5 : DFFR_X1 port map( D => n7729, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_29_port, QN => n_3858);
   clk_r_REG11057_S5 : DFFR_X1 port map( D => n7731, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_27_port, QN => n_3859);
   clk_r_REG11049_S5 : DFFR_X1 port map( D => n7727, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_25_port, QN => n_3860);
   clk_r_REG11040_S5 : DFFR_X1 port map( D => n7725, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_23_port, QN => n_3861);
   clk_r_REG10979_S5 : DFFR_X1 port map( D => n7717, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_15_port, QN => n_3862);
   clk_r_REG11133_S5 : DFFR_X1 port map( D => n7715, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_13_port, QN => n_3863);
   clk_r_REG11012_S5 : DFFR_X1 port map( D => n7723, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_17_port, QN => n_3864);
   clk_r_REG11022_S6 : DFFR_X1 port map( D => n7719, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_19_port, QN => n_3865);
   clk_r_REG11029_S5 : DFFR_X1 port map( D => n7721, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_21_port, QN => n_3866);
   clk_r_REG11147_S5 : DFFR_X1 port map( D => n7713, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_11_port, QN => n_3867);
   clk_r_REG13278_S8 : DFFR_X1 port map( D => n7711, CK => CLK, RN => RST, Q =>
                           n7182, QN => n_3868);
   clk_r_REG13416_S2 : DFFR_X1 port map( D => n7701, CK => CLK, RN => RST, Q =>
                           n7181, QN => n_3869);
   clk_r_REG11354_S6 : DFFR_X1 port map( D => n6113, CK => CLK, RN => RST, Q =>
                           n7180, QN => n_3870);
   clk_r_REG11936_S5 : DFFR_X1 port map( D => n7712, CK => CLK, RN => RST, Q =>
                           n7179, QN => n_3871);
   clk_r_REG13286_S5 : DFFR_X1 port map( D => n7775, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_7_port, QN => n_3872);
   clk_r_REG11154_S5 : DFFR_X1 port map( D => n7774, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_9_port, QN => n_3873);
   clk_r_REG11372_S12 : DFFR_X1 port map( D => n7786, CK => CLK, RN => RST, Q 
                           => IRAM_ADDRESS_5_port, QN => n_3874);
   clk_r_REG13432_S2 : DFFS_X1 port map( D => n7694, CK => CLK, SN => RST, Q =>
                           IRAM_ENABLE, QN => n_3875);
   clk_r_REG11795_S5 : DFFR_X1 port map( D => n7763, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_2_port, QN => n_3876);
   clk_r_REG13437_S3 : DFFR_X1 port map( D => n7361, CK => CLK, RN => RST, Q =>
                           n_3877, QN => n7343);
   clk_r_REG13438_S4 : DFFS_X1 port map( D => n7343, CK => CLK, SN => RST, Q =>
                           n_3878, QN => n7172);
   clk_r_REG11651_S6 : DFFR_X1 port map( D => n6209, CK => CLK, RN => RST, Q =>
                           n7171, QN => n_3879);
   clk_r_REG13635_S1 : DFFR_X1 port map( D => n7347, CK => CLK, RN => RST, Q =>
                           n7170, QN => n_3880);
   clk_r_REG13636_S2 : DFFR_X1 port map( D => n7170, CK => CLK, RN => RST, Q =>
                           n7169, QN => n_3881);
   clk_r_REG13291_S4 : DFFS_X1 port map( D => n7345, CK => CLK, SN => RST, Q =>
                           n7168, QN => n_3882);
   clk_r_REG13288_S3 : DFFR_X1 port map( D => n7333, CK => CLK, RN => RST, Q =>
                           n_3883, QN => n7345);
   clk_r_REG13289_S4 : DFFS_X1 port map( D => n7345, CK => CLK, SN => RST, Q =>
                           n_3884, QN => n7166);
   clk_r_REG11368_S6 : DFFR_X1 port map( D => n6096, CK => CLK, RN => RST, Q =>
                           n7165, QN => n_3885);
   clk_r_REG13378_S1 : DFFR_X1 port map( D => n7342, CK => CLK, RN => RST, Q =>
                           n7164, QN => n_3886);
   clk_r_REG11148_S14 : DFFS_X1 port map( D => n4128, CK => CLK, SN => RST, Q 
                           => n7163, QN => n_3887);
   clk_r_REG11134_S14 : DFFS_X1 port map( D => n7714, CK => CLK, SN => RST, Q 
                           => n7162, QN => n_3888);
   clk_r_REG11122_S15 : DFFS_X1 port map( D => n7716, CK => CLK, SN => RST, Q 
                           => n7161, QN => n_3889);
   clk_r_REG11115_S15 : DFFS_X1 port map( D => n7722, CK => CLK, SN => RST, Q 
                           => n7160, QN => n_3890);
   clk_r_REG11108_S15 : DFFS_X1 port map( D => n7718, CK => CLK, SN => RST, Q 
                           => n7159, QN => n_3891);
   clk_r_REG11102_S15 : DFFS_X1 port map( D => n7720, CK => CLK, SN => RST, Q 
                           => n7158, QN => n_3892);
   clk_r_REG11095_S15 : DFFS_X1 port map( D => n7724, CK => CLK, SN => RST, Q 
                           => n7157, QN => n_3893);
   clk_r_REG11089_S15 : DFFS_X1 port map( D => n7726, CK => CLK, SN => RST, Q 
                           => n7156, QN => n_3894);
   clk_r_REG11083_S15 : DFFS_X1 port map( D => n7730, CK => CLK, SN => RST, Q 
                           => n7155, QN => n_3895);
   clk_r_REG11077_S15 : DFFS_X1 port map( D => n7728, CK => CLK, SN => RST, Q 
                           => n7154, QN => n_3896);
   clk_r_REG13283_S7 : DFFS_X1 port map( D => n7337, CK => CLK, SN => RST, Q =>
                           n7153, QN => n_3897);
   clk_r_REG10960_S14 : DFFS_X1 port map( D => n7336, CK => CLK, SN => RST, Q 
                           => n7152, QN => n_3898);
   clk_r_REG13632_S2 : DFFR_X1 port map( D => n7738, CK => CLK, RN => RST, Q =>
                           n7151, QN => n_3899);
   clk_r_REG13430_S2 : DFFR_X1 port map( D => n7740, CK => CLK, RN => RST, Q =>
                           n7150, QN => n_3900);
   clk_r_REG13292_S3 : DFFS_X1 port map( D => n7702, CK => CLK, SN => RST, Q =>
                           n_3901, QN => n7359);
   clk_r_REG13293_S4 : DFFR_X1 port map( D => n7359, CK => CLK, RN => RST, Q =>
                           n8068, QN => n7148);
   clk_r_REG11080_S16 : DFFR_X1 port map( D => n7358, CK => CLK, RN => RST, Q 
                           => n7147, QN => n_3902);
   clk_r_REG11078_S15 : DFFS_X1 port map( D => n7728, CK => CLK, SN => RST, Q 
                           => n_3903, QN => n7358);
   clk_r_REG11079_S16 : DFFR_X1 port map( D => n7358, CK => CLK, RN => RST, Q 
                           => n_3904, QN => n7145);
   clk_r_REG11086_S16 : DFFR_X1 port map( D => n7357, CK => CLK, RN => RST, Q 
                           => n7144, QN => n_3905);
   clk_r_REG11084_S15 : DFFS_X1 port map( D => n7730, CK => CLK, SN => RST, Q 
                           => n_3906, QN => n7357);
   clk_r_REG11085_S16 : DFFR_X1 port map( D => n7357, CK => CLK, RN => RST, Q 
                           => n_3907, QN => n7142);
   clk_r_REG11092_S16 : DFFR_X1 port map( D => n7356, CK => CLK, RN => RST, Q 
                           => n7141, QN => n_3908);
   clk_r_REG11090_S15 : DFFS_X1 port map( D => n7726, CK => CLK, SN => RST, Q 
                           => n_3909, QN => n7356);
   clk_r_REG11091_S16 : DFFR_X1 port map( D => n7356, CK => CLK, RN => RST, Q 
                           => n_3910, QN => n7139);
   clk_r_REG11098_S16 : DFFR_X1 port map( D => n7355, CK => CLK, RN => RST, Q 
                           => n7138, QN => n_3911);
   clk_r_REG11096_S15 : DFFS_X1 port map( D => n7724, CK => CLK, SN => RST, Q 
                           => n_3912, QN => n7355);
   clk_r_REG11097_S16 : DFFR_X1 port map( D => n7355, CK => CLK, RN => RST, Q 
                           => n_3913, QN => n7136);
   clk_r_REG11105_S16 : DFFR_X1 port map( D => n7354, CK => CLK, RN => RST, Q 
                           => n7135, QN => n_3914);
   clk_r_REG11103_S15 : DFFS_X1 port map( D => n7720, CK => CLK, SN => RST, Q 
                           => n_3915, QN => n7354);
   clk_r_REG11104_S16 : DFFR_X1 port map( D => n7354, CK => CLK, RN => RST, Q 
                           => n_3916, QN => n7133);
   clk_r_REG11111_S16 : DFFR_X1 port map( D => n7353, CK => CLK, RN => RST, Q 
                           => n7132, QN => n_3917);
   clk_r_REG11109_S15 : DFFS_X1 port map( D => n7718, CK => CLK, SN => RST, Q 
                           => n_3918, QN => n7353);
   clk_r_REG11110_S16 : DFFR_X1 port map( D => n7353, CK => CLK, RN => RST, Q 
                           => n_3919, QN => n7130);
   clk_r_REG11118_S16 : DFFR_X1 port map( D => n7352, CK => CLK, RN => RST, Q 
                           => n7129, QN => n_3920);
   clk_r_REG11116_S15 : DFFS_X1 port map( D => n7722, CK => CLK, SN => RST, Q 
                           => n_3921, QN => n7352);
   clk_r_REG11117_S16 : DFFR_X1 port map( D => n7352, CK => CLK, RN => RST, Q 
                           => n_3922, QN => n7127);
   clk_r_REG11125_S16 : DFFR_X1 port map( D => n7351, CK => CLK, RN => RST, Q 
                           => n7126, QN => n_3923);
   clk_r_REG11123_S15 : DFFS_X1 port map( D => n7716, CK => CLK, SN => RST, Q 
                           => n_3924, QN => n7351);
   clk_r_REG11124_S16 : DFFR_X1 port map( D => n7351, CK => CLK, RN => RST, Q 
                           => n_3925, QN => n7124);
   clk_r_REG11137_S15 : DFFR_X1 port map( D => n7350, CK => CLK, RN => RST, Q 
                           => n7123, QN => n_3926);
   clk_r_REG11135_S14 : DFFS_X1 port map( D => n7714, CK => CLK, SN => RST, Q 
                           => n_3927, QN => n7350);
   clk_r_REG11136_S15 : DFFR_X1 port map( D => n7350, CK => CLK, RN => RST, Q 
                           => n_3928, QN => n7121);
   clk_r_REG11151_S15 : DFFR_X1 port map( D => n7338, CK => CLK, RN => RST, Q 
                           => n7120, QN => n_3929);
   clk_r_REG11149_S14 : DFFS_X1 port map( D => n4128, CK => CLK, SN => RST, Q 
                           => n_3930, QN => n7338);
   clk_r_REG11150_S15 : DFFR_X1 port map( D => n7338, CK => CLK, RN => RST, Q 
                           => n_3931, QN => n7118);
   clk_r_REG10963_S15 : DFFR_X1 port map( D => n7349, CK => CLK, RN => RST, Q 
                           => n7117, QN => n_3932);
   clk_r_REG10961_S14 : DFFS_X1 port map( D => n7336, CK => CLK, SN => RST, Q 
                           => n_3933, QN => n7349);
   clk_r_REG10962_S15 : DFFR_X1 port map( D => n7349, CK => CLK, RN => RST, Q 
                           => n_3934, QN => n7115);
   clk_r_REG13285_S8 : DFFR_X1 port map( D => n7360, CK => CLK, RN => RST, Q =>
                           n7114, QN => n_3935);
   clk_r_REG13284_S7 : DFFS_X1 port map( D => n7337, CK => CLK, SN => RST, Q =>
                           n7113, QN => n7360);
   clk_r_REG11376_S7 : DFFS_X1 port map( D => n7344, CK => CLK, SN => RST, Q =>
                           n7112, QN => n_3936);
   clk_r_REG11373_S6 : DFFR_X1 port map( D => n7334, CK => CLK, RN => RST, Q =>
                           n_3937, QN => n7344);
   clk_r_REG11374_S7 : DFFS_X1 port map( D => n7344, CK => CLK, SN => RST, Q =>
                           n_3938, QN => n7110);
   clk_r_REG10316_S4 : DFFR_X1 port map( D => n7348, CK => CLK, RN => RST, Q =>
                           n7109, QN => n_3939);
   clk_r_REG10314_S3 : DFFS_X1 port map( D => n7335, CK => CLK, SN => RST, Q =>
                           n_3940, QN => n7348);
   clk_r_REG13564_S7 : DFFR_X1 port map( D => n7736, CK => CLK, RN => RST, Q =>
                           n7106, QN => n_3941);
   clk_r_REG13295_S3 : DFFS_X1 port map( D => n7702, CK => CLK, SN => RST, Q =>
                           n_3942, QN => n7346);
   clk_r_REG13296_S4 : DFFR_X1 port map( D => n7346, CK => CLK, RN => RST, Q =>
                           n_3943, QN => n7104);
   clk_r_REG13298_S4 : DFFR_X1 port map( D => n7346, CK => CLK, RN => RST, Q =>
                           n7103, QN => n_3944);
   clk_r_REG13536_S2 : DFFS_X1 port map( D => n6178, CK => CLK, SN => RST, Q =>
                           n_3945, QN => n8075);
   clk_r_REG13426_S2 : DFFR_X1 port map( D => n7706, CK => CLK, RN => RST, Q =>
                           DRAM_ENABLE, QN => n_3946);
   clk_r_REG13566_S7 : DFFS_X1 port map( D => n7751, CK => CLK, SN => RST, Q =>
                           n7100, QN => n8069);
   clk_r_REG13568_S7 : DFFS_X1 port map( D => n7750, CK => CLK, SN => RST, Q =>
                           n7099, QN => n8070);
   clk_r_REG13570_S7 : DFFS_X1 port map( D => n7749, CK => CLK, SN => RST, Q =>
                           n7098, QN => n8074);
   clk_r_REG13572_S7 : DFFS_X1 port map( D => n7748, CK => CLK, SN => RST, Q =>
                           n7097, QN => n8073);
   clk_r_REG13480_S6 : DFFS_X1 port map( D => n7703, CK => CLK, SN => RST, Q =>
                           n7096, QN => n_3947);
   clk_r_REG13573_S6 : DFFS_X1 port map( D => n7709, CK => CLK, SN => RST, Q =>
                           n7095, QN => n_3948);
   clk_r_REG10374_S3 : DFFR_X1 port map( D => n7094, CK => CLK, RN => RST, Q =>
                           n7093, QN => n_3949);
   clk_r_REG10385_S2 : DFF_X1 port map( D => n1671, CK => CLK, Q => n7092, QN 
                           => n_3950);
   clk_r_REG10386_S3 : DFFR_X1 port map( D => n7092, CK => CLK, RN => RST, Q =>
                           n7091, QN => n_3951);
   clk_r_REG13019_S2 : DFF_X1 port map( D => n1669, CK => CLK, Q => n7090, QN 
                           => n_3952);
   clk_r_REG13020_S3 : DFFR_X1 port map( D => n7090, CK => CLK, RN => RST, Q =>
                           n7089, QN => n_3953);
   clk_r_REG10477_S2 : DFF_X1 port map( D => n1667, CK => CLK, Q => n7088, QN 
                           => n_3954);
   clk_r_REG10478_S3 : DFFR_X1 port map( D => n7088, CK => CLK, RN => RST, Q =>
                           n7087, QN => n_3955);
   clk_r_REG12384_S2 : DFF_X1 port map( D => n1665, CK => CLK, Q => n7086, QN 
                           => n_3956);
   clk_r_REG12385_S3 : DFFR_X1 port map( D => n7086, CK => CLK, RN => RST, Q =>
                           n7085, QN => n_3957);
   clk_r_REG12448_S2 : DFF_X1 port map( D => n1663, CK => CLK, Q => n7084, QN 
                           => n_3958);
   clk_r_REG12449_S3 : DFFR_X1 port map( D => n7084, CK => CLK, RN => RST, Q =>
                           n7083, QN => n_3959);
   clk_r_REG12512_S2 : DFF_X1 port map( D => n1661, CK => CLK, Q => n7082, QN 
                           => n_3960);
   clk_r_REG12513_S3 : DFFR_X1 port map( D => n7082, CK => CLK, RN => RST, Q =>
                           n7081, QN => n_3961);
   clk_r_REG12576_S2 : DFF_X1 port map( D => n1659, CK => CLK, Q => n7080, QN 
                           => n_3962);
   clk_r_REG12577_S3 : DFFR_X1 port map( D => n7080, CK => CLK, RN => RST, Q =>
                           n7079, QN => n_3963);
   clk_r_REG10410_S2 : DFF_X1 port map( D => n1657, CK => CLK, Q => n7078, QN 
                           => n_3964);
   clk_r_REG10411_S3 : DFFR_X1 port map( D => n7078, CK => CLK, RN => RST, Q =>
                           n7077, QN => n_3965);
   clk_r_REG12767_S2 : DFF_X1 port map( D => n1655, CK => CLK, Q => n7076, QN 
                           => n_3966);
   clk_r_REG12768_S3 : DFFR_X1 port map( D => n7076, CK => CLK, RN => RST, Q =>
                           n7075, QN => n_3967);
   clk_r_REG12831_S2 : DFF_X1 port map( D => n1653, CK => CLK, Q => n7074, QN 
                           => n_3968);
   clk_r_REG12832_S3 : DFFR_X1 port map( D => n7074, CK => CLK, RN => RST, Q =>
                           n7073, QN => n_3969);
   clk_r_REG10495_S2 : DFF_X1 port map( D => n1651, CK => CLK, Q => n7072, QN 
                           => n_3970);
   clk_r_REG10496_S3 : DFFR_X1 port map( D => n7072, CK => CLK, RN => RST, Q =>
                           n7071, QN => n_3971);
   clk_r_REG10310_S2 : DFF_X1 port map( D => n1649, CK => CLK, Q => n7070, QN 
                           => n_3972);
   clk_r_REG13305_S3 : DFFR_X1 port map( D => n7070, CK => CLK, RN => RST, Q =>
                           n7069, QN => n_3973);
   clk_r_REG12258_S2 : DFF_X1 port map( D => n1647, CK => CLK, Q => n7068, QN 
                           => n_3974);
   clk_r_REG12259_S3 : DFFR_X1 port map( D => n7068, CK => CLK, RN => RST, Q =>
                           n7067, QN => n_3975);
   clk_r_REG13083_S2 : DFF_X1 port map( D => n1645, CK => CLK, Q => n7066, QN 
                           => n_3976);
   clk_r_REG13084_S3 : DFFR_X1 port map( D => n7066, CK => CLK, RN => RST, Q =>
                           n7065, QN => n_3977);
   clk_r_REG13147_S2 : DFF_X1 port map( D => n1643, CK => CLK, Q => n7064, QN 
                           => n_3978);
   clk_r_REG13148_S3 : DFFR_X1 port map( D => n7064, CK => CLK, RN => RST, Q =>
                           n7063, QN => n_3979);
   clk_r_REG12003_S2 : DFF_X1 port map( D => n1641, CK => CLK, Q => n7062, QN 
                           => n_3980);
   clk_r_REG12004_S3 : DFFR_X1 port map( D => n7062, CK => CLK, RN => RST, Q =>
                           n7061, QN => n_3981);
   clk_r_REG10647_S2 : DFF_X1 port map( D => n1639, CK => CLK, Q => n7060, QN 
                           => n_3982);
   clk_r_REG10648_S3 : DFFR_X1 port map( D => n7060, CK => CLK, RN => RST, Q =>
                           n7059, QN => n_3983);
   clk_r_REG12067_S2 : DFF_X1 port map( D => n1637, CK => CLK, Q => n7058, QN 
                           => n_3984);
   clk_r_REG12068_S3 : DFFR_X1 port map( D => n7058, CK => CLK, RN => RST, Q =>
                           n7057, QN => n_3985);
   clk_r_REG12131_S2 : DFF_X1 port map( D => n1635, CK => CLK, Q => n7056, QN 
                           => n_3986);
   clk_r_REG12132_S3 : DFFR_X1 port map( D => n7056, CK => CLK, RN => RST, Q =>
                           n7055, QN => n_3987);
   clk_r_REG10741_S2 : DFF_X1 port map( D => n1633, CK => CLK, Q => n7054, QN 
                           => n_3988);
   clk_r_REG10742_S3 : DFFR_X1 port map( D => n7054, CK => CLK, RN => RST, Q =>
                           n7053, QN => n_3989);
   clk_r_REG10782_S2 : DFF_X1 port map( D => n1631, CK => CLK, Q => n7052, QN 
                           => n_3990);
   clk_r_REG10783_S3 : DFFR_X1 port map( D => n7052, CK => CLK, RN => RST, Q =>
                           n7051, QN => n_3991);
   clk_r_REG10849_S2 : DFF_X1 port map( D => n1629, CK => CLK, Q => n7050, QN 
                           => n_3992);
   clk_r_REG10886_S2 : DFF_X1 port map( D => n1627, CK => CLK, Q => n7049, QN 
                           => n_3993);
   clk_r_REG11444_S2 : DFF_X1 port map( D => n1625, CK => CLK, Q => n7048, QN 
                           => n_3994);
   clk_r_REG12641_S2 : DFF_X1 port map( D => n1623, CK => CLK, Q => n7047, QN 
                           => n_3995);
   clk_r_REG11507_S2 : DFF_X1 port map( D => n1621, CK => CLK, Q => n7046, QN 
                           => n_3996);
   clk_r_REG11276_S2 : DFF_X1 port map( D => n1619, CK => CLK, Q => n7045, QN 
                           => n_3997);
   clk_r_REG11581_S2 : DFF_X1 port map( D => n1617, CK => CLK, Q => n7044, QN 
                           => n_3998);
   clk_r_REG11723_S2 : DFF_X1 port map( D => n1615, CK => CLK, Q => n7043, QN 
                           => n_3999);
   clk_r_REG11866_S2 : DFF_X1 port map( D => n1614, CK => CLK, Q => n7042, QN 
                           => n_4000);
   clk_r_REG13211_S2 : DFF_X1 port map( D => n1613, CK => CLK, Q => n7041, QN 
                           => n_4001);
   clk_r_REG10369_S2 : DFF_X1 port map( D => n5229, CK => CLK, Q => n7040, QN 
                           => n_4002);
   clk_r_REG10370_S3 : DFFR_X1 port map( D => n7040, CK => CLK, RN => RST, Q =>
                           n7039, QN => n_4003);
   clk_r_REG10371_S4 : DFFR_X1 port map( D => n7039, CK => CLK, RN => RST, Q =>
                           n7038, QN => n_4004);
   clk_r_REG10379_S2 : DFF_X1 port map( D => n5226, CK => CLK, Q => n7037, QN 
                           => n_4005);
   clk_r_REG10380_S3 : DFFR_X1 port map( D => n7037, CK => CLK, RN => RST, Q =>
                           n7036, QN => n_4006);
   clk_r_REG10381_S4 : DFFR_X1 port map( D => n7036, CK => CLK, RN => RST, Q =>
                           n7035, QN => n_4007);
   clk_r_REG10360_S2 : DFF_X1 port map( D => n5223, CK => CLK, Q => n7034, QN 
                           => n_4008);
   clk_r_REG10361_S3 : DFFR_X1 port map( D => n7034, CK => CLK, RN => RST, Q =>
                           n7033, QN => n_4009);
   clk_r_REG10362_S4 : DFFR_X1 port map( D => n7033, CK => CLK, RN => RST, Q =>
                           n7032, QN => n_4010);
   clk_r_REG10472_S2 : DFF_X1 port map( D => n5220, CK => CLK, Q => n7031, QN 
                           => n_4011);
   clk_r_REG10473_S3 : DFFR_X1 port map( D => n7031, CK => CLK, RN => RST, Q =>
                           n7030, QN => n_4012);
   clk_r_REG10474_S4 : DFFR_X1 port map( D => n7030, CK => CLK, RN => RST, Q =>
                           n7029, QN => n_4013);
   clk_r_REG10465_S2 : DFF_X1 port map( D => n5217, CK => CLK, Q => n7028, QN 
                           => n_4014);
   clk_r_REG10466_S3 : DFFR_X1 port map( D => n7028, CK => CLK, RN => RST, Q =>
                           n7027, QN => n_4015);
   clk_r_REG10467_S4 : DFFR_X1 port map( D => n7027, CK => CLK, RN => RST, Q =>
                           n7026, QN => n_4016);
   clk_r_REG10458_S2 : DFF_X1 port map( D => n5214, CK => CLK, Q => n7025, QN 
                           => n_4017);
   clk_r_REG10459_S3 : DFFR_X1 port map( D => n7025, CK => CLK, RN => RST, Q =>
                           n7024, QN => n_4018);
   clk_r_REG10460_S4 : DFFR_X1 port map( D => n7024, CK => CLK, RN => RST, Q =>
                           n7023, QN => n_4019);
   clk_r_REG10451_S2 : DFF_X1 port map( D => n5211, CK => CLK, Q => n7022, QN 
                           => n_4020);
   clk_r_REG10452_S3 : DFFR_X1 port map( D => n7022, CK => CLK, RN => RST, Q =>
                           n7021, QN => n_4021);
   clk_r_REG10453_S4 : DFFR_X1 port map( D => n7021, CK => CLK, RN => RST, Q =>
                           n7020, QN => n_4022);
   clk_r_REG10442_S2 : DFF_X1 port map( D => n5208, CK => CLK, Q => n7019, QN 
                           => n_4023);
   clk_r_REG10443_S3 : DFFR_X1 port map( D => n7019, CK => CLK, RN => RST, Q =>
                           n7018, QN => n_4024);
   clk_r_REG10444_S4 : DFFR_X1 port map( D => n7018, CK => CLK, RN => RST, Q =>
                           n7017, QN => n_4025);
   clk_r_REG10406_S2 : DFF_X1 port map( D => n5205, CK => CLK, Q => n7016, QN 
                           => n_4026);
   clk_r_REG10407_S3 : DFFR_X1 port map( D => n7016, CK => CLK, RN => RST, Q =>
                           n7015, QN => n_4027);
   clk_r_REG10408_S4 : DFFR_X1 port map( D => n7015, CK => CLK, RN => RST, Q =>
                           n7014, QN => n_4028);
   clk_r_REG10399_S2 : DFF_X1 port map( D => n5202, CK => CLK, Q => n7013, QN 
                           => n_4029);
   clk_r_REG10400_S3 : DFFR_X1 port map( D => n7013, CK => CLK, RN => RST, Q =>
                           n7012, QN => n_4030);
   clk_r_REG10401_S4 : DFFR_X1 port map( D => n7012, CK => CLK, RN => RST, Q =>
                           n7011, QN => n_4031);
   clk_r_REG10392_S2 : DFF_X1 port map( D => n5199, CK => CLK, Q => n7010, QN 
                           => n_4032);
   clk_r_REG10393_S3 : DFFR_X1 port map( D => n7010, CK => CLK, RN => RST, Q =>
                           n7009, QN => n_4033);
   clk_r_REG10394_S4 : DFFR_X1 port map( D => n7009, CK => CLK, RN => RST, Q =>
                           n7008, QN => n_4034);
   clk_r_REG10490_S2 : DFF_X1 port map( D => n5196, CK => CLK, Q => n7007, QN 
                           => n_4035);
   clk_r_REG10491_S3 : DFFR_X1 port map( D => n7007, CK => CLK, RN => RST, Q =>
                           n7006, QN => n_4036);
   clk_r_REG10492_S4 : DFFR_X1 port map( D => n7006, CK => CLK, RN => RST, Q =>
                           n7005, QN => n_4037);
   clk_r_REG10303_S2 : DFF_X1 port map( D => n5193, CK => CLK, Q => n7004, QN 
                           => n_4038);
   clk_r_REG10304_S3 : DFFR_X1 port map( D => n7004, CK => CLK, RN => RST, Q =>
                           n7003, QN => n_4039);
   clk_r_REG10305_S4 : DFFR_X1 port map( D => n7003, CK => CLK, RN => RST, Q =>
                           n7002, QN => n_4040);
   clk_r_REG10483_S2 : DFF_X1 port map( D => n5190, CK => CLK, Q => n7001, QN 
                           => n_4041);
   clk_r_REG10484_S3 : DFFR_X1 port map( D => n7001, CK => CLK, RN => RST, Q =>
                           n7000, QN => n_4042);
   clk_r_REG10485_S4 : DFFR_X1 port map( D => n7000, CK => CLK, RN => RST, Q =>
                           n6999, QN => n_4043);
   clk_r_REG10352_S2 : DFF_X1 port map( D => n5187, CK => CLK, Q => n6998, QN 
                           => n_4044);
   clk_r_REG10353_S3 : DFFR_X1 port map( D => n6998, CK => CLK, RN => RST, Q =>
                           n6997, QN => n_4045);
   clk_r_REG10354_S4 : DFFR_X1 port map( D => n6997, CK => CLK, RN => RST, Q =>
                           n6996, QN => n_4046);
   clk_r_REG10345_S2 : DFF_X1 port map( D => n5184, CK => CLK, Q => n6995, QN 
                           => n_4047);
   clk_r_REG10346_S3 : DFFR_X1 port map( D => n6995, CK => CLK, RN => RST, Q =>
                           n6994, QN => n_4048);
   clk_r_REG10347_S4 : DFFR_X1 port map( D => n6994, CK => CLK, RN => RST, Q =>
                           n6993, QN => n_4049);
   clk_r_REG10621_S2 : DFF_X1 port map( D => n5181, CK => CLK, Q => n6992, QN 
                           => n_4050);
   clk_r_REG10622_S3 : DFFR_X1 port map( D => n6992, CK => CLK, RN => RST, Q =>
                           n6991, QN => n_4051);
   clk_r_REG10623_S4 : DFFR_X1 port map( D => n6991, CK => CLK, RN => RST, Q =>
                           n6990, QN => n_4052);
   clk_r_REG10637_S2 : DFF_X1 port map( D => n5178, CK => CLK, Q => n6989, QN 
                           => n_4053);
   clk_r_REG10638_S3 : DFFR_X1 port map( D => n6989, CK => CLK, RN => RST, Q =>
                           n6988, QN => n_4054);
   clk_r_REG10639_S4 : DFFR_X1 port map( D => n6988, CK => CLK, RN => RST, Q =>
                           n6987, QN => n_4055);
   clk_r_REG10543_S2 : DFF_X1 port map( D => n5175, CK => CLK, Q => n6986, QN 
                           => n_4056);
   clk_r_REG10544_S3 : DFFR_X1 port map( D => n6986, CK => CLK, RN => RST, Q =>
                           n6985, QN => n_4057);
   clk_r_REG10545_S4 : DFFR_X1 port map( D => n6985, CK => CLK, RN => RST, Q =>
                           n6984, QN => n_4058);
   clk_r_REG10524_S2 : DFF_X1 port map( D => n5172, CK => CLK, Q => n6983, QN 
                           => n_4059);
   clk_r_REG10525_S3 : DFFR_X1 port map( D => n6983, CK => CLK, RN => RST, Q =>
                           n6982, QN => n_4060);
   clk_r_REG10526_S4 : DFFR_X1 port map( D => n6982, CK => CLK, RN => RST, Q =>
                           n6981, QN => n_4061);
   clk_r_REG10713_S2 : DFF_X1 port map( D => n5169, CK => CLK, Q => n6980, QN 
                           => n_4062);
   clk_r_REG10714_S3 : DFFR_X1 port map( D => n6980, CK => CLK, RN => RST, Q =>
                           n6979, QN => n_4063);
   clk_r_REG10715_S4 : DFFR_X1 port map( D => n6979, CK => CLK, RN => RST, Q =>
                           n6978, QN => n_4064);
   clk_r_REG10778_S2 : DFF_X1 port map( D => n5166, CK => CLK, Q => n6977, QN 
                           => n_4065);
   clk_r_REG10779_S3 : DFFR_X1 port map( D => n6977, CK => CLK, RN => RST, Q =>
                           n6976, QN => n_4066);
   clk_r_REG10780_S4 : DFFR_X1 port map( D => n6976, CK => CLK, RN => RST, Q =>
                           n6975, QN => n_4067);
   clk_r_REG10841_S2 : DFF_X1 port map( D => n5163, CK => CLK, Q => n6974, QN 
                           => n_4068);
   clk_r_REG10842_S3 : DFFR_X1 port map( D => n6974, CK => CLK, RN => RST, Q =>
                           n6973, QN => n_4069);
   clk_r_REG10843_S4 : DFFR_X1 port map( D => n6973, CK => CLK, RN => RST, Q =>
                           n6972, QN => n_4070);
   clk_r_REG10880_S2 : DFF_X1 port map( D => n5160, CK => CLK, Q => n6971, QN 
                           => n_4071);
   clk_r_REG10881_S3 : DFFR_X1 port map( D => n6971, CK => CLK, RN => RST, Q =>
                           n6970, QN => n_4072);
   clk_r_REG10882_S4 : DFFR_X1 port map( D => n6970, CK => CLK, RN => RST, Q =>
                           n6969, QN => n_4073);
   clk_r_REG10827_S2 : DFF_X1 port map( D => n5157, CK => CLK, Q => n6968, QN 
                           => n_4074);
   clk_r_REG10828_S3 : DFFR_X1 port map( D => n6968, CK => CLK, RN => RST, Q =>
                           n6967, QN => n_4075);
   clk_r_REG10829_S4 : DFFR_X1 port map( D => n6967, CK => CLK, RN => RST, Q =>
                           n6966, QN => n_4076);
   clk_r_REG10418_S2 : DFF_X1 port map( D => n5154, CK => CLK, Q => n6965, QN 
                           => n_4077);
   clk_r_REG10419_S3 : DFFR_X1 port map( D => n6965, CK => CLK, RN => RST, Q =>
                           n6964, QN => n_4078);
   clk_r_REG10420_S4 : DFFR_X1 port map( D => n6964, CK => CLK, RN => RST, Q =>
                           n6963, QN => n_4079);
   clk_r_REG10808_S2 : DFF_X1 port map( D => n5151, CK => CLK, Q => n6962, QN 
                           => n_4080);
   clk_r_REG10809_S3 : DFFR_X1 port map( D => n6962, CK => CLK, RN => RST, Q =>
                           n6961, QN => n_4081);
   clk_r_REG10810_S4 : DFFR_X1 port map( D => n6961, CK => CLK, RN => RST, Q =>
                           n6960, QN => n_4082);
   clk_r_REG10867_S2 : DFF_X1 port map( D => n5148, CK => CLK, Q => n6959, QN 
                           => n_4083);
   clk_r_REG10868_S3 : DFFR_X1 port map( D => n6959, CK => CLK, RN => RST, Q =>
                           n6958, QN => n_4084);
   clk_r_REG10869_S4 : DFFR_X1 port map( D => n6958, CK => CLK, RN => RST, Q =>
                           n6957, QN => n_4085);
   clk_r_REG10794_S2 : DFF_X1 port map( D => n5145, CK => CLK, Q => n6956, QN 
                           => n_4086);
   clk_r_REG10795_S3 : DFFR_X1 port map( D => n6956, CK => CLK, RN => RST, Q =>
                           n6955, QN => n_4087);
   clk_r_REG10796_S4 : DFFR_X1 port map( D => n6955, CK => CLK, RN => RST, Q =>
                           n6954, QN => n_4088);
   clk_r_REG10765_S2 : DFF_X1 port map( D => n5142, CK => CLK, Q => n6953, QN 
                           => n_4089);
   clk_r_REG10766_S3 : DFFR_X1 port map( D => n6953, CK => CLK, RN => RST, Q =>
                           n6952, QN => n_4090);
   clk_r_REG10767_S4 : DFFR_X1 port map( D => n6952, CK => CLK, RN => RST, Q =>
                           n6951, QN => n_4091);
   clk_r_REG10697_S2 : DFF_X1 port map( D => n5139, CK => CLK, Q => n6950, QN 
                           => n_4092);
   clk_r_REG10698_S3 : DFFR_X1 port map( D => n6950, CK => CLK, RN => RST, Q =>
                           n6949, QN => n_4093);
   clk_r_REG10699_S4 : DFFR_X1 port map( D => n6949, CK => CLK, RN => RST, Q =>
                           n6948, QN => n_4094);
   clk_r_REG10324_S2 : DFF_X1 port map( D => n5136, CK => CLK, Q => n6947, QN 
                           => n_4095);
   clk_r_REG10325_S3 : DFFR_X1 port map( D => n6947, CK => CLK, RN => RST, Q =>
                           n6946, QN => n_4096);
   clk_r_REG10326_S4 : DFFR_X1 port map( D => n6946, CK => CLK, RN => RST, Q =>
                           n6945, QN => n_4097);
   clk_r_REG13628_S4 : DFFR_X1 port map( D => n3284, CK => CLK, RN => RST, Q =>
                           n_4098, QN => n7364);
   clk_r_REG13630_S4 : DFFR_X1 port map( D => n4417, CK => CLK, RN => RST, Q =>
                           n_4099, QN => n7365);
   clk_r_REG13434_S4 : DFFR_X1 port map( D => n5131, CK => CLK, RN => RST, Q =>
                           n6942, QN => n8077);
   clk_r_REG13373_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port, CK 
                           => CLK, RN => RST, Q => n6941, QN => n_4100);
   clk_r_REG13371_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port, CK 
                           => CLK, RN => RST, Q => n6940, QN => n_4101);
   clk_r_REG13368_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port, CK 
                           => CLK, RN => RST, Q => n6939, QN => n_4102);
   clk_r_REG13486_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port, CK 
                           => CLK, RN => RST, Q => n6938, QN => n_4103);
   clk_r_REG13427_S2 : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => CLK, 
                           RN => RST, Q => n6936, QN => n_4104);
   clk_r_REG13422_S2 : DFFR_X1 port map( D => n7705, CK => CLK, RN => RST, Q =>
                           n_4105, QN => n6935);
   clk_r_REG13561_S7 : DFFR_X1 port map( D => n7739, CK => CLK, RN => RST, Q =>
                           n_4106, QN => n6934);
   clk_r_REG13414_S1 : DFFR_X1 port map( D => n5122, CK => CLK, RN => RST, Q =>
                           n6933, QN => n_4107);
   clk_r_REG13563_S7 : DFFR_X1 port map( D => n5089, CK => CLK, RN => RST, Q =>
                           n6932, QN => n_4108);
   clk_r_REG13629_S4 : DFFS_X1 port map( D => n7362, CK => CLK, SN => RST, Q =>
                           n_4109, QN => n6931);
   clk_r_REG13559_S7 : DFFS_X1 port map( D => n474, CK => CLK, SN => RST, Q => 
                           n_4110, QN => n7339);
   clk_r_REG13532_S2 : DFFS_X1 port map( D => n7743, CK => CLK, SN => RST, Q =>
                           n_4111, QN => n6929);
   clk_r_REG13433_S2 : DFFS_X1 port map( D => n5117, CK => CLK, SN => RST, Q =>
                           n6928, QN => n_4112);
   clk_r_REG13483_S7 : DFFS_X1 port map( D => n477, CK => CLK, SN => RST, Q => 
                           n6927, QN => n_4113);
   clk_r_REG13531_S2 : DFFR_X1 port map( D => cu_i_n135, CK => CLK, RN => RST, 
                           Q => n6926, QN => n_4114);
   clk_r_REG11152_S14 : DFFS_X1 port map( D => n6082, CK => CLK, SN => RST, Q 
                           => n6925, QN => n_4115);
   clk_r_REG10965_S13 : DFFR_X1 port map( D => n7341, CK => CLK, RN => RST, Q 
                           => n_4116, QN => n6924);
   clk_r_REG13634_S1 : DFFR_X1 port map( D => n7347, CK => CLK, RN => RST, Q =>
                           n_4117, QN => n6923);
   clk_r_REG10318_S6 : DFFR_X1 port map( D => n5507, CK => CLK, RN => RST, Q =>
                           n6922, QN => n7337);
   clk_r_REG10959_S13 : DFFR_X1 port map( D => n5506, CK => CLK, RN => RST, Q 
                           => n6921, QN => n7336);
   clk_r_REG13476_S6 : DFFS_X1 port map( D => n5098, CK => CLK, SN => RST, Q =>
                           n6920, QN => n_4118);
   clk_r_REG13475_S6 : DFFR_X1 port map( D => n5097, CK => CLK, RN => RST, Q =>
                           n6919, QN => n_4119);
   clk_r_REG11146_S5 : DFFR_X1 port map( D => n6081, CK => CLK, RN => RST, Q =>
                           n6918, QN => n_4120);
   clk_r_REG11142_S14 : DFFS_X1 port map( D => n4231, CK => CLK, SN => RST, Q 
                           => n6917, QN => n_4121);
   clk_r_REG11132_S5 : DFFR_X1 port map( D => n5120, CK => CLK, RN => RST, Q =>
                           n6916, QN => n_4122);
   clk_r_REG13287_S3 : DFFR_X1 port map( D => n7333, CK => CLK, RN => RST, Q =>
                           n_4123, QN => n6915);
   clk_r_REG13633_S1 : DFFS_X1 port map( D => n5092, CK => CLK, SN => RST, Q =>
                           n6914, QN => n_4124);
   clk_r_REG10969_S12 : DFFR_X1 port map( D => n6157, CK => CLK, RN => RST, Q 
                           => n6913, QN => n_4125);
   clk_r_REG10971_S12 : DFFR_X1 port map( D => n6159, CK => CLK, RN => RST, Q 
                           => n6912, QN => n_4126);
   clk_r_REG10970_S12 : DFFS_X1 port map( D => n6159, CK => CLK, SN => RST, Q 
                           => n6911, QN => n_4127);
   clk_r_REG10972_S12 : DFFS_X1 port map( D => n4341, CK => CLK, SN => RST, Q 
                           => n6910, QN => n_4128);
   clk_r_REG13484_S7 : DFFS_X1 port map( D => n492, CK => CLK, SN => RST, Q => 
                           n6909, QN => n_4129);
   clk_r_REG11072_S16 : DFFS_X1 port map( D => n5085, CK => CLK, SN => RST, Q 
                           => n6908, QN => n_4130);
   clk_r_REG10311_S2 : DFF_X1 port map( D => n5084, CK => CLK, Q => n6907, QN 
                           => n_4131);
   clk_r_REG13436_S2 : DFFS_X1 port map( D => n3596, CK => CLK, SN => RST, Q =>
                           n_4132, QN => n7361);
   clk_r_REG13367_S1 : DFFS_X1 port map( D => n2299, CK => CLK, SN => RST, Q =>
                           n_4133, QN => n7367);
   clk_r_REG10313_S3 : DFFS_X1 port map( D => n7335, CK => CLK, SN => RST, Q =>
                           n_4134, QN => n6904);
   clk_r_REG13377_S1 : DFFR_X1 port map( D => n7342, CK => CLK, RN => RST, Q =>
                           n8067, QN => n6903);
   clk_r_REG13601_S7 : DFFR_X1 port map( D => n5047, CK => CLK, RN => RST, Q =>
                           n6902, QN => n_4135);
   clk_r_REG13567_S7 : DFFS_X1 port map( D => n7750, CK => CLK, SN => RST, Q =>
                           n_4136, QN => n6901);
   clk_r_REG13482_S7 : DFFR_X1 port map( D => n5076, CK => CLK, RN => RST, Q =>
                           n6900, QN => n8078);
   clk_r_REG13569_S7 : DFFS_X1 port map( D => n7749, CK => CLK, SN => RST, Q =>
                           n_4137, QN => n6899);
   clk_r_REG13487_S7 : DFFR_X1 port map( D => n5077, CK => CLK, RN => RST, Q =>
                           n6898, QN => n_4138);
   clk_r_REG13571_S7 : DFFS_X1 port map( D => n7748, CK => CLK, SN => RST, Q =>
                           n_4139, QN => n6897);
   clk_r_REG13554_S7 : DFFR_X1 port map( D => n5075, CK => CLK, RN => RST, Q =>
                           n6896, QN => n_4140);
   clk_r_REG13616_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_16_port,
                           CK => CLK, RN => RST, Q => n6895, QN => n_4141);
   clk_r_REG13435_S4 : DFFS_X1 port map( D => n5073, CK => CLK, SN => RST, Q =>
                           n6894, QN => n_4142);
   clk_r_REG13617_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_17_port,
                           CK => CLK, RN => RST, Q => n6893, QN => n_4143);
   clk_r_REG13618_S7 : DFFR_X1 port map( D => n5065, CK => CLK, RN => RST, Q =>
                           n6892, QN => n_4144);
   clk_r_REG13619_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_19_port,
                           CK => CLK, RN => RST, Q => n6891, QN => n_4145);
   clk_r_REG13622_S7 : DFFR_X1 port map( D => n5067, CK => CLK, RN => RST, Q =>
                           n6890, QN => n_4146);
   clk_r_REG13489_S7 : DFFR_X1 port map( D => n5071, CK => CLK, RN => RST, Q =>
                           n6889, QN => n_4147);
   clk_r_REG13623_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_20_port,
                           CK => CLK, RN => RST, Q => n6888, QN => n_4148);
   clk_r_REG11648_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_4149);
   clk_r_REG11351_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_4150);
   clk_r_REG11369_S5 : DFFR_X1 port map( D => n1453, CK => CLK, RN => RST, Q =>
                           IRAM_ADDRESS_6_port, QN => n_4151);
   clk_r_REG13530_S2 : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK => CLK, 
                           RN => RST, Q => n6883, QN => n_4152);
   clk_r_REG13376_S1 : DFFR_X1 port map( D => n4052, CK => CLK, RN => RST, Q =>
                           n6882, QN => n_4153);
   clk_r_REG13626_S7 : DFFR_X1 port map( D => n5079, CK => CLK, RN => RST, Q =>
                           n6881, QN => n_4154);
   clk_r_REG13479_S6 : DFFS_X1 port map( D => n7703, CK => CLK, SN => RST, Q =>
                           n_4155, QN => n6880);
   clk_r_REG13429_S3 : DFFR_X1 port map( D => n5053, CK => CLK, RN => RST, Q =>
                           n6879, QN => n_4156);
   clk_r_REG13431_S3 : DFFR_X1 port map( D => n5052, CK => CLK, RN => RST, Q =>
                           n6878, QN => n_4157);
   clk_r_REG13418_S2 : DFFR_X1 port map( D => n5051, CK => CLK, RN => RST, Q =>
                           n6877, QN => n_4158);
   clk_r_REG13491_S7 : DFFR_X1 port map( D => n5049, CK => CLK, RN => RST, Q =>
                           n6876, QN => n_4159);
   clk_r_REG13516_S7 : DFFR_X1 port map( D => n5048, CK => CLK, RN => RST, Q =>
                           n6875, QN => n_4160);
   clk_r_REG13627_S7 : DFFR_X1 port map( D => n5046, CK => CLK, RN => RST, Q =>
                           n6874, QN => n_4161);
   clk_r_REG13520_S7 : DFFR_X1 port map( D => n5045, CK => CLK, RN => RST, Q =>
                           n6873, QN => n_4162);
   clk_r_REG13522_S7 : DFFR_X1 port map( D => n5044, CK => CLK, RN => RST, Q =>
                           n6872, QN => n_4163);
   clk_r_REG13524_S7 : DFFR_X1 port map( D => n5043, CK => CLK, RN => RST, Q =>
                           n6871, QN => n_4164);
   clk_r_REG13526_S7 : DFFR_X1 port map( D => n5042, CK => CLK, RN => RST, Q =>
                           n6870, QN => n_4165);
   clk_r_REG13528_S7 : DFFR_X1 port map( D => n5041, CK => CLK, RN => RST, Q =>
                           n6869, QN => n_4166);
   clk_r_REG13527_S9 : DFFR_X1 port map( D => n5040, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6868, QN => n_4167);
   clk_r_REG13525_S9 : DFFR_X1 port map( D => n5039, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6867, QN => n_4168);
   clk_r_REG13523_S9 : DFFR_X1 port map( D => n5038, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6866, QN => n_4169);
   clk_r_REG13521_S9 : DFFR_X1 port map( D => n5037, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6865, QN => n_4170);
   clk_r_REG13490_S9 : DFFR_X1 port map( D => n5036, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6864, QN => n_4171);
   clk_r_REG13538_S3 : DFFR_X1 port map( D => n5035, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6863, QN => n_4172);
   clk_r_REG13539_S3 : DFFR_X1 port map( D => n5034, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6862, QN => n_4173);
   clk_r_REG13540_S3 : DFFR_X1 port map( D => n5033, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6861, QN => n_4174);
   clk_r_REG13541_S3 : DFFR_X1 port map( D => n5032, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6860, QN => n_4175);
   clk_r_REG13542_S3 : DFFR_X1 port map( D => n5031, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6859, QN => n_4176);
   clk_r_REG13543_S3 : DFFR_X1 port map( D => n5030, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6858, QN => n_4177);
   clk_r_REG13544_S3 : DFFR_X1 port map( D => n5029, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6857, QN => n_4178);
   clk_r_REG13545_S3 : DFFR_X1 port map( D => n5028, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6856, QN => n_4179);
   clk_r_REG13546_S3 : DFFR_X1 port map( D => n5027, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6855, QN => n_4180);
   clk_r_REG13547_S3 : DFFR_X1 port map( D => n5026, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6854, QN => n_4181);
   clk_r_REG13548_S3 : DFFR_X1 port map( D => n5025, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6853, QN => n_4182);
   clk_r_REG13549_S3 : DFFR_X1 port map( D => n5024, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6852, QN => n_4183);
   clk_r_REG13517_S9 : DFFR_X1 port map( D => n5023, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6851, QN => n_4184);
   clk_r_REG13492_S9 : DFFR_X1 port map( D => n5022, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6850, QN => n_4185);
   clk_r_REG13493_S9 : DFFR_X1 port map( D => n5021, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6849, QN => n_4186);
   clk_r_REG13550_S3 : DFFR_X1 port map( D => n5020, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6848, QN => n_4187);
   clk_r_REG13494_S9 : DFFR_X1 port map( D => n5019, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6847, QN => n_4188);
   clk_r_REG13495_S9 : DFFR_X1 port map( D => n5018, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6846, QN => n_4189);
   clk_r_REG13496_S9 : DFFR_X1 port map( D => n5017, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6845, QN => n_4190);
   clk_r_REG13497_S9 : DFFR_X1 port map( D => n5016, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6844, QN => n_4191);
   clk_r_REG13498_S9 : DFFR_X1 port map( D => n5015, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6843, QN => n_4192);
   clk_r_REG13551_S3 : DFFR_X1 port map( D => n5014, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6842, QN => n_4193);
   clk_r_REG13552_S3 : DFFR_X1 port map( D => n5013, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6841, QN => n_4194);
   clk_r_REG13488_S9 : DFFR_X1 port map( D => n5012, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6840, QN => n_4195);
   clk_r_REG13485_S9 : DFFR_X1 port map( D => n5011, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6839, QN => n_4196);
   clk_r_REG13553_S3 : DFFR_X1 port map( D => n5010, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6838, QN => n_4197);
   clk_r_REG13529_S9 : DFFR_X1 port map( D => n5009, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n6837, QN => n_4198);
   clk_r_REG13419_S3 : DFFR_X1 port map( D => n5006, CK => CLK, RN => RST, Q =>
                           n6836, QN => n_4199);
   clk_r_REG13417_S3 : DFFS_X1 port map( D => n5285, CK => CLK, SN => RST, Q =>
                           n6835, QN => n_4200);
   clk_r_REG13474_S6 : DFFR_X1 port map( D => n7708, CK => CLK, RN => RST, Q =>
                           n_4201, QN => n6834);
   clk_r_REG13421_S2 : DFFR_X1 port map( D => n7706, CK => CLK, RN => RST, Q =>
                           n_4202, QN => n8076);
   clk_r_REG13555_S7 : DFFS_X1 port map( D => n5880, CK => CLK, SN => RST, Q =>
                           n6832, QN => n_4203);
   clk_r_REG13562_S7 : DFFR_X1 port map( D => n7736, CK => CLK, RN => RST, Q =>
                           n7363, QN => n6831);
   clk_r_REG13556_S1 : DFFR_X1 port map( D => n4060, CK => CLK, RN => RST, Q =>
                           n_4204, QN => n7369);
   clk_r_REG11935_S5 : DFFR_X1 port map( D => n7712, CK => CLK, RN => RST, Q =>
                           n_4205, QN => n6829);
   clk_r_REG11937_S6 : DFFS_X1 port map( D => n6829, CK => CLK, SN => RST, Q =>
                           n6828, QN => n_4206);
   clk_r_REG11938_S7 : DFFS_X1 port map( D => n6828, CK => CLK, SN => RST, Q =>
                           n6827, QN => n_4207);
   clk_r_REG13277_S8 : DFFR_X1 port map( D => n7711, CK => CLK, RN => RST, Q =>
                           n_4208, QN => n6826);
   clk_r_REG13279_S9 : DFFS_X1 port map( D => n6826, CK => CLK, SN => RST, Q =>
                           n6825, QN => n_4209);
   clk_r_REG13280_S10 : DFFS_X1 port map( D => n6825, CK => CLK, SN => RST, Q 
                           => n6824, QN => n_4210);
   clk_r_REG10850_S3 : DFFS_X1 port map( D => n4989, CK => CLK, SN => RST, Q =>
                           n6823, QN => n_4211);
   clk_r_REG10312_S3 : DFFS_X1 port map( D => n7702, CK => CLK, SN => RST, Q =>
                           n_4212, QN => n6822);
   clk_r_REG10317_S5 : DFFR_X1 port map( D => n4987, CK => CLK, RN => RST, Q =>
                           n6821, QN => n_4213);
   clk_r_REG11357_S5 : DFFR_X1 port map( D => n4986, CK => CLK, RN => RST, Q =>
                           n6820, QN => n_4214);
   clk_r_REG10958_S12 : DFFR_X1 port map( D => n4985, CK => CLK, RN => RST, Q 
                           => n6819, QN => n_4215);
   clk_r_REG11144_S13 : DFFR_X1 port map( D => n4984, CK => CLK, RN => RST, Q 
                           => n6818, QN => n_4216);
   clk_r_REG11127_S13 : DFFR_X1 port map( D => n4983, CK => CLK, RN => RST, Q 
                           => n6817, QN => n_4217);
   clk_r_REG11120_S6 : DFFR_X1 port map( D => n4982, CK => CLK, RN => RST, Q =>
                           n6816, QN => n_4218);
   clk_r_REG11113_S6 : DFFR_X1 port map( D => n4981, CK => CLK, RN => RST, Q =>
                           n6815, QN => n_4219);
   clk_r_REG11107_S7 : DFFR_X1 port map( D => n4980, CK => CLK, RN => RST, Q =>
                           n6814, QN => n_4220);
   clk_r_REG11100_S6 : DFFR_X1 port map( D => n4979, CK => CLK, RN => RST, Q =>
                           n6813, QN => n_4221);
   clk_r_REG11094_S6 : DFFR_X1 port map( D => n4978, CK => CLK, RN => RST, Q =>
                           n6812, QN => n_4222);
   clk_r_REG11088_S6 : DFFR_X1 port map( D => n4977, CK => CLK, RN => RST, Q =>
                           n6811, QN => n_4223);
   clk_r_REG11082_S6 : DFFR_X1 port map( D => n4976, CK => CLK, RN => RST, Q =>
                           n6810, QN => n_4224);
   clk_r_REG11075_S6 : DFFR_X1 port map( D => n4975, CK => CLK, RN => RST, Q =>
                           n6809, QN => n_4225);
   clk_r_REG13374_S1 : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK => CLK, 
                           RN => RST, Q => n6807, QN => n_4226);
   clk_r_REG11649_S5 : DFFS_X1 port map( D => n4972, CK => CLK, SN => RST, Q =>
                           n6806, QN => n_4227);
   clk_r_REG11352_S5 : DFFS_X1 port map( D => n4971, CK => CLK, SN => RST, Q =>
                           n6805, QN => n_4228);
   clk_r_REG11362_S5 : DFFS_X1 port map( D => n4970, CK => CLK, SN => RST, Q =>
                           n6804, QN => n_4229);
   clk_r_REG10954_S12 : DFFS_X1 port map( D => n4969, CK => CLK, SN => RST, Q 
                           => n6803, QN => n_4230);
   clk_r_REG10964_S12 : DFFS_X1 port map( D => n4968, CK => CLK, SN => RST, Q 
                           => n6802, QN => n_4231);
   clk_r_REG11138_S13 : DFFS_X1 port map( D => n4966, CK => CLK, SN => RST, Q 
                           => n6801, QN => n_4232);
   clk_r_REG10973_S13 : DFFS_X1 port map( D => n4965, CK => CLK, SN => RST, Q 
                           => n6800, QN => n_4233);
   clk_r_REG11009_S16 : DFFS_X1 port map( D => n4964, CK => CLK, SN => RST, Q 
                           => n6799, QN => n_4234);
   clk_r_REG11019_S16 : DFFS_X1 port map( D => n4963, CK => CLK, SN => RST, Q 
                           => n6798, QN => n_4235);
   clk_r_REG11026_S16 : DFFS_X1 port map( D => n4962, CK => CLK, SN => RST, Q 
                           => n6797, QN => n_4236);
   clk_r_REG11037_S16 : DFFS_X1 port map( D => n4961, CK => CLK, SN => RST, Q 
                           => n6796, QN => n_4237);
   clk_r_REG11046_S16 : DFFS_X1 port map( D => n4960, CK => CLK, SN => RST, Q 
                           => n6795, QN => n_4238);
   clk_r_REG11054_S16 : DFFS_X1 port map( D => n4959, CK => CLK, SN => RST, Q 
                           => n6794, QN => n_4239);
   clk_r_REG11061_S16 : DFFS_X1 port map( D => n4958, CK => CLK, SN => RST, Q 
                           => n6793, QN => n_4240);
   clk_r_REG11068_S16 : DFFS_X1 port map( D => n4957, CK => CLK, SN => RST, Q 
                           => n6792, QN => n_4241);
   clk_r_REG11790_S5 : DFFR_X1 port map( D => n4956, CK => CLK, RN => RST, Q =>
                           n6791, QN => n_4242);
   clk_r_REG13372_S1 : DFFS_X1 port map( D => n4954, CK => CLK, SN => RST, Q =>
                           n6790, QN => n_4243);
   clk_r_REG13415_S2 : DFFR_X1 port map( D => n7701, CK => CLK, RN => RST, Q =>
                           n_4244, QN => n6789);
   clk_r_REG13413_S1 : DFFR_X1 port map( D => n302, CK => CLK, RN => RST, Q => 
                           n6788, QN => n_4245);
   clk_r_REG10953_S12 : DFFR_X1 port map( D => n1449, CK => CLK, RN => RST, Q 
                           => IRAM_ADDRESS_8_port, QN => n_4246);
   clk_r_REG10968_S14 : DFFR_X1 port map( D => n1447, CK => CLK, RN => RST, Q 
                           => IRAM_ADDRESS_10_port, QN => n_4247);
   clk_r_REG11131_S5 : DFFR_X1 port map( D => n7715, CK => CLK, RN => RST, Q =>
                           n_4248, QN => n6785);
   clk_r_REG11130_S5 : DFFS_X1 port map( D => n7715, CK => CLK, SN => RST, Q =>
                           n_4249, QN => n6784);
   clk_r_REG11145_S5 : DFFS_X1 port map( D => n7713, CK => CLK, SN => RST, Q =>
                           n_4250, QN => n6783);
   clk_r_REG11141_S14 : DFFR_X1 port map( D => n1445, CK => CLK, RN => RST, Q 
                           => n_4251, QN => n7312);
   clk_r_REG10975_S14 : DFFS_X1 port map( D => n7764, CK => CLK, SN => RST, Q 
                           => n_4252, QN => n6781);
   clk_r_REG11007_S15 : DFFS_X1 port map( D => n7753, CK => CLK, SN => RST, Q 
                           => n_4253, QN => n6780);
   clk_r_REG11017_S15 : DFFS_X1 port map( D => n7754, CK => CLK, SN => RST, Q 
                           => n_4254, QN => n6779);
   clk_r_REG11024_S15 : DFFS_X1 port map( D => n7755, CK => CLK, SN => RST, Q 
                           => n_4255, QN => n6778);
   clk_r_REG11035_S15 : DFFS_X1 port map( D => n7757, CK => CLK, SN => RST, Q 
                           => n_4256, QN => n6777);
   clk_r_REG11044_S15 : DFFS_X1 port map( D => n7758, CK => CLK, SN => RST, Q 
                           => n_4257, QN => n6776);
   clk_r_REG11052_S15 : DFFS_X1 port map( D => n7759, CK => CLK, SN => RST, Q 
                           => n_4258, QN => n6775);
   clk_r_REG11059_S15 : DFFS_X1 port map( D => n7760, CK => CLK, SN => RST, Q 
                           => n_4259, QN => n6774);
   clk_r_REG11066_S15 : DFFS_X1 port map( D => n7761, CK => CLK, SN => RST, Q 
                           => n_4260, QN => n6773);
   clk_r_REG11070_S15 : DFFR_X1 port map( D => n5542, CK => CLK, RN => RST, Q 
                           => n6772, QN => n_4261);
   clk_r_REG11063_S5 : DFFR_X1 port map( D => n7729, CK => CLK, RN => RST, Q =>
                           n_4262, QN => n6771);
   clk_r_REG11062_S5 : DFFS_X1 port map( D => n7729, CK => CLK, SN => RST, Q =>
                           n_4263, QN => n6770);
   clk_r_REG11056_S5 : DFFR_X1 port map( D => n7731, CK => CLK, RN => RST, Q =>
                           n_4264, QN => n6769);
   clk_r_REG11055_S5 : DFFS_X1 port map( D => n7731, CK => CLK, SN => RST, Q =>
                           n_4265, QN => n6768);
   clk_r_REG11048_S5 : DFFR_X1 port map( D => n7727, CK => CLK, RN => RST, Q =>
                           n_4266, QN => n6767);
   clk_r_REG11047_S5 : DFFS_X1 port map( D => n7727, CK => CLK, SN => RST, Q =>
                           n_4267, QN => n6766);
   clk_r_REG11039_S5 : DFFR_X1 port map( D => n7725, CK => CLK, RN => RST, Q =>
                           n_4268, QN => n6765);
   clk_r_REG11038_S5 : DFFS_X1 port map( D => n7725, CK => CLK, SN => RST, Q =>
                           n_4269, QN => n6764);
   clk_r_REG11028_S5 : DFFR_X1 port map( D => n7721, CK => CLK, RN => RST, Q =>
                           n_4270, QN => n6763);
   clk_r_REG11027_S5 : DFFS_X1 port map( D => n7721, CK => CLK, SN => RST, Q =>
                           n_4271, QN => n6762);
   clk_r_REG11021_S6 : DFFR_X1 port map( D => n7719, CK => CLK, RN => RST, Q =>
                           n_4272, QN => n6761);
   clk_r_REG11020_S6 : DFFS_X1 port map( D => n7719, CK => CLK, SN => RST, Q =>
                           n_4273, QN => n6760);
   clk_r_REG11011_S5 : DFFR_X1 port map( D => n7723, CK => CLK, RN => RST, Q =>
                           n_4274, QN => n6759);
   clk_r_REG11010_S5 : DFFS_X1 port map( D => n7723, CK => CLK, SN => RST, Q =>
                           n_4275, QN => n6758);
   clk_r_REG10978_S5 : DFFR_X1 port map( D => n7717, CK => CLK, RN => RST, Q =>
                           n_4276, QN => n6757);
   clk_r_REG10977_S5 : DFFS_X1 port map( D => n7717, CK => CLK, SN => RST, Q =>
                           n_4277, QN => n6756);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => n7695, ADD_WR(3) => n7697, ADD_WR(2) =>
                           n4953, ADD_WR(1) => n7698, ADD_WR(0) => n7696, 
                           ADD_RD1(4) => n5049, ADD_RD1(3) => n5048, ADD_RD1(2)
                           => n5079, ADD_RD1(1) => n5047, ADD_RD1(0) => n5046, 
                           ADD_RD2(4) => curr_instruction_to_cu_i_20_port, 
                           ADD_RD2(3) => curr_instruction_to_cu_i_19_port, 
                           ADD_RD2(2) => n7756, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n43, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n44, OUT1(31) => n1673, 
                           OUT1(30) => n1671, OUT1(29) => n1669, OUT1(28) => 
                           n1667, OUT1(27) => n1665, OUT1(26) => n1663, 
                           OUT1(25) => n1661, OUT1(24) => n1659, OUT1(23) => 
                           n1657, OUT1(22) => n1655, OUT1(21) => n1653, 
                           OUT1(20) => n1651, OUT1(19) => n1649, OUT1(18) => 
                           n1647, OUT1(17) => n1645, OUT1(16) => n1643, 
                           OUT1(15) => n1641, OUT1(14) => n1639, OUT1(13) => 
                           n1637, OUT1(12) => n1635, OUT1(11) => n1633, 
                           OUT1(10) => n1631, OUT1(9) => n1629, OUT1(8) => 
                           n1627, OUT1(7) => n1625, OUT1(6) => n1623, OUT1(5) 
                           => n1621, OUT1(4) => n1619, OUT1(3) => n1617, 
                           OUT1(2) => n1615, OUT1(1) => n1614, OUT1(0) => n1613
                           , OUT2(31) => n5229, OUT2(30) => n5226, OUT2(29) => 
                           n5223, OUT2(28) => n5220, OUT2(27) => n5217, 
                           OUT2(26) => n5214, OUT2(25) => n5211, OUT2(24) => 
                           n5208, OUT2(23) => n5205, OUT2(22) => n5202, 
                           OUT2(21) => n5199, OUT2(20) => n5196, OUT2(19) => 
                           n5193, OUT2(18) => n5190, OUT2(17) => n5187, 
                           OUT2(16) => n5184, OUT2(15) => n5181, OUT2(14) => 
                           n5178, OUT2(13) => n5175, OUT2(12) => n5172, 
                           OUT2(11) => n5169, OUT2(10) => n5166, OUT2(9) => 
                           n5163, OUT2(8) => n5160, OUT2(7) => n5157, OUT2(6) 
                           => n5154, OUT2(5) => n5151, OUT2(4) => n5148, 
                           OUT2(3) => n5145, OUT2(2) => n5142, OUT2(1) => n5139
                           , OUT2(0) => n5136, RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_4278, mul_exeception => 
                           n_4279, FUNC(0) => n7700, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_4280, 
                           OUTALU(31) => datapath_i_alu_output_val_i_31_port, 
                           OUTALU(30) => datapath_i_alu_output_val_i_30_port, 
                           OUTALU(29) => datapath_i_alu_output_val_i_29_port, 
                           OUTALU(28) => datapath_i_alu_output_val_i_28_port, 
                           OUTALU(27) => datapath_i_alu_output_val_i_27_port, 
                           OUTALU(26) => datapath_i_alu_output_val_i_26_port, 
                           OUTALU(25) => datapath_i_alu_output_val_i_25_port, 
                           OUTALU(24) => datapath_i_alu_output_val_i_24_port, 
                           OUTALU(23) => datapath_i_alu_output_val_i_23_port, 
                           OUTALU(22) => datapath_i_alu_output_val_i_22_port, 
                           OUTALU(21) => datapath_i_alu_output_val_i_21_port, 
                           OUTALU(20) => datapath_i_alu_output_val_i_20_port, 
                           OUTALU(19) => datapath_i_alu_output_val_i_19_port, 
                           OUTALU(18) => datapath_i_alu_output_val_i_18_port, 
                           OUTALU(17) => datapath_i_alu_output_val_i_17_port, 
                           OUTALU(16) => datapath_i_alu_output_val_i_16_port, 
                           OUTALU(15) => datapath_i_alu_output_val_i_15_port, 
                           OUTALU(14) => datapath_i_alu_output_val_i_14_port, 
                           OUTALU(13) => datapath_i_alu_output_val_i_13_port, 
                           OUTALU(12) => datapath_i_alu_output_val_i_12_port, 
                           OUTALU(11) => datapath_i_alu_output_val_i_11_port, 
                           OUTALU(10) => datapath_i_alu_output_val_i_10_port, 
                           OUTALU(9) => datapath_i_alu_output_val_i_9_port, 
                           OUTALU(8) => datapath_i_alu_output_val_i_8_port, 
                           OUTALU(7) => datapath_i_alu_output_val_i_7_port, 
                           OUTALU(6) => datapath_i_alu_output_val_i_6_port, 
                           OUTALU(5) => datapath_i_alu_output_val_i_5_port, 
                           OUTALU(4) => datapath_i_alu_output_val_i_4_port, 
                           OUTALU(3) => datapath_i_alu_output_val_i_3_port, 
                           OUTALU(2) => datapath_i_alu_output_val_i_2_port, 
                           OUTALU(1) => datapath_i_alu_output_val_i_1_port, 
                           OUTALU(0) => datapath_i_alu_output_val_i_0_port, 
                           rst_BAR => RST);
   U3044 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_31_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(31), ZN => n7525
                           );
   U3046 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_30_port, A2 => 
                           n7557, B1 => n8084, B2 => DRAM_DATA(30), ZN => n7526
                           );
   U3048 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_29_port, A2 => 
                           n8083, B1 => n8084, B2 => DRAM_DATA(29), ZN => n7527
                           );
   U3050 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_28_port, A2 => 
                           n8083, B1 => n8084, B2 => DRAM_DATA(28), ZN => n7528
                           );
   U3052 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_27_port, A2 => 
                           n8083, B1 => n8084, B2 => DRAM_DATA(27), ZN => n7529
                           );
   U3054 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_26_port, A2 => 
                           n8083, B1 => n8084, B2 => DRAM_DATA(26), ZN => n7530
                           );
   U3056 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_25_port, A2 => 
                           n7557, B1 => n8084, B2 => DRAM_DATA(25), ZN => n7531
                           );
   U3058 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_24_port, A2 => 
                           n8083, B1 => n8084, B2 => DRAM_DATA(24), ZN => n7532
                           );
   U3060 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_23_port, A2 => 
                           n8083, B1 => n8084, B2 => DRAM_DATA(23), ZN => n7533
                           );
   U3062 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_22_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(22), ZN => n7534
                           );
   U3064 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_21_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(21), ZN => n7535
                           );
   U3066 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(20), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_20_port, ZN => n7536)
                           ;
   U3068 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(19), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_19_port, ZN => n7537)
                           ;
   U3070 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(18), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_18_port, ZN => n7538)
                           ;
   U3072 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(17), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_17_port, ZN => n7539)
                           ;
   U3074 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(16), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_16_port, ZN => n7540)
                           ;
   U3076 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(15), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_15_port, ZN => n7541)
                           ;
   U3078 : AOI22_X1 port map( A1 => n7556, A2 => DRAM_DATA(14), B1 => n8083, B2
                           => datapath_i_alu_output_val_i_14_port, ZN => n7542)
                           ;
   U3080 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_13_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(13), ZN => n7543
                           );
   U3082 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_12_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(12), ZN => n7544
                           );
   U3084 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_11_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(11), ZN => n7545
                           );
   U3086 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_10_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(10), ZN => n7546
                           );
   U3088 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_9_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(9), ZN => n7547)
                           ;
   U3090 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_8_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(8), ZN => n7548)
                           ;
   U3092 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_7_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(7), ZN => n7549)
                           ;
   U3094 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_6_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(6), ZN => n7550)
                           ;
   U3096 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_5_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(5), ZN => n7551)
                           ;
   U3098 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_4_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(4), ZN => n7552)
                           ;
   U3100 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_3_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(3), ZN => n7553)
                           ;
   U3102 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_2_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(2), ZN => n7554)
                           ;
   U3104 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_1_port, A2 => 
                           n7557, B1 => n7556, B2 => DRAM_DATA(1), ZN => n7555)
                           ;
   U3106 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_0_port, A2 => 
                           n8083, B1 => n7556, B2 => DRAM_DATA(0), ZN => n7558)
                           ;
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => n3284);
   clk_r_REG13299_S4 : DFFS_X1 port map( D => n4337, CK => CLK, SN => RST, Q =>
                           n_4281, QN => n7277);
   clk_r_REG10373_S2 : DFF_X1 port map( D => n1673, CK => CLK, Q => n7094, QN 
                           => n_4282);
   clk_r_REG13535_S2 : DFFS_X1 port map( D => n6178, CK => CLK, SN => RST, Q =>
                           n8072, QN => n7250);
   clk_r_REG13478_S6 : DFFS_X1 port map( D => n4974, CK => CLK, SN => RST, Q =>
                           n6808, QN => n_4283);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => n6894, Q => 
                           n5388);
   clk_r_REG13625_S7 : DFFR_X1 port map( D => n5069, CK => CLK, RN => RST, Q =>
                           n6887, QN => n_4284);
   clk_r_REG13302_S4 : DFFR_X1 port map( D => n7704, CK => CLK, RN => RST, Q =>
                           n7202, QN => n_4285);
   clk_r_REG13300_S4 : DFFR_X1 port map( D => n7704, CK => CLK, RN => RST, Q =>
                           n_4286, QN => n7275);
   clk_r_REG13424_S2 : DFFS_X1 port map( D => n5405, CK => CLK, SN => RST, Q =>
                           n7215, QN => n_4287);
   clk_r_REG10315_S4 : DFFR_X1 port map( D => n7348, CK => CLK, RN => RST, Q =>
                           n_4288, QN => n7107);
   clk_r_REG13481_S6 : DFFR_X1 port map( D => n5388, CK => CLK, RN => RST, Q =>
                           n7200, QN => n_4289);
   clk_r_REG13473_S6 : DFFS_X1 port map( D => n7709, CK => CLK, SN => RST, Q =>
                           n_4290, QN => n6937);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X2 port map( A => 
                           n6990, EN => n7215, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X2 port map( A => 
                           n6987, EN => n6935, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X2 port map( A => 
                           n6999, EN => n7198, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X2 port map( A => 
                           n7005, EN => n7215, Z => DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X2 port map( A => 
                           n7002, EN => n7215, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X2 port map( A => 
                           n6993, EN => n7215, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X2 port map( A => 
                           n6996, EN => n6935, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X2 port map( A => 
                           n7035, EN => n7215, Z => DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X2 port map( A => 
                           n7032, EN => n7215, Z => DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X2 port map( A => 
                           n7029, EN => n7215, Z => DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X2 port map( A => 
                           n7026, EN => n7215, Z => DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X2 port map( A => 
                           n7011, EN => n7215, Z => DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X2 port map( A => 
                           n6984, EN => n7215, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X2 port map( A => 
                           n6969, EN => n7215, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X2 port map( A => 
                           n6960, EN => n7215, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X2 port map( A => 
                           n6957, EN => n7215, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X2 port map( A => 
                           n7020, EN => n6935, Z => DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X2 port map( A => 
                           n6981, EN => n6935, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X2 port map( A => 
                           n6975, EN => n6935, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X2 port map( A => 
                           n6963, EN => n6935, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X2 port map( A => 
                           n6954, EN => n6935, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X2 port map( A => 
                           n6951, EN => n6935, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X2 port map( A => 
                           n6948, EN => n6935, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X2 port map( A => 
                           n7038, EN => n7198, Z => DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X2 port map( A => 
                           n7023, EN => n7198, Z => DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X2 port map( A => 
                           n7017, EN => n7198, Z => DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X2 port map( A => 
                           n7014, EN => n7198, Z => DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X2 port map( A => 
                           n7008, EN => n7198, Z => DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X2 port map( A => 
                           n6978, EN => n7198, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X2 port map( A => 
                           n6972, EN => n7198, Z => DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X2 port map( A => 
                           n6966, EN => n7198, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X2 port map( A => 
                           n6945, EN => n7198, Z => DRAM_DATA(0));
   U3314 : AOI221_X2 port map( B1 => n6880, B2 => n7709, C1 => cu_i_n135, C2 =>
                           n5388, A => n6822, ZN => n4337);
   U3315 : OAI21_X2 port map( B1 => n6920, B2 => n7259, A => n7938, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U3316 : OAI21_X2 port map( B1 => n6920, B2 => n7115, A => n6823, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U3317 : INV_X2 port map( A => n7312, ZN => IRAM_ADDRESS_12_port);
   U3318 : AOI22_X1 port map( A1 => n6937, A2 => cu_i_cmd_alu_op_type_3_port, 
                           B1 => n7095, B2 => n6938, ZN => n7886);
   U3319 : AOI22_X1 port map( A1 => n6937, A2 => cu_i_cmd_alu_op_type_2_port, 
                           B1 => n7095, B2 => n6939, ZN => n7887);
   U3320 : NOR2_X1 port map( A1 => n7887, A2 => n7888, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U3321 : NOR2_X1 port map( A1 => n7890, A2 => n7884, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U3322 : CLKBUF_X1 port map( A => n6808, Z => n8031);
   U3323 : MUX2_X1 port map( A => n6839, B => n6958, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U3324 : MUX2_X1 port map( A => IRAM_DATA(23), B => n6881, S => n6937, Z => 
                           n5079);
   U3325 : INV_X1 port map( A => n5388, ZN => n7709);
   U3326 : NOR2_X1 port map( A1 => n5388, A2 => n6926, ZN => n7858);
   U3327 : AOI21_X1 port map( B1 => n5388, B2 => n7096, A => n7858, ZN => n7789
                           );
   U3328 : INV_X1 port map( A => n7789, ZN => n7703);
   U3329 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(29), B1 => n7200, B2
                           => n7266, ZN => n8020);
   U3330 : INV_X1 port map( A => n8020, ZN => n7746);
   U3331 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(30), B1 => n7200, B2
                           => n7267, ZN => n7796);
   U3332 : INV_X1 port map( A => n7796, ZN => n7747);
   U3333 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(31), B1 => n7200, B2
                           => n7258, ZN => n7800);
   U3334 : NAND3_X1 port map( A1 => n7746, A2 => n7747, A3 => n7800, ZN => 
                           n7799);
   U3335 : INV_X1 port map( A => n7799, ZN => n7745);
   U3336 : CLKBUF_X1 port map( A => n7250, Z => n8080);
   U3337 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(28), B1 => n8070, B2
                           => n8066, ZN => n7750);
   U3338 : NAND3_X1 port map( A1 => n7800, A2 => n7796, A3 => n7746, ZN => 
                           n7985);
   U3339 : OR2_X1 port map( A1 => n7985, A2 => n7750, ZN => n2299);
   U3340 : NAND2_X1 port map( A1 => n6781, A2 => n6916, ZN => n7861);
   U3341 : NOR2_X1 port map( A1 => n6757, A2 => n7861, ZN => n7860);
   U3342 : NAND2_X1 port map( A1 => n7860, A2 => n6780, ZN => n7870);
   U3343 : OAI211_X1 port map( C1 => n7860, C2 => n6780, A => n7201, B => n7870
                           , ZN => n7790);
   U3344 : NAND2_X1 port map( A1 => n6799, A2 => n7790, ZN => n7944);
   U3345 : INV_X1 port map( A => n7944, ZN => n7785);
   U3346 : INV_X1 port map( A => datapath_i_alu_output_val_i_16_port, ZN => 
                           n7791);
   U3347 : OAI222_X1 port map( A1 => n7791, A2 => n7148, B1 => n7107, B2 => 
                           n7261, C1 => n7785, C2 => n7166, ZN => n5342);
   U3348 : INV_X1 port map( A => n5342, ZN => n7753);
   U3349 : NOR2_X1 port map( A1 => n6759, A2 => n7870, ZN => n7869);
   U3350 : NAND2_X1 port map( A1 => n7869, A2 => n6779, ZN => n7873);
   U3351 : OAI211_X1 port map( C1 => n7869, C2 => n6779, A => n7201, B => n7873
                           , ZN => n7792);
   U3352 : NAND2_X1 port map( A1 => n6798, A2 => n7792, ZN => n7937);
   U3353 : INV_X1 port map( A => n7937, ZN => n7784);
   U3354 : INV_X1 port map( A => datapath_i_alu_output_val_i_18_port, ZN => 
                           n7793);
   U3355 : OAI222_X1 port map( A1 => n7793, A2 => n7148, B1 => n7107, B2 => 
                           n7259, C1 => n7784, C2 => n7166, ZN => n5343);
   U3356 : INV_X1 port map( A => n5343, ZN => n7754);
   U3357 : INV_X1 port map( A => n7800, ZN => n7744);
   U3358 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(26), B1 => n8069, B2
                           => n8066, ZN => n7751);
   U3359 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(27), B1 => n7200, B2
                           => n7264, ZN => n7812);
   U3360 : INV_X1 port map( A => n7750, ZN => n8054);
   U3361 : NOR2_X1 port map( A1 => n7812, A2 => n8054, ZN => n7987);
   U3362 : INV_X1 port map( A => n7751, ZN => n7986);
   U3363 : AND4_X1 port map( A1 => n7796, A2 => n7987, A3 => n7744, A4 => n7986
                           , ZN => n7816);
   U3364 : NAND2_X1 port map( A1 => n6903, A2 => n7816, ZN => n8019);
   U3365 : NOR2_X1 port map( A1 => n7746, A2 => n8019, ZN => 
                           cu_i_cmd_word_3_port);
   U3366 : OAI22_X1 port map( A1 => n7709, A2 => cu_i_cmd_word_3_port, B1 => 
                           n6879, B2 => n5388, ZN => n7809);
   U3367 : INV_X1 port map( A => n7809, ZN => n7707);
   U3368 : OAI211_X1 port map( C1 => n6781, C2 => n6916, A => n7201, B => n7861
                           , ZN => n7794);
   U3369 : NAND2_X1 port map( A1 => n6800, A2 => n7794, ZN => n7917);
   U3370 : INV_X1 port map( A => n7917, ZN => n7777);
   U3371 : INV_X1 port map( A => datapath_i_alu_output_val_i_14_port, ZN => 
                           n7795);
   U3372 : OAI222_X1 port map( A1 => n7795, A2 => n7148, B1 => n7107, B2 => 
                           n7218, C1 => n7777, C2 => n7166, ZN => n1443);
   U3373 : INV_X1 port map( A => n1443, ZN => n7764);
   U3374 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(0), B1 => n7200, B2 
                           => n7106, ZN => n7804);
   U3375 : INV_X1 port map( A => n7804, ZN => n7736);
   U3376 : NAND3_X1 port map( A1 => n8020, A2 => n7800, A3 => n7796, ZN => 
                           n7797);
   U3377 : NOR2_X1 port map( A1 => n7797, A2 => n8067, ZN => n7813);
   U3378 : NAND2_X1 port map( A1 => n7813, A2 => n7987, ZN => n6178);
   U3379 : NAND2_X1 port map( A1 => n7812, A2 => n7751, ZN => n7739);
   U3380 : NOR3_X1 port map( A1 => n7797, A2 => n7739, A3 => n8054, ZN => n5880
                           );
   U3381 : INV_X1 port map( A => n5880, ZN => n7900);
   U3382 : NOR2_X1 port map( A1 => n7900, A2 => n8067, ZN => n7738);
   U3383 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(1), B1 => n8073, B2 
                           => n8066, ZN => n7748);
   U3384 : MUX2_X1 port map( A => IRAM_DATA(4), B => n6900, S => n7200, Z => 
                           n5076);
   U3385 : MUX2_X1 port map( A => IRAM_DATA(3), B => n6898, S => n7200, Z => 
                           n5077);
   U3386 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(2), B1 => n8074, B2 
                           => n8066, ZN => n7749);
   U3387 : AOI22_X1 port map( A1 => n7269, A2 => IRAM_DATA(5), B1 => n7200, B2 
                           => n7257, ZN => n7798);
   U3388 : INV_X1 port map( A => n7798, ZN => n7735);
   U3389 : INV_X1 port map( A => n7812, ZN => n7741);
   U3390 : AOI211_X1 port map( C1 => n7750, C2 => n7751, A => n7741, B => n7799
                           , ZN => n4060);
   U3391 : NAND2_X1 port map( A1 => n7800, A2 => n7747, ZN => n7801);
   U3392 : NOR4_X1 port map( A1 => n7750, A2 => n7986, A3 => n7746, A4 => n7801
                           , ZN => n5075);
   U3393 : INV_X1 port map( A => n7738, ZN => n7989);
   U3394 : INV_X1 port map( A => n7749, ZN => n7802);
   U3395 : NAND4_X1 port map( A1 => n5076, A2 => n5077, A3 => n7802, A4 => 
                           n7735, ZN => n7803);
   U3396 : NOR3_X1 port map( A1 => n7804, A2 => n7748, A3 => n7803, ZN => n7848
                           );
   U3397 : NAND2_X1 port map( A1 => n7812, A2 => n8054, ZN => n7805);
   U3398 : AOI21_X1 port map( B1 => n7986, B2 => n7805, A => n7985, ZN => n7806
                           );
   U3399 : NOR3_X1 port map( A1 => n4060, A2 => n5075, A3 => n7806, ZN => n7896
                           );
   U3400 : OAI222_X1 port map( A1 => n6178, A2 => n7751, B1 => n7989, B2 => 
                           n7848, C1 => n7164, C2 => n7896, ZN => n302);
   U3401 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n302, ZN => n5122
                           );
   U3402 : NOR2_X1 port map( A1 => n6761, A2 => n7873, ZN => n7872);
   U3403 : NAND2_X1 port map( A1 => n7872, A2 => n6778, ZN => n7882);
   U3404 : OAI211_X1 port map( C1 => n7872, C2 => n6778, A => n7201, B => n7882
                           , ZN => n7807);
   U3405 : NAND2_X1 port map( A1 => n6797, A2 => n7807, ZN => n7951);
   U3406 : INV_X1 port map( A => n7951, ZN => n7783);
   U3407 : INV_X1 port map( A => datapath_i_alu_output_val_i_20_port, ZN => 
                           n7808);
   U3408 : OAI222_X1 port map( A1 => n7808, A2 => n7148, B1 => n7107, B2 => 
                           n7255, C1 => n7783, C2 => n7166, ZN => n5344);
   U3409 : INV_X1 port map( A => n5344, ZN => n7755);
   U3410 : INV_X1 port map( A => n8019, ZN => n7740);
   U3411 : OAI22_X1 port map( A1 => n7709, A2 => n7740, B1 => n6878, B2 => 
                           n5388, ZN => n5358);
   U3412 : INV_X1 port map( A => n5358, ZN => n7706);
   U3413 : NAND2_X1 port map( A1 => n7706, A2 => n7809, ZN => n5405);
   U3414 : INV_X1 port map( A => n5405, ZN => n7705);
   U3415 : MUX2_X1 port map( A => IRAM_DATA(11), B => n6889, S => n7200, Z => 
                           n5071);
   U3416 : MUX2_X1 port map( A => IRAM_DATA(12), B => n6892, S => n6937, Z => 
                           n5065);
   U3417 : AOI22_X1 port map( A1 => n6937, A2 => n7268, B1 => n7095, B2 => 
                           IRAM_DATA(13), ZN => n7823);
   U3418 : INV_X1 port map( A => n7823, ZN => n7752);
   U3419 : MUX2_X1 port map( A => IRAM_DATA(14), B => n6890, S => n6937, Z => 
                           n5067);
   U3420 : AOI22_X1 port map( A1 => n6937, A2 => n7254, B1 => n7095, B2 => 
                           IRAM_DATA(18), ZN => n7824);
   U3421 : INV_X1 port map( A => n7824, ZN => n7756);
   U3422 : MUX2_X1 port map( A => IRAM_DATA(19), B => n6891, S => n6937, Z => 
                           curr_instruction_to_cu_i_19_port);
   U3423 : NOR2_X1 port map( A1 => n6763, A2 => n7882, ZN => n7881);
   U3424 : NAND2_X1 port map( A1 => n7881, A2 => n6777, ZN => n7879);
   U3425 : OAI211_X1 port map( C1 => n7881, C2 => n6777, A => n7201, B => n7879
                           , ZN => n7810);
   U3426 : NAND2_X1 port map( A1 => n6796, A2 => n7810, ZN => n8036);
   U3427 : INV_X1 port map( A => n8036, ZN => n7782);
   U3428 : INV_X1 port map( A => datapath_i_alu_output_val_i_22_port, ZN => 
                           n7811);
   U3429 : OAI222_X1 port map( A1 => n7811, A2 => n7148, B1 => n7107, B2 => 
                           n7252, C1 => n7782, C2 => n7166, ZN => n5345);
   U3430 : INV_X1 port map( A => n5345, ZN => n7757);
   U3431 : NAND2_X1 port map( A1 => n7812, A2 => n7986, ZN => n474);
   U3432 : NAND2_X1 port map( A1 => n7813, A2 => n8054, ZN => n7847);
   U3433 : NOR2_X1 port map( A1 => n7847, A2 => n474, ZN => n8055);
   U3434 : INV_X1 port map( A => n8055, ZN => n7743);
   U3435 : NOR3_X1 port map( A1 => n7750, A2 => n7739, A3 => n7744, ZN => n7815
                           );
   U3436 : INV_X1 port map( A => n7896, ZN => n7814);
   U3437 : NOR3_X1 port map( A1 => n7816, A2 => n7815, A3 => n7814, ZN => n7901
                           );
   U3438 : OAI211_X1 port map( C1 => n7901, C2 => n8067, A => n7743, B => n6178
                           , ZN => n7737);
   U3439 : CLKBUF_X1 port map( A => n7737, Z => n8082);
   U3440 : NOR2_X1 port map( A1 => n6765, A2 => n7879, ZN => n7878);
   U3441 : NAND2_X1 port map( A1 => n7878, A2 => n6776, ZN => n7876);
   U3442 : OAI211_X1 port map( C1 => n7878, C2 => n6776, A => n7201, B => n7876
                           , ZN => n7817);
   U3443 : NAND2_X1 port map( A1 => n6795, A2 => n7817, ZN => n7935);
   U3444 : INV_X1 port map( A => n7935, ZN => n7781);
   U3445 : INV_X1 port map( A => datapath_i_alu_output_val_i_24_port, ZN => 
                           n7818);
   U3446 : OAI222_X1 port map( A1 => n7818, A2 => n7148, B1 => n7107, B2 => 
                           n7246, C1 => n7781, C2 => n7166, ZN => n5346);
   U3447 : INV_X1 port map( A => n5346, ZN => n7758);
   U3448 : NOR2_X1 port map( A1 => n4417, A2 => n3284, ZN => n7819);
   U3449 : NAND3_X1 port map( A1 => n5131, A2 => n7819, A3 => cu_i_n151, ZN => 
                           n5073);
   U3450 : INV_X1 port map( A => cu_i_n151, ZN => n7699);
   U3451 : OR2_X1 port map( A1 => n7819, A2 => n7699, ZN => n7362);
   U3452 : MUX2_X1 port map( A => IRAM_DATA(20), B => n6888, S => n6937, Z => 
                           curr_instruction_to_cu_i_20_port);
   U3453 : MUX2_X1 port map( A => IRAM_DATA(15), B => n6887, S => n6937, Z => 
                           n5069);
   U3454 : INV_X1 port map( A => n6178, ZN => n7742);
   U3455 : CLKBUF_X1 port map( A => n7742, Z => n8081);
   U3456 : NAND2_X1 port map( A1 => n5073, A2 => n7362, ZN => n7849);
   U3457 : AOI21_X1 port map( B1 => n7848, B2 => n7849, A => n7989, ZN => n7825
                           );
   U3458 : INV_X1 port map( A => n7825, ZN => n8018);
   U3459 : AOI221_X1 port map( B1 => n8018, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n7825, C2 =>
                           n5069, A => n8081, ZN => n7820);
   U3460 : INV_X1 port map( A => n7820, ZN => n7695);
   U3461 : MUX2_X1 port map( A => IRAM_DATA(16), B => n6895, S => n6937, Z => 
                           curr_instruction_to_cu_i_16_port);
   U3462 : AOI221_X1 port map( B1 => n8018, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n7825, C2 =>
                           n5071, A => n8081, ZN => n7821);
   U3463 : INV_X1 port map( A => n7821, ZN => n7696);
   U3464 : MUX2_X1 port map( A => IRAM_DATA(17), B => n6893, S => n6937, Z => 
                           curr_instruction_to_cu_i_17_port);
   U3465 : AOI221_X1 port map( B1 => n8018, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n7825, C2 =>
                           n5065, A => n8081, ZN => n7822);
   U3466 : INV_X1 port map( A => n7822, ZN => n7698);
   U3467 : OAI221_X1 port map( B1 => n7825, B2 => n7824, C1 => n8018, C2 => 
                           n7823, A => n6178, ZN => n4953);
   U3468 : AOI221_X1 port map( B1 => n8018, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n7825, C2 =>
                           n5067, A => n8081, ZN => n7826);
   U3469 : INV_X1 port map( A => n7826, ZN => n7697);
   U3470 : NAND2_X1 port map( A1 => n7738, A2 => n7848, ZN => n5117);
   U3471 : NOR2_X1 port map( A1 => n7362, A2 => n5117, ZN => n7827);
   U3472 : NOR2_X1 port map( A1 => n7827, A2 => n6836, ZN => n7830);
   U3473 : AND3_X1 port map( A1 => n7830, A2 => n7270, A3 => DRAM_READY, ZN => 
                           n7556);
   U3474 : CLKBUF_X1 port map( A => n7556, Z => n8084);
   U3475 : AOI222_X1 port map( A1 => n7204, A2 => n6921, B1 => n7109, B2 => 
                           n7117, C1 => n7205, C2 => 
                           datapath_i_alu_output_val_i_9_port, ZN => n7959);
   U3476 : INV_X1 port map( A => n7959, ZN => n7774);
   U3477 : NOR2_X1 port map( A1 => n6767, A2 => n7876, ZN => n7875);
   U3478 : NAND2_X1 port map( A1 => n7875, A2 => n6775, ZN => n7867);
   U3479 : OAI211_X1 port map( C1 => n7875, C2 => n6775, A => n7201, B => n7867
                           , ZN => n7828);
   U3480 : NAND2_X1 port map( A1 => n6794, A2 => n7828, ZN => n7931);
   U3481 : INV_X1 port map( A => n7931, ZN => n7780);
   U3482 : INV_X1 port map( A => datapath_i_alu_output_val_i_26_port, ZN => 
                           n7829);
   U3483 : OAI222_X1 port map( A1 => n7829, A2 => n7148, B1 => n7107, B2 => 
                           n7244, C1 => n7780, C2 => n7166, ZN => n5347);
   U3484 : INV_X1 port map( A => n5347, ZN => n7759);
   U3485 : AOI222_X1 port map( A1 => n7204, A2 => n6922, B1 => n7109, B2 => 
                           n7114, C1 => n7205, C2 => 
                           datapath_i_alu_output_val_i_7_port, ZN => n7957);
   U3486 : INV_X1 port map( A => n7957, ZN => n7775);
   U3487 : OAI211_X1 port map( C1 => n7901, C2 => n7164, A => n7743, B => n8018
                           , ZN => enable_rf_i);
   U3488 : OAI21_X1 port map( B1 => n7362, B2 => n5117, A => n6835, ZN => 
                           write_rf_i);
   U3489 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U3490 : AOI21_X1 port map( B1 => datapath_i_alu_output_val_i_5_port, B2 => 
                           n7103, A => n7194, ZN => n7958);
   U3491 : INV_X1 port map( A => n7958, ZN => n7786);
   U3492 : NOR2_X1 port map( A1 => n7830, A2 => n7172, ZN => n7557);
   U3493 : CLKBUF_X1 port map( A => n7557, Z => n8083);
   U3494 : NOR2_X1 port map( A1 => n6769, A2 => n7867, ZN => n7866);
   U3495 : NAND2_X1 port map( A1 => n7866, A2 => n6774, ZN => n7864);
   U3496 : OAI211_X1 port map( C1 => n7866, C2 => n6774, A => n7201, B => n7864
                           , ZN => n7831);
   U3497 : NAND2_X1 port map( A1 => n6793, A2 => n7831, ZN => n7929);
   U3498 : INV_X1 port map( A => n7929, ZN => n7779);
   U3499 : INV_X1 port map( A => datapath_i_alu_output_val_i_28_port, ZN => 
                           n7832);
   U3500 : OAI222_X1 port map( A1 => n7832, A2 => n7148, B1 => n7107, B2 => 
                           n7242, C1 => n7779, C2 => n7166, ZN => n5348);
   U3501 : INV_X1 port map( A => n5348, ZN => n7760);
   U3502 : NOR2_X1 port map( A1 => n6771, A2 => n7864, ZN => n7863);
   U3503 : NAND2_X1 port map( A1 => n7863, A2 => n6773, ZN => n7835);
   U3504 : OAI211_X1 port map( C1 => n7863, C2 => n6773, A => n7201, B => n7835
                           , ZN => n7833);
   U3505 : NAND2_X1 port map( A1 => n6792, A2 => n7833, ZN => n7927);
   U3506 : INV_X1 port map( A => n7927, ZN => n7778);
   U3507 : INV_X1 port map( A => datapath_i_alu_output_val_i_30_port, ZN => 
                           n7834);
   U3508 : OAI222_X1 port map( A1 => n7834, A2 => n7148, B1 => n7107, B2 => 
                           n7238, C1 => n7778, C2 => n7166, ZN => n5349);
   U3509 : INV_X1 port map( A => n5349, ZN => n7761);
   U3510 : XOR2_X1 port map( A => n6772, B => n7835, Z => n7836);
   U3511 : AOI22_X1 port map( A1 => n7201, A2 => n7836, B1 => n7274, B2 => 
                           n6908, ZN => n8043);
   U3512 : INV_X1 port map( A => n8043, ZN => n7732);
   U3513 : AOI22_X1 port map( A1 => n7195, A2 => n7168, B1 => 
                           datapath_i_alu_output_val_i_2_port, B2 => n8068, ZN 
                           => n7837);
   U3514 : OAI21_X1 port map( B1 => n7107, B2 => n7235, A => n7837, ZN => n7763
                           );
   U3515 : INV_X1 port map( A => n7311, ZN => IRAM_ADDRESS_1_port);
   U3516 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_1_port, B1 => n7168, B2 
                           => n7179, ZN => n7838);
   U3517 : OAI21_X1 port map( B1 => n7107, B2 => n6827, A => n7838, ZN => n5478
                           );
   U3518 : AOI22_X1 port map( A1 => n7275, A2 => IRAM_ADDRESS_1_port, B1 => 
                           n7197, B2 => n5478, ZN => n7839);
   U3519 : INV_X1 port map( A => n7839, ZN => n7712);
   U3520 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n7168, B2 
                           => n7171, ZN => n7840);
   U3521 : OAI21_X1 port map( B1 => n7107, B2 => n7232, A => n7840, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U3522 : AOI22_X1 port map( A1 => n7205, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n7168, B2 
                           => n7180, ZN => n7841);
   U3523 : OAI21_X1 port map( B1 => n7107, B2 => n7229, A => n7841, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U3524 : NAND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_3_port,
                           A2 => n7763, ZN => n8048);
   U3525 : INV_X1 port map( A => n8048, ZN => n7954);
   U3526 : NAND2_X1 port map( A1 => n7954, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n7953);
   U3527 : NOR2_X1 port map( A1 => n7958, A2 => n7953, ZN => n7940);
   U3528 : AOI211_X1 port map( C1 => n7958, C2 => n7953, A => n7275, B => n7940
                           , ZN => n7842);
   U3529 : OR2_X1 port map( A1 => n6820, A2 => n7842, ZN => n7334);
   U3530 : AOI22_X1 port map( A1 => n7110, A2 => n6904, B1 => n6915, B2 => 
                           n7334, ZN => n7843);
   U3531 : INV_X1 port map( A => n7843, ZN => n7710);
   U3532 : AOI22_X1 port map( A1 => n7205, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n7168, B2 
                           => n7165, ZN => n7844);
   U3533 : OAI21_X1 port map( B1 => n7107, B2 => n7226, A => n7844, ZN => n1453
                           );
   U3534 : INV_X1 port map( A => datapath_i_alu_output_val_i_8_port, ZN => 
                           n7845);
   U3535 : OAI222_X1 port map( A1 => n7845, A2 => n7104, B1 => n7107, B2 => 
                           n7223, C1 => n7225, C2 => n7166, ZN => n1449);
   U3536 : NAND2_X1 port map( A1 => n7940, A2 => n1453, ZN => n7939);
   U3537 : NOR2_X1 port map( A1 => n7957, A2 => n7939, ZN => n7894);
   U3538 : NAND2_X1 port map( A1 => n7894, A2 => n1449, ZN => n7908);
   U3539 : OAI211_X1 port map( C1 => n7894, C2 => n1449, A => n7202, B => n7908
                           , ZN => n7846);
   U3540 : NAND2_X1 port map( A1 => n6803, A2 => n7846, ZN => n7947);
   U3541 : INV_X1 port map( A => n7947, ZN => n7762);
   U3542 : OAI21_X1 port map( B1 => n7739, B2 => n7847, A => n6178, ZN => 
                           cu_i_cmd_word_6_port);
   U3543 : NOR2_X1 port map( A1 => cu_i_cmd_word_6_port, A2 => n8055, ZN => 
                           n7904);
   U3544 : INV_X1 port map( A => n7904, ZN => cu_i_n135);
   U3545 : INV_X1 port map( A => n4337, ZN => n7704);
   U3546 : NAND2_X1 port map( A1 => n5880, A2 => n7848, ZN => n477);
   U3547 : AOI22_X1 port map( A1 => n6903, A2 => n477, B1 => n7738, B2 => n7849
                           , ZN => n7850);
   U3548 : AOI21_X1 port map( B1 => n6914, B2 => n7850, A => n5388, ZN => n7694
                           );
   U3549 : INV_X1 port map( A => n7319, ZN => IRAM_ADDRESS_0_port);
   U3550 : AOI22_X1 port map( A1 => n7205, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n7168, B2 
                           => n7182, ZN => n7851);
   U3551 : OAI21_X1 port map( B1 => n7107, B2 => n6824, A => n7851, ZN => n5479
                           );
   U3552 : AOI22_X1 port map( A1 => n7275, A2 => IRAM_ADDRESS_0_port, B1 => 
                           n7197, B2 => n5479, ZN => n7852);
   U3553 : INV_X1 port map( A => n7852, ZN => n7711);
   U3554 : OAI211_X1 port map( C1 => n6918, C2 => IRAM_ADDRESS_12_port, A => 
                           n6917, B => n7201, ZN => n7853);
   U3555 : NAND2_X1 port map( A1 => n6801, A2 => n7853, ZN => n7912);
   U3556 : INV_X1 port map( A => n7912, ZN => n7776);
   U3557 : AOI211_X1 port map( C1 => n6783, C2 => n6925, A => n7274, B => n6918
                           , ZN => n7854);
   U3558 : NOR2_X1 port map( A1 => n6818, A2 => n7854, ZN => n4128);
   U3559 : AOI22_X1 port map( A1 => n7109, A2 => n7120, B1 => n7205, B2 => 
                           datapath_i_alu_output_val_i_11_port, ZN => n7855);
   U3560 : OAI21_X1 port map( B1 => n4128, B2 => n8071, A => n7855, ZN => n7713
                           );
   U3561 : AOI211_X1 port map( C1 => n6917, C2 => n6784, A => n6916, B => n7274
                           , ZN => n7856);
   U3562 : NOR2_X1 port map( A1 => n6817, A2 => n7856, ZN => n7714);
   U3563 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n7109, B2
                           => n7123, ZN => n7857);
   U3564 : OAI21_X1 port map( B1 => n7714, B2 => n8071, A => n7857, ZN => n7715
                           );
   U3565 : NOR2_X1 port map( A1 => n7709, A2 => cu_i_n135, ZN => n7859);
   U3566 : NOR2_X1 port map( A1 => n7859, A2 => n7858, ZN => n7708);
   U3567 : AOI211_X1 port map( C1 => n6756, C2 => n7861, A => n7274, B => n7860
                           , ZN => n7862);
   U3568 : NOR2_X1 port map( A1 => n6816, A2 => n7862, ZN => n7716);
   U3569 : AOI211_X1 port map( C1 => n6770, C2 => n7864, A => n7274, B => n7863
                           , ZN => n7865);
   U3570 : NOR2_X1 port map( A1 => n6809, A2 => n7865, ZN => n7728);
   U3571 : AOI211_X1 port map( C1 => n6768, C2 => n7867, A => n7274, B => n7866
                           , ZN => n7868);
   U3572 : NOR2_X1 port map( A1 => n6810, A2 => n7868, ZN => n7730);
   U3573 : AOI211_X1 port map( C1 => n6758, C2 => n7870, A => n7274, B => n7869
                           , ZN => n7871);
   U3574 : NOR2_X1 port map( A1 => n6815, A2 => n7871, ZN => n7722);
   U3575 : AOI211_X1 port map( C1 => n6760, C2 => n7873, A => n7274, B => n7872
                           , ZN => n7874);
   U3576 : NOR2_X1 port map( A1 => n6814, A2 => n7874, ZN => n7718);
   U3577 : AOI211_X1 port map( C1 => n6766, C2 => n7876, A => n7274, B => n7875
                           , ZN => n7877);
   U3578 : NOR2_X1 port map( A1 => n6811, A2 => n7877, ZN => n7726);
   U3579 : AOI211_X1 port map( C1 => n6764, C2 => n7879, A => n7274, B => n7878
                           , ZN => n7880);
   U3580 : NOR2_X1 port map( A1 => n6812, A2 => n7880, ZN => n7724);
   U3581 : AOI211_X1 port map( C1 => n6762, C2 => n7882, A => n7274, B => n7881
                           , ZN => n7883);
   U3582 : NOR2_X1 port map( A1 => n6813, A2 => n7883, ZN => n7720);
   U3583 : MUX2_X1 port map( A => n6838, B => n6961, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U3584 : AOI22_X1 port map( A1 => n6937, A2 => cu_i_cmd_alu_op_type_0_port, 
                           B1 => n7095, B2 => n6941, ZN => n7890);
   U3585 : AOI22_X1 port map( A1 => n6937, A2 => cu_i_cmd_alu_op_type_1_port, 
                           B1 => n7095, B2 => n6940, ZN => n7889);
   U3586 : AOI21_X1 port map( B1 => n7887, B2 => n7889, A => n7886, ZN => n7884
                           );
   U3587 : AOI21_X1 port map( B1 => n7887, B2 => n7890, A => n7886, ZN => n7885
                           );
   U3588 : NOR2_X1 port map( A1 => n7889, A2 => n7885, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U3589 : INV_X1 port map( A => n7886, ZN => n7888);
   U3590 : OAI211_X1 port map( C1 => n7890, C2 => n7889, A => n7888, B => n7887
                           , ZN => n7891);
   U3591 : INV_X1 port map( A => n7891, ZN => n7700);
   U3592 : INV_X1 port map( A => datapath_i_alu_output_val_i_10_port, ZN => 
                           n7892);
   U3593 : OAI222_X1 port map( A1 => n7892, A2 => n7104, B1 => n7107, B2 => 
                           n7220, C1 => n7222, C2 => n7166, ZN => n1447);
   U3594 : NOR2_X1 port map( A1 => n7959, A2 => n7908, ZN => n7907);
   U3595 : NAND2_X1 port map( A1 => n7907, A2 => n1447, ZN => n6082);
   U3596 : OAI211_X1 port map( C1 => n7907, C2 => n1447, A => n7202, B => n6082
                           , ZN => n7893);
   U3597 : AND2_X1 port map( A1 => n6802, A2 => n7893, ZN => n7341);
   U3598 : CLKBUF_X1 port map( A => n8076, Z => n8079);
   U3599 : AOI211_X1 port map( C1 => n7957, C2 => n7939, A => n7275, B => n7894
                           , ZN => n7895);
   U3600 : OR2_X1 port map( A1 => n6821, A2 => n7895, ZN => n5507);
   U3601 : INV_X1 port map( A => curr_instruction_to_cu_i_19_port, ZN => n7898)
                           ;
   U3602 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_20_port, A2 => 
                           curr_instruction_to_cu_i_16_port, A3 => 
                           curr_instruction_to_cu_i_17_port, A4 => n7756, ZN =>
                           n7897);
   U3603 : AOI21_X1 port map( B1 => n7898, B2 => n7897, A => n7896, ZN => n7899
                           );
   U3604 : AOI21_X1 port map( B1 => n7901, B2 => n7900, A => n7899, ZN => n7905
                           );
   U3605 : OR4_X1 port map( A1 => n5071, A2 => n5065, A3 => n7752, A4 => n5067,
                           ZN => n7902);
   U3606 : OAI21_X1 port map( B1 => n5069, B2 => n7902, A => n7738, ZN => n7903
                           );
   U3607 : OAI211_X1 port map( C1 => n7905, C2 => n8067, A => n7904, B => n7903
                           , ZN => n7906);
   U3608 : AOI211_X1 port map( C1 => n6882, C2 => n7169, A => n7740, B => n7906
                           , ZN => n4052);
   U3609 : OR2_X1 port map( A1 => n4052, A2 => n7170, ZN => n7342);
   U3610 : AOI211_X1 port map( C1 => n7959, C2 => n7908, A => n7275, B => n7907
                           , ZN => n7909);
   U3611 : OR2_X1 port map( A1 => n6819, A2 => n7909, ZN => n5506);
   U3612 : OR2_X1 port map( A1 => n7248, A2 => n7151, ZN => cu_i_N278);
   U3613 : INV_X1 port map( A => n7313, ZN => IRAM_ADDRESS_14_port);
   U3614 : INV_X1 port map( A => n7314, ZN => IRAM_ADDRESS_16_port);
   U3615 : INV_X1 port map( A => n7315, ZN => IRAM_ADDRESS_18_port);
   U3616 : INV_X1 port map( A => n7316, ZN => IRAM_ADDRESS_20_port);
   U3617 : INV_X1 port map( A => n7317, ZN => IRAM_ADDRESS_22_port);
   U3618 : INV_X1 port map( A => n7309, ZN => IRAM_ADDRESS_24_port);
   U3619 : INV_X1 port map( A => n7307, ZN => IRAM_ADDRESS_26_port);
   U3620 : INV_X1 port map( A => n7310, ZN => IRAM_ADDRESS_28_port);
   U3621 : INV_X1 port map( A => n7318, ZN => IRAM_ADDRESS_30_port);
   U3622 : INV_X1 port map( A => n7708, ZN => n8050);
   U3623 : NOR2_X1 port map( A1 => n7249, A2 => n8050, ZN => n5097);
   U3624 : INV_X1 port map( A => n4128, ZN => n7910);
   U3625 : AOI22_X1 port map( A1 => n6919, A2 => n7910, B1 => n6834, B2 => 
                           n7053, ZN => n7911);
   U3626 : OAI21_X1 port map( B1 => n6920, B2 => n7118, A => n7911, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U3627 : AOI22_X1 port map( A1 => n6919, A2 => n7912, B1 => n6834, B2 => 
                           n7055, ZN => n7913);
   U3628 : OAI21_X1 port map( B1 => n6920, B2 => n7216, A => n7913, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U3629 : INV_X1 port map( A => n7714, ZN => n7914);
   U3630 : AOI22_X1 port map( A1 => n6919, A2 => n7914, B1 => n6834, B2 => 
                           n7057, ZN => n7915);
   U3631 : OAI21_X1 port map( B1 => n6920, B2 => n7121, A => n7915, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U3632 : MUX2_X1 port map( A => n6842, B => n6949, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U3633 : MUX2_X1 port map( A => n6840, B => n6955, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U3634 : MUX2_X1 port map( A => n6841, B => n6952, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U3635 : NAND2_X1 port map( A1 => n7708, A2 => n7249, ZN => n5098);
   U3636 : AOI22_X1 port map( A1 => n6919, A2 => n6924, B1 => n6834, B2 => 
                           n7051, ZN => n7916);
   U3637 : OAI21_X1 port map( B1 => n6920, B2 => n7220, A => n7916, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U3638 : MUX2_X1 port map( A => IRAM_DATA(22), B => n6902, S => n6937, Z => 
                           n5047);
   U3639 : MUX2_X1 port map( A => n6848, B => n6946, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U3640 : AOI22_X1 port map( A1 => n6919, A2 => n7917, B1 => n6834, B2 => 
                           n7059, ZN => n7918);
   U3641 : OAI21_X1 port map( B1 => n6920, B2 => n7218, A => n7918, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U3642 : INV_X1 port map( A => n7716, ZN => n7919);
   U3643 : AOI22_X1 port map( A1 => n6919, A2 => n7919, B1 => n6834, B2 => 
                           n7061, ZN => n7920);
   U3644 : OAI21_X1 port map( B1 => n6920, B2 => n7124, A => n7920, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U3645 : INV_X1 port map( A => n7718, ZN => n7921);
   U3646 : AOI22_X1 port map( A1 => n6919, A2 => n7921, B1 => n6834, B2 => 
                           n7069, ZN => n7922);
   U3647 : OAI21_X1 port map( B1 => n6920, B2 => n7130, A => n7922, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U3648 : INV_X1 port map( A => n7713, ZN => n7960);
   U3649 : NOR2_X1 port map( A1 => n7960, A2 => n6082, ZN => n6081);
   U3650 : INV_X1 port map( A => datapath_i_alu_output_val_i_12_port, ZN => 
                           n7923);
   U3651 : OAI222_X1 port map( A1 => n7923, A2 => n7104, B1 => n7107, B2 => 
                           n7216, C1 => n7776, C2 => n7166, ZN => n1445);
   U3652 : NAND2_X1 port map( A1 => n6081, A2 => n1445, ZN => n4231);
   U3653 : INV_X1 port map( A => n7715, ZN => n7924);
   U3654 : NOR2_X1 port map( A1 => n7924, A2 => n4231, ZN => n5120);
   U3655 : INV_X1 port map( A => n7728, ZN => n7925);
   U3656 : AOI22_X1 port map( A1 => n6919, A2 => n7925, B1 => n6834, B2 => 
                           n7089, ZN => n7926);
   U3657 : OAI21_X1 port map( B1 => n6920, B2 => n7145, A => n7926, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U3658 : AOI22_X1 port map( A1 => n6919, A2 => n7927, B1 => n6834, B2 => 
                           n7091, ZN => n7928);
   U3659 : OAI21_X1 port map( B1 => n6920, B2 => n7238, A => n7928, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U3660 : AOI22_X1 port map( A1 => n6919, A2 => n7929, B1 => n6834, B2 => 
                           n7087, ZN => n7930);
   U3661 : OAI21_X1 port map( B1 => n6920, B2 => n7242, A => n7930, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U3662 : AOI22_X1 port map( A1 => n6919, A2 => n7931, B1 => n6834, B2 => 
                           n7083, ZN => n7932);
   U3663 : OAI21_X1 port map( B1 => n6920, B2 => n7244, A => n7932, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U3664 : INV_X1 port map( A => n7726, ZN => n7933);
   U3665 : AOI22_X1 port map( A1 => n6919, A2 => n7933, B1 => n6834, B2 => 
                           n7081, ZN => n7934);
   U3666 : OAI21_X1 port map( B1 => n6920, B2 => n7139, A => n7934, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U3667 : AOI22_X1 port map( A1 => n6919, A2 => n7935, B1 => n6834, B2 => 
                           n7079, ZN => n7936);
   U3668 : OAI21_X1 port map( B1 => n6920, B2 => n7246, A => n7936, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U3669 : AOI22_X1 port map( A1 => n6919, A2 => n7937, B1 => n6834, B2 => 
                           n7067, ZN => n7938);
   U3670 : OAI211_X1 port map( C1 => n7940, C2 => n1453, A => n7202, B => n7939
                           , ZN => n7941);
   U3671 : NAND2_X1 port map( A1 => n6804, A2 => n7941, ZN => n6096);
   U3672 : AOI22_X1 port map( A1 => n5097, A2 => n6096, B1 => n7047, B2 => 
                           n8050, ZN => n7942);
   U3673 : OAI21_X1 port map( B1 => n7227, B2 => n5098, A => n7942, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);
   U3674 : AOI22_X1 port map( A1 => n5097, A2 => n5507, B1 => n7048, B2 => 
                           n8050, ZN => n7943);
   U3675 : OAI21_X1 port map( B1 => n7113, B2 => n5098, A => n7943, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U3676 : AOI22_X1 port map( A1 => n5097, A2 => n5506, B1 => n7050, B2 => 
                           n8050, ZN => n4989);
   U3677 : AOI22_X1 port map( A1 => n6919, A2 => n7944, B1 => n6834, B2 => 
                           n7063, ZN => n7945);
   U3678 : OAI21_X1 port map( B1 => n6920, B2 => n7261, A => n7945, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U3679 : NOR2_X1 port map( A1 => n8077, A2 => n7364, ZN => n7982);
   U3680 : INV_X1 port map( A => n7982, ZN => n7984);
   U3681 : NOR2_X1 port map( A1 => n7365, A2 => n7984, ZN => n7983);
   U3682 : NOR2_X1 port map( A1 => n7983, A2 => n7366, ZN => n7946);
   U3683 : AOI211_X1 port map( C1 => n7983, C2 => n7366, A => n6928, B => n7946
                           , ZN => cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U3685 : AOI22_X1 port map( A1 => n5097, A2 => n7947, B1 => n7049, B2 => 
                           n8050, ZN => n7948);
   U3686 : OAI21_X1 port map( B1 => n7224, B2 => n5098, A => n7948, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U3687 : AOI22_X1 port map( A1 => n5097, A2 => n7712, B1 => n7042, B2 => 
                           n8050, ZN => n7949);
   U3688 : OAI21_X1 port map( B1 => n6828, B2 => n5098, A => n7949, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U3689 : AOI22_X1 port map( A1 => n5097, A2 => n7334, B1 => n7046, B2 => 
                           n8050, ZN => n7950);
   U3690 : OAI21_X1 port map( B1 => n7196, B2 => n5098, A => n7950, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U3691 : AOI22_X1 port map( A1 => n6919, A2 => n7951, B1 => n6834, B2 => 
                           n7071, ZN => n7952);
   U3692 : OAI21_X1 port map( B1 => n6920, B2 => n7255, A => n7952, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U3693 : OAI211_X1 port map( C1 => n7954, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n7202, B => n7953, ZN => n7955);
   U3694 : NAND2_X1 port map( A1 => n6805, A2 => n7955, ZN => n6113);
   U3695 : AOI22_X1 port map( A1 => n5097, A2 => n6113, B1 => n7045, B2 => 
                           n8050, ZN => n7956);
   U3696 : OAI21_X1 port map( B1 => n7230, B2 => n5098, A => n7956, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U3697 : NAND2_X1 port map( A1 => n4052, A2 => n7170, ZN => n5092);
   U3698 : INV_X1 port map( A => n7694, ZN => n8045);
   U3699 : NOR2_X1 port map( A1 => n8048, A2 => n8045, ZN => n7994);
   U3700 : NAND2_X1 port map( A1 => n7994, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n7993);
   U3701 : NOR2_X1 port map( A1 => n7958, A2 => n7993, ZN => n7996);
   U3702 : NAND2_X1 port map( A1 => n7996, A2 => n1453, ZN => n7995);
   U3703 : NOR2_X1 port map( A1 => n7957, A2 => n7995, ZN => n7998);
   U3704 : AOI211_X1 port map( C1 => n7957, C2 => n7995, A => n7998, B => n7704
                           , ZN => n4987);
   U3705 : AOI211_X1 port map( C1 => n7958, C2 => n7993, A => n7996, B => n7704
                           , ZN => n4986);
   U3706 : NAND2_X1 port map( A1 => n7998, A2 => n1449, ZN => n7997);
   U3707 : NOR2_X1 port map( A1 => n7959, A2 => n7997, ZN => n7999);
   U3708 : AOI211_X1 port map( C1 => n7959, C2 => n7997, A => n7999, B => n7704
                           , ZN => n4985);
   U3709 : AOI211_X1 port map( C1 => n6913, C2 => n6783, A => n6911, B => n7277
                           , ZN => n4984);
   U3710 : NAND2_X1 port map( A1 => n7999, A2 => n1447, ZN => n6157);
   U3711 : NOR2_X1 port map( A1 => n7960, A2 => n6157, ZN => n6159);
   U3712 : NAND2_X1 port map( A1 => n6159, A2 => n1445, ZN => n4341);
   U3713 : NOR2_X1 port map( A1 => n6910, A2 => n6785, ZN => n8001);
   U3714 : AOI211_X1 port map( C1 => n6785, C2 => n6910, A => n8001, B => n7202
                           , ZN => n4983);
   U3715 : NAND2_X1 port map( A1 => n6781, A2 => n8001, ZN => n8000);
   U3716 : NOR2_X1 port map( A1 => n6757, A2 => n8000, ZN => n8003);
   U3717 : AOI211_X1 port map( C1 => n6757, C2 => n8000, A => n8003, B => n7202
                           , ZN => n4982);
   U3718 : NAND2_X1 port map( A1 => n6780, A2 => n8003, ZN => n8002);
   U3719 : NOR2_X1 port map( A1 => n6759, A2 => n8002, ZN => n8005);
   U3720 : AOI211_X1 port map( C1 => n6759, C2 => n8002, A => n8005, B => n7202
                           , ZN => n4981);
   U3721 : NAND2_X1 port map( A1 => n6779, A2 => n8005, ZN => n8004);
   U3722 : NOR2_X1 port map( A1 => n6761, A2 => n8004, ZN => n8007);
   U3723 : AOI211_X1 port map( C1 => n6761, C2 => n8004, A => n8007, B => n7202
                           , ZN => n4980);
   U3724 : NAND2_X1 port map( A1 => n6778, A2 => n8007, ZN => n8006);
   U3725 : NOR2_X1 port map( A1 => n6763, A2 => n8006, ZN => n8009);
   U3726 : AOI211_X1 port map( C1 => n6763, C2 => n8006, A => n8009, B => n7202
                           , ZN => n4979);
   U3727 : NAND2_X1 port map( A1 => n6777, A2 => n8009, ZN => n8008);
   U3728 : NOR2_X1 port map( A1 => n6765, A2 => n8008, ZN => n8011);
   U3729 : AOI211_X1 port map( C1 => n6765, C2 => n8008, A => n8011, B => n7202
                           , ZN => n4978);
   U3730 : NAND2_X1 port map( A1 => n6776, A2 => n8011, ZN => n8010);
   U3731 : NOR2_X1 port map( A1 => n6767, A2 => n8010, ZN => n8013);
   U3732 : AOI211_X1 port map( C1 => n6767, C2 => n8010, A => n8013, B => n7202
                           , ZN => n4977);
   U3733 : NAND2_X1 port map( A1 => n6775, A2 => n8013, ZN => n8012);
   U3734 : NOR2_X1 port map( A1 => n6769, A2 => n8012, ZN => n8015);
   U3735 : AOI211_X1 port map( C1 => n6769, C2 => n8012, A => n8015, B => n7202
                           , ZN => n4976);
   U3736 : NAND2_X1 port map( A1 => n6774, A2 => n8015, ZN => n8014);
   U3737 : NOR2_X1 port map( A1 => n6771, A2 => n8014, ZN => n8016);
   U3738 : AOI211_X1 port map( C1 => n6771, C2 => n8014, A => n8016, B => n7202
                           , ZN => n4975);
   U3739 : AOI22_X1 port map( A1 => n5388, A2 => n8082, B1 => n7248, B2 => 
                           n7709, ZN => n4974);
   U3740 : INV_X1 port map( A => datapath_i_alu_output_val_i_31_port, ZN => 
                           n7961);
   U3741 : OAI222_X1 port map( A1 => n7732, A2 => n7166, B1 => n7961, B2 => 
                           n7104, C1 => n7240, C2 => n7107, ZN => n5542);
   U3742 : NAND3_X1 port map( A1 => n7257, A2 => n6832, A3 => n8078, ZN => 
                           n7962);
   U3743 : NOR2_X1 port map( A1 => n6898, A2 => n7962, ZN => n7977);
   U3744 : NOR2_X1 port map( A1 => n7098, A2 => n7363, ZN => n7974);
   U3745 : NAND2_X1 port map( A1 => n6832, A2 => n6909, ZN => n7969);
   U3746 : INV_X1 port map( A => n7962, ZN => n7963);
   U3747 : NAND3_X1 port map( A1 => n6898, A2 => n7097, A3 => n7963, ZN => 
                           n7981);
   U3748 : INV_X1 port map( A => n7977, ZN => n7964);
   U3749 : OAI211_X1 port map( C1 => n7097, C2 => n7969, A => n7981, B => n7964
                           , ZN => n7965);
   U3750 : AOI22_X1 port map( A1 => n7977, A2 => n6932, B1 => n7974, B2 => 
                           n7965, ZN => n7968);
   U3751 : NAND3_X1 port map( A1 => n7265, A2 => n6934, A3 => n6901, ZN => 
                           n7967);
   U3752 : NAND2_X1 port map( A1 => n7264, A2 => n6896, ZN => n7966);
   U3753 : NAND4_X1 port map( A1 => n6790, A2 => n7968, A3 => n7967, A4 => 
                           n7966, ZN => cu_i_N264);
   U3754 : NOR2_X1 port map( A1 => n7969, A2 => n7257, ZN => n7970);
   U3755 : AOI21_X1 port map( B1 => n7970, B2 => n7974, A => n6896, ZN => n7979
                           );
   U3756 : NOR3_X1 port map( A1 => n6831, A2 => n6899, A3 => n7981, ZN => n7973
                           );
   U3757 : NAND3_X1 port map( A1 => n7265, A2 => n7339, A3 => n7099, ZN => 
                           n7971);
   U3758 : NAND2_X1 port map( A1 => n7971, A2 => n6927, ZN => n7972);
   U3759 : AOI211_X1 port map( C1 => n6934, C2 => n7367, A => n7973, B => n7972
                           , ZN => n7976);
   U3760 : NAND3_X1 port map( A1 => n7097, A2 => n7977, A3 => n7974, ZN => 
                           n7975);
   U3761 : NAND3_X1 port map( A1 => n7979, A2 => n7976, A3 => n7975, ZN => 
                           cu_i_N265);
   U3762 : OAI221_X1 port map( B1 => n6932, B2 => n7097, C1 => n6932, C2 => 
                           n7363, A => n7977, ZN => n7980);
   U3763 : OAI221_X1 port map( B1 => n7339, B2 => n7264, C1 => n7339, C2 => 
                           n7100, A => n7367, ZN => n7978);
   U3764 : OAI211_X1 port map( C1 => n7098, C2 => n7980, A => n7979, B => n7978
                           , ZN => cu_i_N266);
   U3765 : OAI221_X1 port map( B1 => n7981, B2 => n6831, C1 => n7981, C2 => 
                           n7098, A => n7369, ZN => cu_i_N267);
   U3766 : NAND2_X1 port map( A1 => n6937, A2 => n6928, ZN => cu_i_N274);
   U3767 : AOI211_X1 port map( C1 => n7364, C2 => n8077, A => n6928, B => n7982
                           , ZN => cu_i_N275);
   U3768 : NOR2_X1 port map( A1 => n6928, A2 => n6942, ZN => cu_i_N273);
   U3769 : AOI211_X1 port map( C1 => n7365, C2 => n7984, A => n6928, B => n7983
                           , ZN => cu_i_N276);
   U3770 : AOI211_X1 port map( C1 => n6937, C2 => n6894, A => n6928, B => n6931
                           , ZN => cu_i_N279);
   U3771 : NOR2_X1 port map( A1 => n7748, A2 => n7736, ZN => n5089);
   U3772 : NOR2_X1 port map( A1 => n5076, A2 => n5077, ZN => n492);
   U3773 : NAND4_X1 port map( A1 => n7749, A2 => n5089, A3 => n492, A4 => n7735
                           , ZN => n7990);
   U3774 : NOR2_X1 port map( A1 => n7986, A2 => n7985, ZN => n8053);
   U3775 : NAND3_X1 port map( A1 => n6903, A2 => n7987, A3 => n8053, ZN => 
                           n7988);
   U3776 : OAI21_X1 port map( B1 => n7990, B2 => n7989, A => n7988, ZN => 
                           cu_i_cmd_word_8_port);
   U3777 : MUX2_X1 port map( A => n6807, B => cu_i_cmd_word_8_port, S => n5388,
                           Z => alu_cin_i);
   U3778 : MUX2_X1 port map( A => n6936, B => n6879, S => n5388, Z => n5053);
   U3779 : MUX2_X1 port map( A => n7150, B => n6878, S => n5388, Z => n5052);
   U3780 : MUX2_X1 port map( A => n6788, B => n6877, S => n5388, Z => n5051);
   U3781 : MUX2_X1 port map( A => IRAM_DATA(25), B => n6876, S => n7200, Z => 
                           n5049);
   U3782 : MUX2_X1 port map( A => IRAM_DATA(24), B => n6875, S => n7200, Z => 
                           n5048);
   U3783 : MUX2_X1 port map( A => IRAM_DATA(21), B => n6874, S => n6937, Z => 
                           n5046);
   U3784 : MUX2_X1 port map( A => IRAM_DATA(10), B => n6873, S => n7200, Z => 
                           n5045);
   U3785 : MUX2_X1 port map( A => IRAM_DATA(9), B => n6872, S => n7200, Z => 
                           n5044);
   U3786 : MUX2_X1 port map( A => IRAM_DATA(8), B => n6871, S => n7200, Z => 
                           n5043);
   U3787 : MUX2_X1 port map( A => IRAM_DATA(7), B => n6870, S => n7200, Z => 
                           n5042);
   U3788 : MUX2_X1 port map( A => IRAM_DATA(6), B => n6869, S => n7200, Z => 
                           n5041);
   U3789 : INV_X1 port map( A => n7763, ZN => n8046);
   U3790 : NOR2_X1 port map( A1 => n8046, A2 => n8045, ZN => n7992);
   U3791 : INV_X1 port map( A => n7994, ZN => n7991);
   U3792 : OAI211_X1 port map( C1 => n7992, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n4337, B => n7991, ZN => n4972);
   U3793 : OAI211_X1 port map( C1 => n7994, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n4337, B => n7993, ZN => n4971);
   U3794 : OAI211_X1 port map( C1 => n7996, C2 => n1453, A => n4337, B => n7995
                           , ZN => n4970);
   U3795 : OAI211_X1 port map( C1 => n7998, C2 => n1449, A => n4337, B => n7997
                           , ZN => n4969);
   U3796 : OAI211_X1 port map( C1 => n7999, C2 => n1447, A => n4337, B => n6157
                           , ZN => n4968);
   U3797 : OAI211_X1 port map( C1 => n6912, C2 => IRAM_ADDRESS_12_port, A => 
                           n7275, B => n6910, ZN => n4966);
   U3798 : OAI211_X1 port map( C1 => n8001, C2 => IRAM_ADDRESS_14_port, A => 
                           n7275, B => n8000, ZN => n4965);
   U3799 : OAI211_X1 port map( C1 => n8003, C2 => IRAM_ADDRESS_16_port, A => 
                           n7275, B => n8002, ZN => n4964);
   U3800 : OAI211_X1 port map( C1 => n8005, C2 => IRAM_ADDRESS_18_port, A => 
                           n7275, B => n8004, ZN => n4963);
   U3801 : OAI211_X1 port map( C1 => n8007, C2 => IRAM_ADDRESS_20_port, A => 
                           n7275, B => n8006, ZN => n4962);
   U3802 : OAI211_X1 port map( C1 => n8009, C2 => IRAM_ADDRESS_22_port, A => 
                           n7275, B => n8008, ZN => n4961);
   U3803 : OAI211_X1 port map( C1 => n8011, C2 => IRAM_ADDRESS_24_port, A => 
                           n7275, B => n8010, ZN => n4960);
   U3804 : OAI211_X1 port map( C1 => n8013, C2 => IRAM_ADDRESS_26_port, A => 
                           n7275, B => n8012, ZN => n4959);
   U3805 : OAI211_X1 port map( C1 => n8015, C2 => IRAM_ADDRESS_28_port, A => 
                           n7275, B => n8014, ZN => n4958);
   U3806 : NAND2_X1 port map( A1 => n6773, A2 => n8016, ZN => n8017);
   U3807 : OAI211_X1 port map( C1 => n8016, C2 => IRAM_ADDRESS_30_port, A => 
                           n7275, B => n8017, ZN => n4957);
   U3808 : XOR2_X1 port map( A => n6772, B => n8017, Z => n5085);
   U3809 : AND2_X1 port map( A1 => n7248, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U3810 : OAI21_X1 port map( B1 => n8020, B2 => n8019, A => n8018, ZN => 
                           read_rf_p2_i);
   U3811 : OAI21_X1 port map( B1 => n6825, B2 => n7270, A => n7558, ZN => 
                           datapath_i_decode_stage_dp_n44);
   U3812 : OAI21_X1 port map( B1 => n6828, B2 => n7270, A => n7555, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U3813 : OAI21_X1 port map( B1 => n7236, B2 => n7270, A => n7554, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U3814 : OAI21_X1 port map( B1 => n7233, B2 => n7270, A => n7553, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U3815 : OAI21_X1 port map( B1 => n7230, B2 => n7270, A => n7552, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U3816 : OAI21_X1 port map( B1 => n7270, B2 => n7112, A => n7551, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U3817 : OAI21_X1 port map( B1 => n7227, B2 => n7270, A => n7550, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U3818 : OAI21_X1 port map( B1 => n7270, B2 => n7153, A => n7549, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U3819 : OAI21_X1 port map( B1 => n7224, B2 => n7270, A => n7548, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U3820 : OAI21_X1 port map( B1 => n7199, B2 => n7152, A => n7547, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U3821 : OAI21_X1 port map( B1 => n7199, B2 => n7221, A => n7546, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U3822 : OAI21_X1 port map( B1 => n7270, B2 => n7163, A => n7545, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U3823 : OAI21_X1 port map( B1 => n7270, B2 => n7217, A => n7544, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U3824 : OAI21_X1 port map( B1 => n7199, B2 => n7162, A => n7543, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U3825 : OAI21_X1 port map( B1 => n7199, B2 => n7219, A => n7542, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U3826 : OAI21_X1 port map( B1 => n7270, B2 => n7161, A => n7541, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U3827 : OAI21_X1 port map( B1 => n7270, B2 => n7262, A => n7540, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U3828 : OAI21_X1 port map( B1 => n7199, B2 => n7160, A => n7539, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U3829 : OAI21_X1 port map( B1 => n7199, B2 => n7260, A => n7538, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U3830 : OAI21_X1 port map( B1 => n7270, B2 => n7159, A => n7537, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U3831 : OAI21_X1 port map( B1 => n7270, B2 => n7256, A => n7536, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U3832 : OAI21_X1 port map( B1 => n7199, B2 => n7158, A => n7535, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U3833 : OAI21_X1 port map( B1 => n7199, B2 => n7253, A => n7534, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U3834 : OAI21_X1 port map( B1 => n7270, B2 => n7157, A => n7533, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U3835 : OAI21_X1 port map( B1 => n7270, B2 => n7247, A => n7532, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U3836 : OAI21_X1 port map( B1 => n7199, B2 => n7156, A => n7531, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U3837 : OAI21_X1 port map( B1 => n7199, B2 => n7245, A => n7530, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U3838 : OAI21_X1 port map( B1 => n7270, B2 => n7155, A => n7529, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U3839 : OAI21_X1 port map( B1 => n7270, B2 => n7243, A => n7528, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U3840 : OAI21_X1 port map( B1 => n7199, B2 => n7154, A => n7527, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U3841 : OAI21_X1 port map( B1 => n7199, B2 => n7239, A => n7526, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U3842 : OAI21_X1 port map( B1 => n7270, B2 => n7241, A => n7525, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U3843 : NOR4_X1 port map( A1 => n1641, A2 => n1643, A3 => n1645, A4 => n1647
                           , ZN => n8024);
   U3844 : NOR4_X1 port map( A1 => n1649, A2 => n1651, A3 => n1653, A4 => n1655
                           , ZN => n8023);
   U3845 : NOR4_X1 port map( A1 => n1625, A2 => n1627, A3 => n1629, A4 => n1631
                           , ZN => n8022);
   U3846 : NOR4_X1 port map( A1 => n1633, A2 => n1635, A3 => n1637, A4 => n1639
                           , ZN => n8021);
   U3847 : NAND4_X1 port map( A1 => n8024, A2 => n8023, A3 => n8022, A4 => 
                           n8021, ZN => n8030);
   U3848 : NOR4_X1 port map( A1 => n1663, A2 => n1617, A3 => n1619, A4 => n1621
                           , ZN => n8028);
   U3849 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1661
                           , ZN => n8027);
   U3850 : NOR4_X1 port map( A1 => n1667, A2 => n1669, A3 => n1657, A4 => n1659
                           , ZN => n8026);
   U3851 : NOR4_X1 port map( A1 => n1623, A2 => n1671, A3 => n1673, A4 => n1665
                           , ZN => n8025);
   U3852 : NAND4_X1 port map( A1 => n8028, A2 => n8027, A3 => n8026, A4 => 
                           n8025, ZN => n8029);
   U3853 : NOR2_X1 port map( A1 => n8030, A2 => n8029, ZN => n5084);
   U3854 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n8080, Z => n5040);
   U3855 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n8080, Z => n5039);
   U3856 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n7250, Z => n5038);
   U3857 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n7250, Z => n5037);
   U3858 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n8080, Z => n5036);
   U3859 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n8080, Z => n5035);
   U3860 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n7250, Z => n5034);
   U3861 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n7250, Z => n5033);
   U3862 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, S 
                           => n8080, Z => n5032);
   U3863 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, S 
                           => n8080, Z => n5031);
   U3864 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, S 
                           => n7250, Z => n5030);
   U3865 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, S 
                           => n7250, Z => n5029);
   U3866 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, S 
                           => n8080, Z => n5028);
   U3867 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, S 
                           => n8080, Z => n5027);
   U3868 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, S 
                           => n7250, Z => n5026);
   U3869 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, S 
                           => n7250, Z => n5025);
   U3870 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, S 
                           => n8080, Z => n5024);
   U3871 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, S 
                           => n8080, Z => n5023);
   U3872 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, S 
                           => n7250, Z => n5022);
   U3873 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, S 
                           => n7250, Z => n5021);
   U3874 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n8080, Z => n5020);
   U3875 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, S 
                           => n8080, Z => n5019);
   U3876 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, S 
                           => n7250, Z => n5018);
   U3877 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, S 
                           => n7250, Z => n5017);
   U3878 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, S 
                           => n8080, Z => n5016);
   U3879 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, S 
                           => n8080, Z => n5015);
   U3880 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n7250, Z => n5014);
   U3881 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n8080, Z => n5013);
   U3882 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n8080, Z => n5012);
   U3883 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n8080, Z => n5011);
   U3884 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n8080, Z => n5010);
   U3885 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n8080, Z => n5009);
   U3886 : MUX2_X1 port map( A => n6868, B => n6967, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U3887 : MUX2_X1 port map( A => n6867, B => n6970, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U3888 : MUX2_X1 port map( A => n6866, B => n6973, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U3889 : MUX2_X1 port map( A => n6865, B => n6976, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U3890 : MUX2_X1 port map( A => n6864, B => n6979, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U3891 : MUX2_X1 port map( A => n6863, B => n6982, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U3892 : MUX2_X1 port map( A => n6862, B => n6985, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U3893 : MUX2_X1 port map( A => n6861, B => n6988, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U3894 : MUX2_X1 port map( A => n6860, B => n6991, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U3895 : MUX2_X1 port map( A => n6859, B => n6994, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U3896 : MUX2_X1 port map( A => n6858, B => n6997, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U3897 : MUX2_X1 port map( A => n6857, B => n7000, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U3898 : MUX2_X1 port map( A => n6856, B => n7003, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U3899 : MUX2_X1 port map( A => n6855, B => n7006, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U3900 : MUX2_X1 port map( A => n6854, B => n7009, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U3901 : MUX2_X1 port map( A => n6853, B => n7012, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U3902 : MUX2_X1 port map( A => n6852, B => n7015, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U3903 : MUX2_X1 port map( A => n6851, B => n7018, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U3904 : MUX2_X1 port map( A => n6850, B => n7021, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U3905 : MUX2_X1 port map( A => n6849, B => n7024, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U3906 : MUX2_X1 port map( A => n6847, B => n7027, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U3907 : MUX2_X1 port map( A => n6846, B => n7030, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U3908 : MUX2_X1 port map( A => n6845, B => n7033, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U3909 : MUX2_X1 port map( A => n6844, B => n7036, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U3910 : MUX2_X1 port map( A => n6843, B => n7039, S => n6808, Z => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U3911 : MUX2_X1 port map( A => n6837, B => n6964, S => n8031, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U3912 : INV_X1 port map( A => n7722, ZN => n8032);
   U3913 : AOI22_X1 port map( A1 => n6919, A2 => n8032, B1 => n6834, B2 => 
                           n7065, ZN => n8033);
   U3914 : OAI21_X1 port map( B1 => n6920, B2 => n7127, A => n8033, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U3915 : INV_X1 port map( A => n7720, ZN => n8034);
   U3916 : AOI22_X1 port map( A1 => n6919, A2 => n8034, B1 => n6834, B2 => 
                           n7073, ZN => n8035);
   U3917 : OAI21_X1 port map( B1 => n6920, B2 => n7133, A => n8035, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U3918 : AOI22_X1 port map( A1 => n6919, A2 => n8036, B1 => n6834, B2 => 
                           n7075, ZN => n8037);
   U3919 : OAI21_X1 port map( B1 => n6920, B2 => n7252, A => n8037, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U3920 : INV_X1 port map( A => n7724, ZN => n8038);
   U3921 : AOI22_X1 port map( A1 => n6919, A2 => n8038, B1 => n6834, B2 => 
                           n7077, ZN => n8039);
   U3922 : OAI21_X1 port map( B1 => n6920, B2 => n7136, A => n8039, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U3923 : AOI22_X1 port map( A1 => n5097, A2 => n7711, B1 => n7041, B2 => 
                           n8050, ZN => n8040);
   U3924 : OAI21_X1 port map( B1 => n6825, B2 => n5098, A => n8040, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U3925 : INV_X1 port map( A => n7730, ZN => n8041);
   U3926 : AOI22_X1 port map( A1 => n6919, A2 => n8041, B1 => n6834, B2 => 
                           n7085, ZN => n8042);
   U3927 : OAI21_X1 port map( B1 => n6920, B2 => n7142, A => n8042, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U3928 : AOI22_X1 port map( A1 => n8043, A2 => n6919, B1 => n6834, B2 => 
                           n7093, ZN => n8044);
   U3929 : OAI21_X1 port map( B1 => n7240, B2 => n6920, A => n8044, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U3930 : AOI22_X1 port map( A1 => n8046, A2 => n7694, B1 => n8045, B2 => 
                           n7763, ZN => n4956);
   U3931 : AOI22_X1 port map( A1 => n6791, A2 => n7275, B1 => n7202, B2 => 
                           n7763, ZN => n6207);
   U3932 : AOI22_X1 port map( A1 => n6207, A2 => n5097, B1 => n7043, B2 => 
                           n8050, ZN => n8047);
   U3933 : OAI21_X1 port map( B1 => n7236, B2 => n5098, A => n8047, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U3934 : OAI211_X1 port map( C1 => n7763, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n7202, B => n8048, ZN => n8049);
   U3935 : NAND2_X1 port map( A1 => n6806, A2 => n8049, ZN => n6209);
   U3936 : AOI22_X1 port map( A1 => n5097, A2 => n6209, B1 => n7044, B2 => 
                           n8050, ZN => n8051);
   U3937 : OAI21_X1 port map( B1 => n7233, B2 => n5098, A => n8051, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U3938 : MUX2_X1 port map( A => n6877, B => n6836, S => n5388, Z => n5006);
   U3939 : AND4_X1 port map( A1 => n7696, A2 => n7698, A3 => n4953, A4 => n7697
                           , ZN => n8052);
   U3940 : NAND2_X1 port map( A1 => n8052, A2 => n7695, ZN => n3596);
   U3941 : OAI21_X1 port map( B1 => n7741, B2 => n8054, A => n8053, ZN => n4954
                           );
   U3942 : MUX2_X1 port map( A => n6789, B => n6835, S => n5388, Z => n5285);
   U3943 : OAI221_X1 port map( B1 => n5388, B2 => n6883, C1 => n7709, C2 => 
                           cu_i_cmd_word_6_port, A => n6907, ZN => n8057);
   U3944 : AOI22_X1 port map( A1 => n5388, A2 => n8055, B1 => n6929, B2 => 
                           n7709, ZN => n8056);
   U3945 : MUX2_X1 port map( A => n6907, B => n8057, S => n8056, Z => n7702);
   U3946 : NAND2_X1 port map( A1 => n7702, A2 => n8072, ZN => n7333);
   U3947 : NAND2_X1 port map( A1 => n8075, A2 => n7702, ZN => n7335);
   U3948 : NOR2_X1 port map( A1 => n4052, A2 => n6923, ZN => n7347);
   U3949 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n7109, B2
                           => n7144, ZN => n8058);
   U3950 : OAI21_X1 port map( B1 => n7730, B2 => n8071, A => n8058, ZN => n7731
                           );
   U3951 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n7109, B2
                           => n7147, ZN => n8059);
   U3952 : OAI21_X1 port map( B1 => n7728, B2 => n8071, A => n8059, ZN => n7729
                           );
   U3953 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n7109, B2
                           => n7141, ZN => n8060);
   U3954 : OAI21_X1 port map( B1 => n7726, B2 => n8071, A => n8060, ZN => n7727
                           );
   U3955 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n7109, B2
                           => n7138, ZN => n8061);
   U3956 : OAI21_X1 port map( B1 => n7724, B2 => n8071, A => n8061, ZN => n7725
                           );
   U3957 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n7109, B2
                           => n7129, ZN => n8062);
   U3958 : OAI21_X1 port map( B1 => n7722, B2 => n8071, A => n8062, ZN => n7723
                           );
   U3959 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n7109, B2
                           => n7135, ZN => n8063);
   U3960 : OAI21_X1 port map( B1 => n7720, B2 => n8071, A => n8063, ZN => n7721
                           );
   U3961 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n7109, B2
                           => n7132, ZN => n8064);
   U3962 : OAI21_X1 port map( B1 => n7718, B2 => n8071, A => n8064, ZN => n7719
                           );
   U3963 : AOI22_X1 port map( A1 => n7203, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n7109, B2
                           => n7126, ZN => n8065);
   U3964 : OAI21_X1 port map( B1 => n7716, B2 => n8071, A => n8065, ZN => n7717
                           );
   U3965 : MUX2_X1 port map( A => n6933, B => n7181, S => n5388, Z => n7701);

end SYN_dlx_rtl;
