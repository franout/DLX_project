--------------------------------------------------------------------------------
-- Title       : write back stage of datapath 
-- Project     : DLX for Microelectronic Systems
--------------------------------------------------------------------------------
-- File        : a.b.e-Write_back.stage.vhd
-- Author      : Francesco Angione <s262620@studenti.polito.it> franout@github.com
-- Company     : Politecnico di Torino, Italy
-- Created     : Wed Jul 22 23:00:39 2020
-- Last update : Wed Jul 22 23:00:44 2020
-- Platform    : Default Part Number
-- Standard    : VHDL-2008 
--------------------------------------------------------------------------------
-- Copyright (c) 2020 Politecnico di Torino, Italy
-------------------------------------------------------------------------------
-- Description: 
--------------------------------------------------------------------------------


library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity write_back_stage is
  port (
	clock
  ) ;
end entity ; -- write_back_stage

architecture arch of write_back_stage is

begin

end architecture ; -- arch