
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n3076, 
      n3077, n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n1995, n1996, 
      n1997, n5121, n5122, n5123, n5124, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n1991, n1992, n7164, n7165, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n7170, n7171, n7172, 
      n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, 
      n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, 
      n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, 
      n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, 
      n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
      n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, 
      n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, 
      n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, 
      n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, 
      n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, 
      n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, 
      n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, 
      n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, 
      n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, 
      n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, 
      n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, 
      n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, 
      n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, 
      n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, 
      n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, 
      n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, 
      n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, 
      n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, 
      n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
      n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, 
      n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, 
      n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, 
      n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, 
      n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, 
      n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, 
      n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, 
      n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, 
      n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, 
      n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, 
      n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, 
      n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, 
      n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, 
      n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, 
      n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, 
      n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, 
      n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, 
      n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, 
      n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, 
      n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, 
      n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, 
      n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, 
      n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, 
      n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, 
      n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, 
      n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, 
      n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, 
      n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, 
      n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, 
      n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, 
      n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, 
      n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, 
      n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, 
      n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, 
      n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, 
      n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, 
      n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, 
      n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, 
      n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, 
      n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, 
      n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, 
      n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, 
      n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, 
      n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, 
      n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, 
      n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, 
      n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, 
      n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, 
      n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, 
      n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, 
      n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, 
      n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, 
      n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, 
      n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, 
      n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, 
      n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, 
      n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, 
      n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, 
      n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, 
      n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, 
      n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, 
      n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, 
      n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, 
      n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, 
      n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, 
      n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, 
      n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, 
      n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, 
      n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, 
      n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, 
      n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, 
      n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, 
      n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, 
      n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, 
      n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, 
      n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, 
      n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, 
      n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, 
      n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, 
      n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, 
      n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, 
      n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, 
      n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, 
      n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, 
      n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, 
      n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, 
      n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, 
      n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, 
      n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, 
      n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, 
      n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, 
      n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, 
      n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, 
      n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, 
      n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, 
      n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, 
      n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, 
      n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, 
      n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, 
      n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, 
      n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, 
      n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, 
      n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, 
      n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, 
      n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, 
      n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, 
      n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, 
      n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, 
      n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, 
      n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, 
      n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, 
      n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, 
      n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, 
      n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, 
      n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, 
      n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, 
      n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, 
      n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, 
      n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, 
      n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, 
      n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, 
      n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, 
      n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, 
      n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, 
      n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, 
      n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, 
      n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, 
      n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, 
      n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, 
      n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, 
      n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, 
      n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, 
      n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, 
      n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, 
      n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, 
      n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, 
      n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, 
      n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, 
      n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, 
      n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, 
      n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, 
      n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, 
      n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, 
      n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, 
      n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, 
      n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, 
      n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, 
      n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, 
      n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, 
      n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, 
      n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, 
      n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, 
      n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, 
      n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, 
      n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, 
      n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, 
      n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, 
      n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, 
      n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, 
      n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, 
      n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, 
      n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, 
      n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, 
      n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, 
      n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, 
      n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, 
      n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, 
      n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, 
      n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, 
      n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, 
      n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, 
      n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, 
      n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, 
      n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, 
      n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, 
      n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, 
      n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, 
      n9193, n9194, n9195, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348 : std_logic;

begin
   
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n1992, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n9190, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n1992, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n9190, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n9190, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n1992, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n1992, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n9190, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n9190, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n1992, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n9190, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n1992, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n9190, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n9190, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n1992, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n1992, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n9190, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n1992, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n9190, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n1992, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n9190, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n1992, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n1992, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n1992, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n1992, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n1992, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n1992, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n1992, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => n9195, GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => n9194, GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => n9193, GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => n9192, GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => n9191, GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => n7182, Q => n9189, QN => n7165);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => n7172, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => n7178, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => n7176, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => n7179, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3080);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => n7174, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => n7181, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => n7171, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => n7171, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => n7182, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => n7184, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => n7184, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3079);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => n7183, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => n7176, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => n7175, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => n7175, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => n7175, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => n7172, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3078);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => n7179, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => n7181, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => n7182, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => n7174, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => n7170, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => n7170, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => n7177, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => n7178, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => n7184, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3082);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => n7183, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => n7170, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => n7178, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => n7181, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => n7178, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => n7183, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => n7177, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => n7172, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => n7173, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => n7174, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => n7178, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => n7182, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3076);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => n7174, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => n7171, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => n7177, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => n7172, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => n7171, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => n7184, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => n7171, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => n7179, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => n7175, Q => n_1060, QN => n5126);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => n7181, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3095, CK => clk, RN => n7179, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => n7171, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => n7173, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => n7174, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => n7183, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => n7182, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => n7181, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => n7179, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => n7172, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => n7170, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => n7178, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => n7176, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n7182, Q => n_1106, QN => n5134);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => n7171, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => n7183, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => n7184, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => n7179, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => n7173, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => n7177, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => n7179, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => n7183, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1120);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => n7180, Q => n_1121, QN => n5133);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1122
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3094, CK => clk, RN => n7171, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1123
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => n7181, Q => boothmul_pipelined_i_sum_out_6_9_port
                           , QN => n_1124);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => n7174, Q => boothmul_pipelined_i_sum_out_6_8_port
                           , QN => n_1125);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => n7174, Q => boothmul_pipelined_i_sum_out_6_7_port
                           , QN => n_1126);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => n7176, Q => boothmul_pipelined_i_sum_out_6_6_port
                           , QN => n_1127);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => n7175, Q => boothmul_pipelined_i_sum_out_6_5_port
                           , QN => n_1128);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => n7179, Q => boothmul_pipelined_i_sum_out_6_4_port
                           , QN => n_1129);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => n7184, Q => boothmul_pipelined_i_sum_out_6_3_port
                           , QN => n_1130);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => n7180, Q => boothmul_pipelined_i_sum_out_6_2_port
                           , QN => n_1131);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => n7177, Q => boothmul_pipelined_i_sum_out_6_1_port
                           , QN => n_1132);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => n7172, Q => boothmul_pipelined_i_sum_out_6_0_port
                           , QN => n_1133);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => n5129
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => n5123
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1156);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1157);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1158);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1159);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1160);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1161);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1162);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1163);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1164);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => n7172, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1165);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => n7173, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1166);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1167);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => n7173, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => n7174, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => n7173, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => n7177, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => n7183, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1177);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => n7172, Q => n_1178, QN => n5132);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => n7179, Q => boothmul_pipelined_i_sum_out_5_9_port
                           , QN => n_1179);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3093, CK => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1180)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => n7182, Q => boothmul_pipelined_i_sum_out_5_7_port
                           , QN => n_1181);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => n7182, Q => boothmul_pipelined_i_sum_out_5_6_port
                           , QN => n_1182);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => n7177, Q => boothmul_pipelined_i_sum_out_5_5_port
                           , QN => n_1183);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => n7177, Q => boothmul_pipelined_i_sum_out_5_4_port
                           , QN => n_1184);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => n7171, Q => boothmul_pipelined_i_sum_out_5_3_port
                           , QN => n_1185);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => n7177, Q => boothmul_pipelined_i_sum_out_5_2_port
                           , QN => n_1186);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => n7175, Q => boothmul_pipelined_i_sum_out_5_1_port
                           , QN => n_1187);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => n7176, Q => boothmul_pipelined_i_sum_out_5_0_port
                           , QN => n_1188);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => n5128
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1189);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1190);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1191);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n5122);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => n7171, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => n7183, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => n7170, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => n7172, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => n7173, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1231);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => n7184, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1232
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => n7174, Q => n_1233, QN => n5131);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => n7175, Q => boothmul_pipelined_i_sum_out_4_7_port
                           , QN => n_1234);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3092, CK => clk, RN => n7170, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1235)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => n7177, Q => boothmul_pipelined_i_sum_out_4_5_port
                           , QN => n_1236);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => n7183, Q => boothmul_pipelined_i_sum_out_4_4_port
                           , QN => n_1237);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => n7183, Q => boothmul_pipelined_i_sum_out_4_3_port
                           , QN => n_1238);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => n7173, Q => boothmul_pipelined_i_sum_out_4_2_port
                           , QN => n_1239);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => n7177, Q => boothmul_pipelined_i_sum_out_4_1_port
                           , QN => n_1240);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => n7176, Q => boothmul_pipelined_i_sum_out_4_0_port
                           , QN => n_1241);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => n5127
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1242);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1243);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1244);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => n7175, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1245);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1246);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1249);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1250);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1251);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1252);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1253);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1254);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1255);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => n5121
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1256);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1257);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1258);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => n7179, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => n7182, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => n7174, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => n7177, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => n7176, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => n7184, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => n7180, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => n7174, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => n7170, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1282);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => n7170, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1283
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => n7174, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1284
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1285
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => rst_BAR, Q => n_1286, QN => n5124);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => n7176, Q => boothmul_pipelined_i_sum_out_3_5_port
                           , QN => n_1287);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3091, CK => clk, RN => n7179, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1288)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_3_port, QN => n_1289)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => n7181, Q => boothmul_pipelined_i_sum_out_3_2_port
                           , QN => n_1290);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => n7182, Q => boothmul_pipelined_i_sum_out_3_1_port
                           , QN => n_1291);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => n7176, Q => boothmul_pipelined_i_sum_out_3_0_port
                           , QN => n_1292);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => n7164
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1293);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1294);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1295);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1296);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1297);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => n7172, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1298);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => n7182, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => n7181, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => n7173, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => n7171, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => n7183, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => n7177, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => n7179, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => n7184, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => n7178, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => n7174, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => n7176, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => n7184, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => n7171, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => n7183, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => n7172, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => n7178, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => n7170, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => n7177, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => n7183, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1332
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => n7181, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1333
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => n7182, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1334
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1335
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => n7175, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1336
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => n7183, Q => n_1337, QN => n5130);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => n7173, Q => boothmul_pipelined_i_sum_out_2_3_port
                           , QN => n_1338);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3086, CK => clk, RN => n7173, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1339)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           n1981, CK => clk, RN => n7180, Q => 
                           boothmul_pipelined_i_sum_out_2_1_port, QN => n_1340)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => n7178, Q => boothmul_pipelined_i_sum_out_2_0_port
                           , QN => n_1341);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => n7170, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n3077);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n9190, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1982, B => n1983, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1980, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1979, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1977, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1975, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1973, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1971, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1969, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1967, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1965, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1963, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1961, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1959, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1957, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1955, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => n1978, 
                           CI => n3083, CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => n1976, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => n1974, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => n1972, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => n1970, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => n1968, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => n1966, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => n1964, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => n1962, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => n1960, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => n1958, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => n1956, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1342, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3085,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1343, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3084,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n1991, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1344, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3090,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n1997, B => boothmul_pipelined_i_sum_B_in_4_24_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1345, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3089
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n1996, B => boothmul_pipelined_i_sum_B_in_5_26_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1346, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3088
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n1995, B => boothmul_pipelined_i_sum_B_in_6_28_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1347, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3087
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1348, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n9190, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n1992, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n1992, Q => 
                           DATA2_I_28_port);
   U3 : CLKBUF_X1 port map( A => n7173, Z => n7170);
   U4 : CLKBUF_X1 port map( A => n7173, Z => n7171);
   U5 : CLKBUF_X1 port map( A => n7173, Z => n7172);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n7173);
   U7 : CLKBUF_X1 port map( A => n7177, Z => n7174);
   U8 : CLKBUF_X1 port map( A => n7170, Z => n7175);
   U9 : CLKBUF_X1 port map( A => n7171, Z => n7176);
   U10 : CLKBUF_X1 port map( A => n7171, Z => n7177);
   U11 : CLKBUF_X1 port map( A => n7171, Z => n7178);
   U12 : CLKBUF_X1 port map( A => n7171, Z => n7179);
   U13 : CLKBUF_X1 port map( A => n7172, Z => n7180);
   U14 : CLKBUF_X1 port map( A => n7172, Z => n7181);
   U15 : CLKBUF_X1 port map( A => n7172, Z => n7182);
   U16 : CLKBUF_X1 port map( A => n7172, Z => n7183);
   U17 : CLKBUF_X1 port map( A => n7172, Z => n7184);
   U18 : NOR2_X2 port map( A1 => n7234, A2 => DATA2(2), ZN => n7978);
   U19 : AOI211_X4 port map( C1 => n8890, C2 => n7439, A => n8889, B => n8888, 
                           ZN => n8832);
   U20 : INV_X1 port map( A => n1992, ZN => n8858);
   U21 : CLKBUF_X1 port map( A => n8893, Z => n8883);
   U22 : CLKBUF_X1 port map( A => DATA1(14), Z => n9195);
   U23 : CLKBUF_X1 port map( A => DATA1(6), Z => n9192);
   U24 : CLKBUF_X1 port map( A => DATA1(3), Z => n9191);
   U25 : CLKBUF_X1 port map( A => DATA1(7), Z => n9193);
   U26 : NOR2_X1 port map( A1 => FUNC(2), A2 => FUNC(0), ZN => n7219);
   U27 : INV_X1 port map( A => FUNC(1), ZN => n8709);
   U28 : NAND2_X1 port map( A1 => n7219, A2 => n8709, ZN => n1992);
   U29 : CLKBUF_X1 port map( A => n1992, Z => n9190);
   U30 : CLKBUF_X1 port map( A => DATA1(13), Z => n9194);
   U31 : INV_X1 port map( A => data1_mul_0_port, ZN => n1983);
   U32 : INV_X1 port map( A => data2_mul_1_port, ZN => n7185);
   U33 : NOR2_X1 port map( A1 => boothmul_pipelined_i_encoder_out_0_0_port, A2 
                           => n7185, ZN => n7196);
   U34 : CLKBUF_X1 port map( A => n7196, Z => n9165);
   U35 : NAND2_X1 port map( A1 => n7185, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n9168);
   U36 : INV_X1 port map( A => n9168, ZN => n7202);
   U37 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n8895);
   U38 : NOR2_X1 port map( A1 => n7185, A2 => n8895, ZN => n9166);
   U39 : CLKBUF_X1 port map( A => n9166, Z => n7199);
   U40 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, A2
                           => n9165, B1 => data1_mul_14_port, B2 => n7202, C1 
                           => boothmul_pipelined_i_muxes_in_0_103_port, C2 => 
                           n7199, ZN => n7186);
   U41 : INV_X1 port map( A => n7186, ZN => n1956);
   U42 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, A2
                           => n9165, B1 => data1_mul_13_port, B2 => n7202, C1 
                           => boothmul_pipelined_i_muxes_in_0_104_port, C2 => 
                           n9166, ZN => n7187);
   U43 : INV_X1 port map( A => n7187, ZN => n1958);
   U44 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, A2
                           => n9165, B1 => data1_mul_12_port, B2 => n7202, C1 
                           => boothmul_pipelined_i_muxes_in_0_105_port, C2 => 
                           n7199, ZN => n7188);
   U45 : INV_X1 port map( A => n7188, ZN => n1960);
   U46 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, A2
                           => n9165, B1 => data1_mul_11_port, B2 => n7202, C1 
                           => boothmul_pipelined_i_muxes_in_0_106_port, C2 => 
                           n9166, ZN => n7189);
   U47 : INV_X1 port map( A => n7189, ZN => n1962);
   U48 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, A2
                           => n7196, B1 => data1_mul_10_port, B2 => n7202, C1 
                           => boothmul_pipelined_i_muxes_in_0_107_port, C2 => 
                           n7199, ZN => n7190);
   U49 : INV_X1 port map( A => n7190, ZN => n1964);
   U50 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, A2
                           => n7196, B1 => data1_mul_9_port, B2 => n7202, C1 =>
                           boothmul_pipelined_i_muxes_in_0_108_port, C2 => 
                           n7199, ZN => n7191);
   U51 : INV_X1 port map( A => n7191, ZN => n1966);
   U52 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, A2
                           => n7196, B1 => data1_mul_8_port, B2 => n7202, C1 =>
                           boothmul_pipelined_i_muxes_in_0_109_port, C2 => 
                           n7199, ZN => n7192);
   U53 : INV_X1 port map( A => n7192, ZN => n1968);
   U54 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, A2
                           => n7196, B1 => data1_mul_7_port, B2 => n7202, C1 =>
                           boothmul_pipelined_i_muxes_in_0_110_port, C2 => 
                           n9166, ZN => n7193);
   U55 : INV_X1 port map( A => n7193, ZN => n1970);
   U56 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, A2
                           => n7196, B1 => data1_mul_6_port, B2 => n7202, C1 =>
                           boothmul_pipelined_i_muxes_in_0_111_port, C2 => 
                           n7199, ZN => n7194);
   U57 : INV_X1 port map( A => n7194, ZN => n1972);
   U58 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, A2
                           => n7196, B1 => data1_mul_5_port, B2 => n7202, C1 =>
                           boothmul_pipelined_i_muxes_in_0_112_port, C2 => 
                           n7199, ZN => n7195);
   U59 : INV_X1 port map( A => n7195, ZN => n1974);
   U60 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, A2
                           => n7196, B1 => data1_mul_4_port, B2 => n7202, C1 =>
                           boothmul_pipelined_i_muxes_in_0_113_port, C2 => 
                           n9166, ZN => n7197);
   U61 : INV_X1 port map( A => n7197, ZN => n1976);
   U62 : AOI222_X1 port map( A1 => n9165, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           data1_mul_3_port, B2 => n7202, C1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, C2 => 
                           n9166, ZN => n7198);
   U63 : INV_X1 port map( A => n7198, ZN => n1978);
   U64 : AOI222_X1 port map( A1 => data1_mul_0_port, A2 => n9165, B1 => 
                           data1_mul_1_port, B2 => n7202, C1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C2 => 
                           n7199, ZN => n7200);
   U65 : INV_X1 port map( A => n7200, ZN => n1981);
   U66 : INV_X1 port map( A => FUNC(2), ZN => n7220);
   U67 : NOR3_X1 port map( A1 => FUNC(1), A2 => FUNC(0), A3 => n7220, ZN => 
                           n7395);
   U68 : INV_X1 port map( A => FUNC(3), ZN => n8857);
   U69 : NAND2_X1 port map( A1 => n7395, A2 => n8857, ZN => n553);
   U70 : INV_X1 port map( A => data1_mul_15_port, ZN => n1955);
   U71 : INV_X1 port map( A => data1_mul_14_port, ZN => n1957);
   U72 : INV_X1 port map( A => data1_mul_13_port, ZN => n1959);
   U73 : INV_X1 port map( A => data1_mul_12_port, ZN => n1961);
   U74 : INV_X1 port map( A => data1_mul_11_port, ZN => n1963);
   U75 : INV_X1 port map( A => data1_mul_10_port, ZN => n1965);
   U76 : INV_X1 port map( A => data1_mul_9_port, ZN => n1967);
   U77 : INV_X1 port map( A => data1_mul_8_port, ZN => n1969);
   U78 : INV_X1 port map( A => data1_mul_7_port, ZN => n1971);
   U79 : INV_X1 port map( A => data1_mul_6_port, ZN => n1973);
   U80 : INV_X1 port map( A => data1_mul_5_port, ZN => n1975);
   U81 : INV_X1 port map( A => data1_mul_4_port, ZN => n1977);
   U82 : INV_X1 port map( A => data1_mul_3_port, ZN => n1979);
   U83 : INV_X1 port map( A => data1_mul_2_port, ZN => n1980);
   U84 : INV_X1 port map( A => data1_mul_1_port, ZN => n1982);
   U85 : XOR2_X1 port map( A => n1955, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => boothmul_pipelined_i_muxes_in_0_119_port);
   U86 : AOI22_X1 port map( A1 => n9166, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n9165, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n7201);
   U87 : OAI21_X1 port map( B1 => n9168, B2 => n1955, A => n7201, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U88 : AOI222_X1 port map( A1 => n7202, A2 => data1_mul_2_port, B1 => n9166, 
                           B2 => boothmul_pipelined_i_muxes_in_0_115_port, C1 
                           => n9165, C2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n7204);
   U89 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n8936);
   U90 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n8936, ZN => n8896);
   U91 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n8896, ZN => n7203);
   U92 : NOR2_X1 port map( A1 => n7204, A2 => n7203, ZN => n3083);
   U93 : AOI21_X1 port map( B1 => n7204, B2 => n7203, A => n3083, ZN => n3086);
   U94 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n7205);
   U95 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n7205, ZN => n8938);
   U96 : NOR3_X1 port map( A1 => n5130, A2 => n8938, A3 => n1983, ZN => n3085);
   U97 : OR2_X1 port map( A1 => n1983, A2 => n8938, ZN => n7206);
   U98 : AOI21_X1 port map( B1 => n5130, B2 => n7206, A => n3085, ZN => n3091);
   U99 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n7207);
   U100 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, A
                           => n7207, ZN => n8979);
   U101 : NOR3_X1 port map( A1 => n3077, A2 => n5124, A3 => n8979, ZN => n3084)
                           ;
   U102 : AOI221_X1 port map( B1 => n3077, B2 => n5124, C1 => n8979, C2 => 
                           n5124, A => n3084, ZN => n3092);
   U103 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n7208);
   U104 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, A
                           => n7208, ZN => n9015);
   U105 : NOR3_X1 port map( A1 => n5121, A2 => n5131, A3 => n9015, ZN => n3090)
                           ;
   U106 : AOI221_X1 port map( B1 => n5121, B2 => n5131, C1 => n9015, C2 => 
                           n5131, A => n3090, ZN => n3093);
   U107 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n7209);
   U108 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           A => n7209, ZN => n9051);
   U109 : NOR3_X1 port map( A1 => n5122, A2 => n5132, A3 => n9051, ZN => n3089)
                           ;
   U110 : AOI221_X1 port map( B1 => n5122, B2 => n5132, C1 => n9051, C2 => 
                           n5132, A => n3089, ZN => n3094);
   U111 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n7210);
   U112 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           A => n7210, ZN => n9087);
   U113 : NOR3_X1 port map( A1 => n5123, A2 => n5133, A3 => n9087, ZN => n3088)
                           ;
   U114 : AOI221_X1 port map( B1 => n5123, B2 => n5133, C1 => n9087, C2 => 
                           n5133, A => n3088, ZN => n3095);
   U115 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(8), A3 => DATA2(6), A4 
                           => DATA2(7), ZN => n7218);
   U116 : NOR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n7439);
   U117 : INV_X1 port map( A => DATA2(3), ZN => n8889);
   U118 : OR2_X1 port map( A1 => DATA2(4), A2 => DATA2(5), ZN => n8051);
   U119 : INV_X1 port map( A => n8051, ZN => n8101);
   U120 : NAND2_X1 port map( A1 => n8889, A2 => n8101, ZN => n7234);
   U121 : NAND2_X1 port map( A1 => n7439, A2 => n7978, ZN => n7893);
   U122 : INV_X1 port map( A => DATA2(12), ZN => n8878);
   U123 : INV_X1 port map( A => DATA2(10), ZN => n8880);
   U124 : INV_X1 port map( A => DATA2(11), ZN => n8879);
   U125 : INV_X1 port map( A => DATA2(13), ZN => n8877);
   U126 : NAND4_X1 port map( A1 => n8878, A2 => n8880, A3 => n8879, A4 => n8877
                           , ZN => n7211);
   U127 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n7893, A4 
                           => n7211, ZN => n7217);
   U128 : NOR4_X1 port map( A1 => DATA1(15), A2 => n9195, A3 => n9194, A4 => 
                           DATA1(12), ZN => n7215);
   U129 : NOR4_X1 port map( A1 => DATA1(11), A2 => DATA1(10), A3 => DATA1(9), 
                           A4 => DATA1(8), ZN => n7214);
   U130 : NOR4_X1 port map( A1 => DATA1(7), A2 => DATA1(6), A3 => DATA1(5), A4 
                           => DATA1(4), ZN => n7213);
   U131 : NOR4_X1 port map( A1 => n9191, A2 => DATA1(2), A3 => DATA1(1), A4 => 
                           DATA1(0), ZN => n7212);
   U132 : AND4_X1 port map( A1 => n7215, A2 => n7214, A3 => n7213, A4 => n7212,
                           ZN => n7216);
   U133 : AOI211_X1 port map( C1 => n7218, C2 => n7217, A => n7216, B => n553, 
                           ZN => n8514);
   U134 : CLKBUF_X1 port map( A => n8514, Z => n8575);
   U135 : NAND2_X1 port map( A1 => FUNC(1), A2 => n7219, ZN => n8525);
   U136 : INV_X1 port map( A => n8525, ZN => n8567);
   U137 : INV_X1 port map( A => DATA1(9), ZN => n7679);
   U138 : NOR2_X1 port map( A1 => n7679, A2 => DATA2(9), ZN => n8656);
   U139 : INV_X1 port map( A => n8656, ZN => n8598);
   U140 : NAND2_X1 port map( A1 => DATA2(9), A2 => n7679, ZN => n8657);
   U141 : NAND2_X1 port map( A1 => n8598, A2 => n8657, ZN => n8725);
   U142 : AOI22_X1 port map( A1 => dataout_mul_9_port, A2 => n8575, B1 => n8567
                           , B2 => n8725, ZN => n7399);
   U143 : INV_X1 port map( A => DATA2(2), ZN => n8890);
   U144 : INV_X1 port map( A => DATA2(4), ZN => n8888);
   U145 : NOR2_X1 port map( A1 => n8890, A2 => n8888, ZN => n7420);
   U146 : NAND2_X1 port map( A1 => DATA2(3), A2 => n7420, ZN => n8021);
   U147 : INV_X1 port map( A => DATA2(1), ZN => n8891);
   U148 : NOR2_X1 port map( A1 => n8021, A2 => n8891, ZN => n8842);
   U149 : OR4_X1 port map( A1 => DATA2(5), A2 => FUNC(0), A3 => n8709, A4 => 
                           n7220, ZN => n8036);
   U150 : AOI21_X1 port map( B1 => DATA2(0), B2 => n8842, A => n8036, ZN => 
                           n7393);
   U151 : NAND2_X1 port map( A1 => FUNC(3), A2 => n7393, ZN => n8536);
   U152 : INV_X1 port map( A => n8536, ZN => n8848);
   U153 : INV_X1 port map( A => n7420, ZN => n7282);
   U154 : NAND2_X1 port map( A1 => DATA2(0), A2 => n8891, ZN => n8020);
   U155 : NOR3_X1 port map( A1 => DATA2(3), A2 => n7282, A3 => n8020, ZN => 
                           n8351);
   U156 : INV_X1 port map( A => n8351, ZN => n8821);
   U157 : NAND2_X1 port map( A1 => n7439, A2 => n8890, ZN => n7221);
   U158 : OAI21_X1 port map( B1 => DATA2(3), B2 => n7221, A => n8051, ZN => 
                           n8805);
   U159 : CLKBUF_X1 port map( A => n8805, Z => n8485);
   U160 : NAND2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n7315);
   U161 : INV_X1 port map( A => n7315, ZN => n7419);
   U162 : NAND2_X1 port map( A1 => DATA2(3), A2 => n7419, ZN => n7525);
   U163 : OAI21_X1 port map( B1 => n8890, B2 => n7525, A => n8101, ZN => n7862)
                           ;
   U164 : INV_X1 port map( A => n7862, ZN => n8456);
   U165 : NOR2_X1 port map( A1 => n8051, A2 => n8456, ZN => n8431);
   U166 : CLKBUF_X1 port map( A => n8431, Z => n7943);
   U167 : INV_X1 port map( A => n7943, ZN => n8803);
   U168 : INV_X1 port map( A => n7439, ZN => n7606);
   U169 : OR4_X1 port map( A1 => n8889, A2 => n8890, A3 => n8051, A4 => n7606, 
                           ZN => n8788);
   U170 : INV_X1 port map( A => n8788, ZN => n8496);
   U171 : CLKBUF_X1 port map( A => DATA1(19), Z => n8365);
   U172 : INV_X1 port map( A => n7893, ZN => n8323);
   U173 : INV_X1 port map( A => n7978, ZN => n8087);
   U174 : CLKBUF_X1 port map( A => n8087, Z => n7776);
   U175 : AOI22_X1 port map( A1 => n8365, A2 => n8323, B1 => DATA1(23), B2 => 
                           n7776, ZN => n7222);
   U176 : INV_X1 port map( A => DATA2(0), ZN => n8892);
   U177 : NAND3_X1 port map( A1 => n8892, A2 => DATA2(1), A3 => n7978, ZN => 
                           n8130);
   U178 : INV_X1 port map( A => n8130, ZN => n8152);
   U179 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(21), ZN => n7748);
   U180 : NOR2_X1 port map( A1 => n8087, A2 => n8020, ZN => n7896);
   U181 : INV_X1 port map( A => n7896, ZN => n8312);
   U182 : INV_X1 port map( A => n8312, ZN => n8153);
   U183 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(20), ZN => n7666);
   U184 : NAND2_X1 port map( A1 => n7978, A2 => n7419, ZN => n7680);
   U185 : INV_X1 port map( A => n7680, ZN => n7832);
   U186 : NAND2_X1 port map( A1 => n7832, A2 => DATA1(22), ZN => n7779);
   U187 : NAND4_X1 port map( A1 => n7222, A2 => n7748, A3 => n7666, A4 => n7779
                           , ZN => n7256);
   U188 : OAI21_X1 port map( B1 => n7234, B2 => DATA2(1), A => n8087, ZN => 
                           n7982);
   U189 : INV_X1 port map( A => n7982, ZN => n8772);
   U190 : CLKBUF_X1 port map( A => DATA1(17), Z => n8403);
   U191 : CLKBUF_X1 port map( A => n8323, Z => n8762);
   U192 : AOI22_X1 port map( A1 => n8403, A2 => n8762, B1 => DATA1(21), B2 => 
                           n7776, ZN => n7223);
   U193 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(19), ZN => n7667);
   U194 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(18), ZN => n7641);
   U195 : CLKBUF_X1 port map( A => n7832, Z => n8763);
   U196 : NAND2_X1 port map( A1 => n8763, A2 => DATA1(20), ZN => n7749);
   U197 : NAND4_X1 port map( A1 => n7223, A2 => n7667, A3 => n7641, A4 => n7749
                           , ZN => n7235);
   U198 : OAI21_X1 port map( B1 => n8892, B2 => n8890, A => n7982, ZN => n7224)
                           ;
   U199 : INV_X1 port map( A => n7224, ZN => n8770);
   U200 : INV_X1 port map( A => DATA1(20), ZN => n8681);
   U201 : NOR2_X1 port map( A1 => n8130, A2 => n8681, ZN => n7711);
   U202 : INV_X1 port map( A => DATA1(22), ZN => n8618);
   U203 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(18), ZN => n7646);
   U204 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(19), ZN => n7661);
   U205 : OAI211_X1 port map( C1 => n7978, C2 => n8618, A => n7646, B => n7661,
                           ZN => n7225);
   U206 : AOI211_X1 port map( C1 => DATA1(21), C2 => n8763, A => n7711, B => 
                           n7225, ZN => n7226);
   U207 : INV_X1 port map( A => n7226, ZN => n7254);
   U208 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(0), ZN => n7263);
   U209 : NOR3_X1 port map( A1 => DATA2(1), A2 => n7263, A3 => n7234, ZN => 
                           n7506);
   U210 : CLKBUF_X1 port map( A => n7506, Z => n8768);
   U211 : AOI222_X1 port map( A1 => n7256, A2 => n8772, B1 => n7235, B2 => 
                           n8770, C1 => n7254, C2 => n8768, ZN => n7276);
   U212 : NAND2_X1 port map( A1 => n8101, A2 => n8890, ZN => n7250);
   U213 : OAI21_X1 port map( B1 => DATA2(1), B2 => n7250, A => n7234, ZN => 
                           n7227);
   U214 : INV_X1 port map( A => n7227, ZN => n8785);
   U215 : INV_X1 port map( A => n8785, ZN => n8331);
   U216 : NOR3_X1 port map( A1 => n8889, A2 => n7606, A3 => n7250, ZN => n8272)
                           ;
   U217 : CLKBUF_X1 port map( A => n8272, Z => n8229);
   U218 : INV_X1 port map( A => n7982, ZN => n7586);
   U219 : AOI22_X1 port map( A1 => n8762, A2 => DATA1(15), B1 => n8365, B2 => 
                           n7776, ZN => n7228);
   U220 : NAND2_X1 port map( A1 => n8152, A2 => n8403, ZN => n7642);
   U221 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(16), ZN => n7638);
   U222 : NAND2_X1 port map( A1 => n8763, A2 => DATA1(18), ZN => n7668);
   U223 : NAND4_X1 port map( A1 => n7228, A2 => n7642, A3 => n7638, A4 => n7668
                           , ZN => n7233);
   U224 : AOI22_X1 port map( A1 => n8323, A2 => DATA1(16), B1 => DATA1(20), B2 
                           => n7776, ZN => n7229);
   U225 : NAND2_X1 port map( A1 => n8763, A2 => n8365, ZN => n7713);
   U226 : NAND2_X1 port map( A1 => n7896, A2 => DATA1(17), ZN => n7647);
   U227 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(18), ZN => n7662);
   U228 : NAND4_X1 port map( A1 => n7229, A2 => n7713, A3 => n7647, A4 => n7662
                           , ZN => n7236);
   U229 : AOI222_X1 port map( A1 => n7235, A2 => n7586, B1 => n7233, B2 => 
                           n8770, C1 => n7236, C2 => n7506, ZN => n7252);
   U230 : INV_X1 port map( A => n7252, ZN => n7262);
   U231 : AOI22_X1 port map( A1 => DATA1(13), A2 => n8762, B1 => DATA1(17), B2 
                           => n7776, ZN => n7230);
   U232 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(15), ZN => n7639);
   U233 : NAND2_X1 port map( A1 => n9195, A2 => n7896, ZN => n7656);
   U234 : NAND2_X1 port map( A1 => DATA1(16), A2 => n8763, ZN => n7644);
   U235 : NAND4_X1 port map( A1 => n7230, A2 => n7639, A3 => n7656, A4 => n7644
                           , ZN => n7242);
   U236 : INV_X1 port map( A => DATA1(15), ZN => n8434);
   U237 : NOR2_X1 port map( A1 => n8434, A2 => n8312, ZN => n7655);
   U238 : INV_X1 port map( A => n9195, ZN => n8454);
   U239 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(16), ZN => n7648);
   U240 : NAND2_X1 port map( A1 => DATA1(18), A2 => n8087, ZN => n7714);
   U241 : OAI211_X1 port map( C1 => n7893, C2 => n8454, A => n7648, B => n7714,
                           ZN => n7231);
   U242 : AOI211_X1 port map( C1 => DATA1(17), C2 => n7832, A => n7655, B => 
                           n7231, ZN => n7232);
   U243 : INV_X1 port map( A => n7232, ZN => n7241);
   U244 : AOI222_X1 port map( A1 => n7233, A2 => n7586, B1 => n7242, B2 => 
                           n8770, C1 => n7241, C2 => n7506, ZN => n7353);
   U245 : INV_X1 port map( A => n7353, ZN => n7243);
   U246 : OAI21_X1 port map( B1 => DATA2(0), B2 => n7234, A => n7586, ZN => 
                           n8231);
   U247 : INV_X1 port map( A => n8231, ZN => n8777);
   U248 : INV_X1 port map( A => n8777, ZN => n8203);
   U249 : AOI22_X1 port map( A1 => n8229, A2 => n7262, B1 => n7243, B2 => n8203
                           , ZN => n7238);
   U250 : NOR2_X1 port map( A1 => n7234, A2 => n8203, ZN => n7919);
   U251 : AOI222_X1 port map( A1 => n7236, A2 => n7586, B1 => n7241, B2 => 
                           n8770, C1 => n7233, C2 => n8768, ZN => n7269);
   U252 : INV_X1 port map( A => n7269, ZN => n7247);
   U253 : NAND3_X1 port map( A1 => n7606, A2 => n7234, A3 => n8331, ZN => n8780
                           );
   U254 : INV_X1 port map( A => n8780, ZN => n8335);
   U255 : AOI222_X1 port map( A1 => n8770, A2 => n7236, B1 => n8768, B2 => 
                           n7235, C1 => n7586, C2 => n7254, ZN => n7259);
   U256 : INV_X1 port map( A => n7259, ZN => n7279);
   U257 : AOI22_X1 port map( A1 => n7919, A2 => n7247, B1 => n8335, B2 => n7279
                           , ZN => n7237);
   U258 : OAI211_X1 port map( C1 => n7276, C2 => n8331, A => n7238, B => n7237,
                           ZN => n7357);
   U259 : CLKBUF_X1 port map( A => DATA1(12), Z => n8504);
   U260 : AOI22_X1 port map( A1 => n8504, A2 => n8323, B1 => DATA1(16), B2 => 
                           n8087, ZN => n7239);
   U261 : NAND2_X1 port map( A1 => n8152, A2 => n9195, ZN => n7653);
   U262 : NAND2_X1 port map( A1 => n8153, A2 => n9194, ZN => n7691);
   U263 : NAND2_X1 port map( A1 => DATA1(15), A2 => n7832, ZN => n7649);
   U264 : NAND4_X1 port map( A1 => n7239, A2 => n7653, A3 => n7691, A4 => n7649
                           , ZN => n7268);
   U265 : AOI22_X1 port map( A1 => DATA1(14), A2 => n7832, B1 => n8762, B2 => 
                           DATA1(11), ZN => n7240);
   U266 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(13), ZN => n7657);
   U267 : NAND2_X1 port map( A1 => n7896, A2 => n8504, ZN => n7677);
   U268 : NAND2_X1 port map( A1 => DATA1(15), A2 => n8087, ZN => n7643);
   U269 : NAND4_X1 port map( A1 => n7240, A2 => n7657, A3 => n7677, A4 => n7643
                           , ZN => n7352);
   U270 : AOI222_X1 port map( A1 => n7242, A2 => n7586, B1 => n7268, B2 => 
                           n7506, C1 => n7352, C2 => n8770, ZN => n7445);
   U271 : INV_X1 port map( A => n7445, ZN => n7408);
   U272 : AOI22_X1 port map( A1 => n8335, A2 => n7247, B1 => n7408, B2 => n8203
                           , ZN => n7245);
   U273 : CLKBUF_X1 port map( A => n7919, Z => n8230);
   U274 : AOI222_X1 port map( A1 => n7506, A2 => n7242, B1 => n8770, B2 => 
                           n7268, C1 => n7586, C2 => n7241, ZN => n7405);
   U275 : INV_X1 port map( A => n7405, ZN => n7246);
   U276 : AOI22_X1 port map( A1 => n8229, A2 => n7243, B1 => n8230, B2 => n7246
                           , ZN => n7244);
   U277 : OAI211_X1 port map( C1 => n7252, C2 => n8331, A => n7245, B => n7244,
                           ZN => n7448);
   U278 : INV_X1 port map( A => n7448, ZN => n7413);
   U279 : INV_X1 port map( A => n8051, ZN => n8798);
   U280 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(2), ZN => n7251);
   U281 : NAND3_X1 port map( A1 => n8798, A2 => n7251, A3 => n7525, ZN => n8786
                           );
   U282 : INV_X1 port map( A => n7919, ZN => n8044);
   U283 : AOI22_X1 port map( A1 => n8229, A2 => n7247, B1 => n8231, B2 => n7246
                           , ZN => n7249);
   U284 : AOI22_X1 port map( A1 => n8785, A2 => n7279, B1 => n8335, B2 => n7262
                           , ZN => n7248);
   U285 : OAI211_X1 port map( C1 => n7353, C2 => n8044, A => n7249, B => n7248,
                           ZN => n7409);
   U286 : INV_X1 port map( A => n7409, ZN => n7360);
   U287 : OR2_X1 port map( A1 => n7250, A2 => n7525, ZN => n8790);
   U288 : OAI22_X1 port map( A1 => n7413, A2 => n8786, B1 => n7360, B2 => n8790
                           , ZN => n7265);
   U289 : OAI21_X1 port map( B1 => n8891, B2 => n7251, A => n8101, ZN => n8339)
                           ;
   U290 : INV_X1 port map( A => n8339, ZN => n8793);
   U291 : INV_X1 port map( A => n7276, ZN => n7287);
   U292 : OAI22_X1 port map( A1 => n8777, A2 => n7252, B1 => n7259, B2 => n8044
                           , ZN => n7258);
   U293 : AOI22_X1 port map( A1 => n8763, A2 => DATA1(23), B1 => n8762, B2 => 
                           DATA1(20), ZN => n7253);
   U294 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(22), ZN => n7765);
   U295 : CLKBUF_X1 port map( A => DATA1(21), Z => n8286);
   U296 : NAND2_X1 port map( A1 => n8153, A2 => n8286, ZN => n7712);
   U297 : CLKBUF_X1 port map( A => DATA1(24), Z => n8692);
   U298 : NAND2_X1 port map( A1 => n8692, A2 => n8087, ZN => n7850);
   U299 : NAND4_X1 port map( A1 => n7253, A2 => n7765, A3 => n7712, A4 => n7850
                           , ZN => n7275);
   U300 : AOI222_X1 port map( A1 => n7275, A2 => n8772, B1 => n7254, B2 => 
                           n8770, C1 => n7256, C2 => n8768, ZN => n7291);
   U301 : AOI22_X1 port map( A1 => n7832, A2 => DATA1(24), B1 => n8762, B2 => 
                           DATA1(21), ZN => n7255);
   U302 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(23), ZN => n7778);
   U303 : NAND2_X1 port map( A1 => n7896, A2 => DATA1(22), ZN => n7747);
   U304 : NAND2_X1 port map( A1 => DATA1(25), A2 => n8087, ZN => n7874);
   U305 : NAND4_X1 port map( A1 => n7255, A2 => n7778, A3 => n7747, A4 => n7874
                           , ZN => n7284);
   U306 : AOI222_X1 port map( A1 => n7284, A2 => n8772, B1 => n7256, B2 => 
                           n8770, C1 => n7275, C2 => n7506, ZN => n7293);
   U307 : OAI22_X1 port map( A1 => n7291, A2 => n8780, B1 => n7293, B2 => n8331
                           , ZN => n7257);
   U308 : AOI211_X1 port map( C1 => n8229, C2 => n7287, A => n7258, B => n7257,
                           ZN => n7304);
   U309 : OAI22_X1 port map( A1 => n8777, A2 => n7269, B1 => n7291, B2 => n8331
                           , ZN => n7261);
   U310 : INV_X1 port map( A => n8272, ZN => n8774);
   U311 : CLKBUF_X1 port map( A => n8774, Z => n8330);
   U312 : OAI22_X1 port map( A1 => n7259, A2 => n8330, B1 => n7276, B2 => n8780
                           , ZN => n7260);
   U313 : AOI211_X1 port map( C1 => n7919, C2 => n7262, A => n7261, B => n7260,
                           ZN => n7299);
   U314 : CLKBUF_X1 port map( A => n8339, Z => n7995);
   U315 : NOR3_X1 port map( A1 => n8889, A2 => n7263, A3 => n7995, ZN => n8797)
                           ;
   U316 : INV_X1 port map( A => n8797, ZN => n8477);
   U317 : OAI22_X1 port map( A1 => n8793, A2 => n7304, B1 => n7299, B2 => n8477
                           , ZN => n7264);
   U318 : AOI211_X1 port map( C1 => n8496, C2 => n7357, A => n7265, B => n7264,
                           ZN => n7361);
   U319 : CLKBUF_X1 port map( A => n7862, Z => n8801);
   U320 : INV_X1 port map( A => n8786, ZN => n8522);
   U321 : INV_X1 port map( A => DATA1(11), ZN => n8526);
   U322 : NOR2_X1 port map( A1 => n8312, A2 => n8526, ZN => n7684);
   U323 : NAND2_X1 port map( A1 => n8762, A2 => DATA1(10), ZN => n7727);
   U324 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(12), ZN => n7690);
   U325 : OAI211_X1 port map( C1 => n7978, C2 => n8454, A => n7727, B => n7690,
                           ZN => n7266);
   U326 : AOI211_X1 port map( C1 => n9194, C2 => n8763, A => n7684, B => n7266,
                           ZN => n7267);
   U327 : INV_X1 port map( A => n7267, ZN => n7404);
   U328 : AOI222_X1 port map( A1 => n8770, A2 => n7404, B1 => n8768, B2 => 
                           n7352, C1 => n7586, C2 => n7268, ZN => n7473);
   U329 : OAI22_X1 port map( A1 => n7473, A2 => n8777, B1 => n7353, B2 => n8780
                           , ZN => n7271);
   U330 : OAI22_X1 port map( A1 => n7405, A2 => n8774, B1 => n7269, B2 => n8331
                           , ZN => n7270);
   U331 : AOI211_X1 port map( C1 => n7919, C2 => n7408, A => n7271, B => n7270,
                           ZN => n7477);
   U332 : INV_X1 port map( A => n7477, ZN => n7410);
   U333 : INV_X1 port map( A => n7357, ZN => n7300);
   U334 : OAI22_X1 port map( A1 => n8793, A2 => n7299, B1 => n7300, B2 => n8477
                           , ZN => n7272);
   U335 : AOI21_X1 port map( B1 => n8522, B2 => n7410, A => n7272, ZN => n7273)
                           ;
   U336 : OAI21_X1 port map( B1 => n7413, B2 => n8790, A => n7273, ZN => n7414)
                           ;
   U337 : AOI21_X1 port map( B1 => n8496, B2 => n7409, A => n7414, ZN => n7363)
                           ;
   U338 : INV_X1 port map( A => n7299, ZN => n7298);
   U339 : OAI22_X1 port map( A1 => n7360, A2 => n8786, B1 => n7300, B2 => n8790
                           , ZN => n7281);
   U340 : OAI22_X1 port map( A1 => n7291, A2 => n8330, B1 => n7293, B2 => n8780
                           , ZN => n7278);
   U341 : AOI22_X1 port map( A1 => n8763, A2 => DATA1(25), B1 => n8762, B2 => 
                           DATA1(22), ZN => n7274);
   U342 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(24), ZN => n7815);
   U343 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(23), ZN => n7764);
   U344 : NAND2_X1 port map( A1 => DATA1(26), A2 => n8087, ZN => n7891);
   U345 : NAND4_X1 port map( A1 => n7274, A2 => n7815, A3 => n7764, A4 => n7891
                           , ZN => n7290);
   U346 : AOI222_X1 port map( A1 => n7290, A2 => n8772, B1 => n7275, B2 => 
                           n8770, C1 => n7284, C2 => n7506, ZN => n7325);
   U347 : OAI22_X1 port map( A1 => n7276, A2 => n8044, B1 => n7325, B2 => n8331
                           , ZN => n7277);
   U348 : AOI211_X1 port map( C1 => n8203, C2 => n7279, A => n7278, B => n7277,
                           ZN => n7332);
   U349 : OAI22_X1 port map( A1 => n8793, A2 => n7332, B1 => n7304, B2 => n8477
                           , ZN => n7280);
   U350 : AOI211_X1 port map( C1 => n8496, C2 => n7298, A => n7281, B => n7280,
                           ZN => n7318);
   U351 : OAI222_X1 port map( A1 => n8803, A2 => n7361, B1 => n8801, B2 => 
                           n7363, C1 => n7318, C2 => n8101, ZN => n7483);
   U352 : NOR2_X1 port map( A1 => n8889, A2 => n8101, ZN => n8111);
   U353 : INV_X1 port map( A => n8111, ZN => n8819);
   U354 : NAND2_X1 port map( A1 => n7282, A2 => n8819, ZN => n8809);
   U355 : NOR4_X1 port map( A1 => n8891, A2 => n8809, A3 => n8101, A4 => 
                           DATA2(0), ZN => n8103);
   U356 : CLKBUF_X1 port map( A => n8103, Z => n8807);
   U357 : OAI22_X1 port map( A1 => n7291, A2 => n8044, B1 => n7325, B2 => n8780
                           , ZN => n7286);
   U358 : AOI22_X1 port map( A1 => DATA1(23), A2 => n8762, B1 => DATA1(27), B2 
                           => n7776, ZN => n7283);
   U359 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(25), ZN => n7829);
   U360 : NAND2_X1 port map( A1 => n7896, A2 => n8692, ZN => n7777);
   U361 : NAND2_X1 port map( A1 => n7832, A2 => DATA1(26), ZN => n7873);
   U362 : NAND4_X1 port map( A1 => n7283, A2 => n7829, A3 => n7777, A4 => n7873
                           , ZN => n7307);
   U363 : AOI222_X1 port map( A1 => n7307, A2 => n8772, B1 => n7284, B2 => 
                           n8770, C1 => n7290, C2 => n8768, ZN => n7324);
   U364 : OAI22_X1 port map( A1 => n7293, A2 => n8774, B1 => n7324, B2 => n8331
                           , ZN => n7285);
   U365 : AOI211_X1 port map( C1 => n8203, C2 => n7287, A => n7286, B => n7285,
                           ZN => n7329);
   U366 : NAND2_X1 port map( A1 => n7832, A2 => DATA1(27), ZN => n7892);
   U367 : INV_X1 port map( A => n7892, ZN => n7289);
   U368 : INV_X1 port map( A => DATA1(28), ZN => n8700);
   U369 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(25), ZN => n7814);
   U370 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(26), ZN => n7848);
   U371 : OAI211_X1 port map( C1 => n7978, C2 => n8700, A => n7814, B => n7848,
                           ZN => n7288);
   U372 : AOI211_X1 port map( C1 => n8692, C2 => n8762, A => n7289, B => n7288,
                           ZN => n7323);
   U373 : INV_X1 port map( A => n7323, ZN => n7306);
   U374 : AOI222_X1 port map( A1 => n8770, A2 => n7290, B1 => n8768, B2 => 
                           n7307, C1 => n7586, C2 => n7306, ZN => n8270);
   U375 : OAI22_X1 port map( A1 => n8331, A2 => n8270, B1 => n8777, B2 => n7291
                           , ZN => n7292);
   U376 : INV_X1 port map( A => n7292, ZN => n7295);
   U377 : INV_X1 port map( A => n7293, ZN => n7310);
   U378 : INV_X1 port map( A => n7324, ZN => n7340);
   U379 : AOI22_X1 port map( A1 => n8230, A2 => n7310, B1 => n8335, B2 => n7340
                           , ZN => n7294);
   U380 : OAI211_X1 port map( C1 => n7325, C2 => n8330, A => n7295, B => n7294,
                           ZN => n8384);
   U381 : INV_X1 port map( A => n8384, ZN => n7311);
   U382 : OAI22_X1 port map( A1 => n8477, A2 => n7329, B1 => n8793, B2 => n7311
                           , ZN => n7297);
   U383 : OAI22_X1 port map( A1 => n8788, A2 => n7332, B1 => n8790, B2 => n7304
                           , ZN => n7296);
   U384 : AOI211_X1 port map( C1 => n7298, C2 => n8522, A => n7297, B => n7296,
                           ZN => n7320);
   U385 : OAI22_X1 port map( A1 => n7299, A2 => n8790, B1 => n7332, B2 => n8477
                           , ZN => n7302);
   U386 : OAI22_X1 port map( A1 => n8793, A2 => n7329, B1 => n7300, B2 => n8786
                           , ZN => n7301);
   U387 : NOR2_X1 port map( A1 => n7302, A2 => n7301, ZN => n7317);
   U388 : OAI21_X1 port map( B1 => n7304, B2 => n8788, A => n7317, ZN => n7303)
                           ;
   U389 : INV_X1 port map( A => n7303, ZN => n7314);
   U390 : OAI222_X1 port map( A1 => n7320, A2 => n8101, B1 => n7314, B2 => 
                           n8803, C1 => n7318, C2 => n8801, ZN => n8497);
   U391 : OAI22_X1 port map( A1 => n7304, A2 => n8786, B1 => n7332, B2 => n8790
                           , ZN => n7313);
   U392 : AOI22_X1 port map( A1 => DATA1(25), A2 => n8323, B1 => DATA1(29), B2 
                           => n7776, ZN => n7305);
   U393 : NAND2_X1 port map( A1 => n7896, A2 => DATA1(26), ZN => n7828);
   U394 : NAND2_X1 port map( A1 => n8763, A2 => DATA1(28), ZN => n7977);
   U395 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(27), ZN => n7872);
   U396 : NAND4_X1 port map( A1 => n7305, A2 => n7828, A3 => n7977, A4 => n7872
                           , ZN => n7321);
   U397 : AOI222_X1 port map( A1 => n7321, A2 => n8772, B1 => n7307, B2 => 
                           n8770, C1 => n7306, C2 => n8768, ZN => n8269);
   U398 : OAI22_X1 port map( A1 => n8270, A2 => n8780, B1 => n8269, B2 => n8331
                           , ZN => n7309);
   U399 : OAI22_X1 port map( A1 => n7325, A2 => n8044, B1 => n7324, B2 => n8774
                           , ZN => n7308);
   U400 : AOI211_X1 port map( C1 => n8203, C2 => n7310, A => n7309, B => n7308,
                           ZN => n7328);
   U401 : OAI22_X1 port map( A1 => n8793, A2 => n7328, B1 => n7311, B2 => n8477
                           , ZN => n7312);
   U402 : NOR2_X1 port map( A1 => n7313, A2 => n7312, ZN => n7319);
   U403 : OAI222_X1 port map( A1 => n8803, A2 => n7320, B1 => n7862, B2 => 
                           n7314, C1 => n7319, C2 => n8798, ZN => n8501);
   U404 : INV_X1 port map( A => n8501, ZN => n7335);
   U405 : NOR3_X1 port map( A1 => n8888, A2 => n8809, A3 => n7315, ZN => n7316)
                           ;
   U406 : CLKBUF_X1 port map( A => n7316, Z => n8500);
   U407 : INV_X1 port map( A => n8500, ZN => n8814);
   U408 : INV_X1 port map( A => n8485, ZN => n8463);
   U409 : NAND4_X1 port map( A1 => n8890, A2 => n8891, A3 => n8819, A4 => n8463
                           , ZN => n8461);
   U410 : INV_X1 port map( A => n8461, ZN => n8811);
   U411 : OAI222_X1 port map( A1 => n8803, A2 => n7318, B1 => n7862, B2 => 
                           n7361, C1 => n7317, C2 => n8798, ZN => n7440);
   U412 : OAI21_X1 port map( B1 => n8788, B2 => n7329, A => n7319, ZN => n7347)
                           ;
   U413 : INV_X1 port map( A => n7320, ZN => n7333);
   U414 : INV_X1 port map( A => n8770, ZN => n7986);
   U415 : INV_X1 port map( A => n8768, ZN => n7984);
   U416 : INV_X1 port map( A => n7321, ZN => n7339);
   U417 : INV_X1 port map( A => n8772, ZN => n7898);
   U418 : NOR2_X1 port map( A1 => n8130, A2 => n8700, ZN => n7895);
   U419 : INV_X1 port map( A => DATA1(30), ZN => n8577);
   U420 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(26), ZN => n7813);
   U421 : NAND2_X1 port map( A1 => n7896, A2 => DATA1(27), ZN => n7847);
   U422 : OAI211_X1 port map( C1 => n7978, C2 => n8577, A => n7813, B => n7847,
                           ZN => n7322);
   U423 : AOI211_X1 port map( C1 => DATA1(29), C2 => n7832, A => n7895, B => 
                           n7322, ZN => n8188);
   U424 : OAI222_X1 port map( A1 => n7986, A2 => n7323, B1 => n7984, B2 => 
                           n7339, C1 => n7898, C2 => n8188, ZN => n8273);
   U425 : OAI22_X1 port map( A1 => n8270, A2 => n8774, B1 => n8269, B2 => n8780
                           , ZN => n7327);
   U426 : OAI22_X1 port map( A1 => n8777, A2 => n7325, B1 => n7324, B2 => n8044
                           , ZN => n7326);
   U427 : AOI211_X1 port map( C1 => n8785, C2 => n8273, A => n7327, B => n7326,
                           ZN => n7346);
   U428 : INV_X1 port map( A => n7346, ZN => n8386);
   U429 : INV_X1 port map( A => n7328, ZN => n8385);
   U430 : CLKBUF_X1 port map( A => n8797, Z => n8100);
   U431 : AOI22_X1 port map( A1 => n8339, A2 => n8386, B1 => n8385, B2 => n8100
                           , ZN => n7331);
   U432 : INV_X1 port map( A => n7329, ZN => n7343);
   U433 : INV_X1 port map( A => n8790, ZN => n8524);
   U434 : AOI22_X1 port map( A1 => n7343, A2 => n8524, B1 => n8384, B2 => n8496
                           , ZN => n7330);
   U435 : OAI211_X1 port map( C1 => n8786, C2 => n7332, A => n7331, B => n7330,
                           ZN => n8417);
   U436 : AOI222_X1 port map( A1 => n7943, A2 => n7347, B1 => n8456, B2 => 
                           n7333, C1 => n8417, C2 => n8051, ZN => n8462);
   U437 : INV_X1 port map( A => n8462, ZN => n8498);
   U438 : AOI22_X1 port map( A1 => n8811, A2 => n7440, B1 => n8809, B2 => n8498
                           , ZN => n7334);
   U439 : OAI21_X1 port map( B1 => n7335, B2 => n8814, A => n7334, ZN => n7336)
                           ;
   U440 : AOI21_X1 port map( B1 => n8807, B2 => n8497, A => n7336, ZN => n7486)
                           ;
   U441 : INV_X1 port map( A => n7486, ZN => n7337);
   U442 : AOI21_X1 port map( B1 => n8485, B2 => n7483, A => n7337, ZN => n8552)
                           ;
   U443 : NAND4_X1 port map( A1 => n8819, A2 => n8892, A3 => DATA2(1), A4 => 
                           n7420, ZN => n8817);
   U444 : INV_X1 port map( A => n8809, ZN => n8052);
   U445 : INV_X1 port map( A => n8269, ZN => n8232);
   U446 : INV_X1 port map( A => n8768, ZN => n8186);
   U447 : INV_X1 port map( A => DATA1(29), ZN => n8131);
   U448 : NOR2_X1 port map( A1 => n8130, A2 => n8131, ZN => n7980);
   U449 : INV_X1 port map( A => DATA1(31), ZN => n8128);
   U450 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(27), ZN => n7827);
   U451 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(28), ZN => n7871);
   U452 : OAI211_X1 port map( C1 => n7978, C2 => n8128, A => n7827, B => n7871,
                           ZN => n7338);
   U453 : AOI211_X1 port map( C1 => DATA1(30), C2 => n8763, A => n7980, B => 
                           n7338, ZN => n8187);
   U454 : OAI222_X1 port map( A1 => n7986, A2 => n7339, B1 => n8186, B2 => 
                           n8188, C1 => n7898, C2 => n8187, ZN => n8271);
   U455 : AOI22_X1 port map( A1 => n8229, A2 => n8232, B1 => n8785, B2 => n8271
                           , ZN => n7342);
   U456 : AOI22_X1 port map( A1 => n8335, A2 => n8273, B1 => n8203, B2 => n7340
                           , ZN => n7341);
   U457 : OAI211_X1 port map( C1 => n8270, C2 => n8044, A => n7342, B => n7341,
                           ZN => n8387);
   U458 : AOI22_X1 port map( A1 => n8524, A2 => n8384, B1 => n7995, B2 => n8387
                           , ZN => n7345);
   U459 : AOI22_X1 port map( A1 => n8496, A2 => n8385, B1 => n8522, B2 => n7343
                           , ZN => n7344);
   U460 : OAI211_X1 port map( C1 => n7346, C2 => n8477, A => n7345, B => n7344,
                           ZN => n8416);
   U461 : AOI222_X1 port map( A1 => n8416, A2 => n8051, B1 => n8417, B2 => 
                           n7943, C1 => n7347, C2 => n8456, ZN => n8484);
   U462 : INV_X1 port map( A => n7440, ZN => n7415);
   U463 : OAI22_X1 port map( A1 => n8052, A2 => n8484, B1 => n8463, B2 => n7415
                           , ZN => n7349);
   U464 : INV_X1 port map( A => n8497, ZN => n7366);
   U465 : OAI22_X1 port map( A1 => n7366, A2 => n8461, B1 => n8462, B2 => n8814
                           , ZN => n7348);
   U466 : AOI211_X1 port map( C1 => n8807, C2 => n8501, A => n7349, B => n7348,
                           ZN => n8551);
   U467 : INV_X1 port map( A => n7473, ZN => n7356);
   U468 : INV_X1 port map( A => DATA1(10), ZN => n8599);
   U469 : NOR2_X1 port map( A1 => n8312, A2 => n8599, ZN => n7688);
   U470 : INV_X1 port map( A => DATA1(13), ZN => n8474);
   U471 : NAND2_X1 port map( A1 => n8762, A2 => DATA1(9), ZN => n7379);
   U472 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(11), ZN => n7676);
   U473 : OAI211_X1 port map( C1 => n7978, C2 => n8474, A => n7379, B => n7676,
                           ZN => n7350);
   U474 : AOI211_X1 port map( C1 => n8504, C2 => n7832, A => n7688, B => n7350,
                           ZN => n7351);
   U475 : INV_X1 port map( A => n7351, ZN => n7444);
   U476 : AOI222_X1 port map( A1 => n8770, A2 => n7444, B1 => n8768, B2 => 
                           n7404, C1 => n7586, C2 => n7352, ZN => n7508);
   U477 : OAI22_X1 port map( A1 => n8777, A2 => n7508, B1 => n7405, B2 => n8780
                           , ZN => n7355);
   U478 : OAI22_X1 port map( A1 => n7445, A2 => n8774, B1 => n7353, B2 => n8331
                           , ZN => n7354);
   U479 : AOI211_X1 port map( C1 => n8230, C2 => n7356, A => n7355, B => n7354,
                           ZN => n7511);
   U480 : INV_X1 port map( A => n7511, ZN => n7480);
   U481 : AOI22_X1 port map( A1 => n8524, A2 => n7410, B1 => n8522, B2 => n7480
                           , ZN => n7359);
   U482 : AOI22_X1 port map( A1 => n8496, A2 => n7448, B1 => n7995, B2 => n7357
                           , ZN => n7358);
   U483 : OAI211_X1 port map( C1 => n7360, C2 => n8477, A => n7359, B => n7358,
                           ZN => n7451);
   U484 : INV_X1 port map( A => n7451, ZN => n7362);
   U485 : OAI222_X1 port map( A1 => n8803, A2 => n7363, B1 => n7862, B2 => 
                           n7362, C1 => n7361, C2 => n8798, ZN => n7516);
   U486 : AOI22_X1 port map( A1 => n8807, A2 => n7440, B1 => n8485, B2 => n7516
                           , ZN => n7365);
   U487 : AOI22_X1 port map( A1 => n8811, A2 => n7483, B1 => n8809, B2 => n8501
                           , ZN => n7364);
   U488 : OAI211_X1 port map( C1 => n7366, C2 => n8814, A => n7365, B => n7364,
                           ZN => n7523);
   U489 : INV_X1 port map( A => n7523, ZN => n7487);
   U490 : OAI21_X1 port map( B1 => n7606, B2 => n8111, A => n8809, ZN => n8828)
                           ;
   U491 : INV_X1 port map( A => n8828, ZN => n8553);
   U492 : OAI222_X1 port map( A1 => n8821, A2 => n8552, B1 => n8817, B2 => 
                           n8551, C1 => n7487, C2 => n8553, ZN => n7378);
   U493 : NOR2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n7400);
   U494 : XNOR2_X1 port map( A => DATA2_I_9_port, B => DATA1(9), ZN => n7620);
   U495 : NOR2_X1 port map( A1 => n7400, A2 => n7620, ZN => n8556);
   U496 : NAND2_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, ZN => n7372)
                           ;
   U497 : OAI21_X1 port map( B1 => n9193, B2 => DATA2_I_7_port, A => n7372, ZN 
                           => n7463);
   U498 : NAND2_X1 port map( A1 => n9192, A2 => DATA2_I_6_port, ZN => n7435);
   U499 : NAND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n7369)
                           ;
   U500 : INV_X1 port map( A => n7369, ZN => n7434);
   U501 : XOR2_X1 port map( A => DATA2_I_3_port, B => n9191, Z => n7611);
   U502 : NAND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n7431)
                           ;
   U503 : OAI21_X1 port map( B1 => DATA1(2), B2 => DATA2_I_2_port, A => n7431, 
                           ZN => n8125);
   U504 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n7429)
                           ;
   U505 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n8566)
                           ;
   U506 : INV_X1 port map( A => n8566, ZN => n8316);
   U507 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n8320);
   U508 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n7429, 
                           ZN => n8319);
   U509 : NOR2_X1 port map( A1 => n8320, A2 => n8319, ZN => n8318);
   U510 : OAI21_X1 port map( B1 => n8316, B2 => cin, A => n8318, ZN => n7367);
   U511 : OAI221_X1 port map( B1 => n8125, B2 => n7429, C1 => n8125, C2 => 
                           n7367, A => n7431, ZN => n7368);
   U512 : AND2_X1 port map( A1 => n9191, A2 => DATA2_I_3_port, ZN => n7432);
   U513 : AOI21_X1 port map( B1 => n7611, B2 => n7368, A => n7432, ZN => n7370)
                           ;
   U514 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n7433)
                           ;
   U515 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n7433, 
                           ZN => n7572);
   U516 : OAI21_X1 port map( B1 => DATA1(5), B2 => DATA2_I_5_port, A => n7369, 
                           ZN => n7535);
   U517 : AOI221_X1 port map( B1 => n7370, B2 => n7433, C1 => n7572, C2 => 
                           n7433, A => n7535, ZN => n7371);
   U518 : XOR2_X1 port map( A => DATA2_I_6_port, B => n9192, Z => n7499);
   U519 : OAI21_X1 port map( B1 => n7434, B2 => n7371, A => n7499, ZN => n7373)
                           ;
   U520 : OAI221_X1 port map( B1 => n7463, B2 => n7435, C1 => n7463, C2 => 
                           n7373, A => n7372, ZN => n8486);
   U521 : NAND2_X1 port map( A1 => n8858, A2 => n8486, ZN => n8451);
   U522 : AOI211_X1 port map( C1 => n7400, C2 => n7620, A => n8556, B => n8451,
                           ZN => n7377);
   U523 : NAND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n7375)
                           ;
   U524 : INV_X1 port map( A => DATA1(8), ZN => n8654);
   U525 : INV_X1 port map( A => DATA2_I_8_port, ZN => n7374);
   U526 : NOR3_X1 port map( A1 => n8654, A2 => n7620, A3 => n7374, ZN => n8545)
                           ;
   U527 : NOR2_X1 port map( A1 => n9190, A2 => n8486, ZN => n8506);
   U528 : INV_X1 port map( A => n8506, ZN => n8543);
   U529 : AOI211_X1 port map( C1 => n7620, C2 => n7375, A => n8545, B => n8543,
                           ZN => n7376);
   U530 : AOI211_X1 port map( C1 => n8848, C2 => n7378, A => n7377, B => n7376,
                           ZN => n7398);
   U531 : NOR2_X1 port map( A1 => n8312, A2 => n8654, ZN => n7441);
   U532 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(7), ZN => n7504);
   U533 : NAND2_X1 port map( A1 => n7832, A2 => DATA1(6), ZN => n7579);
   U534 : NAND2_X1 port map( A1 => DATA1(5), A2 => n7776, ZN => n8325);
   U535 : NAND4_X1 port map( A1 => n7379, A2 => n7504, A3 => n7579, A4 => n8325
                           , ZN => n7380);
   U536 : NOR2_X1 port map( A1 => n7441, A2 => n7380, ZN => n7800);
   U537 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(8), ZN => n7401);
   U538 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(6), ZN => n7542);
   U539 : NAND2_X1 port map( A1 => n8763, A2 => DATA1(5), ZN => n8090);
   U540 : NAND2_X1 port map( A1 => DATA1(4), A2 => n7776, ZN => n8764);
   U541 : AND4_X1 port map( A1 => n7401, A2 => n7542, A3 => n8090, A4 => n8764,
                           ZN => n7381);
   U542 : NAND2_X1 port map( A1 => n7896, A2 => n9193, ZN => n7470);
   U543 : AND2_X1 port map( A1 => n7381, A2 => n7470, ZN => n7802);
   U544 : INV_X1 port map( A => DATA1(5), ZN => n7526);
   U545 : NOR2_X1 port map( A1 => n8130, A2 => n7526, ZN => n7583);
   U546 : INV_X1 port map( A => n9191, ZN => n7575);
   U547 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(6), ZN => n7503);
   U548 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(7), ZN => n7382);
   U549 : OAI211_X1 port map( C1 => n7978, C2 => n7575, A => n7503, B => n7382,
                           ZN => n7383);
   U550 : AOI211_X1 port map( C1 => DATA1(4), C2 => n7832, A => n7583, B => 
                           n7383, ZN => n7392);
   U551 : OAI222_X1 port map( A1 => n7986, A2 => n7800, B1 => n8186, B2 => 
                           n7802, C1 => n7898, C2 => n7392, ZN => n7955);
   U552 : INV_X1 port map( A => n7955, ZN => n8045);
   U553 : NOR2_X1 port map( A1 => n8312, A2 => n7526, ZN => n7544);
   U554 : INV_X1 port map( A => DATA1(2), ZN => n8585);
   U555 : CLKBUF_X1 port map( A => DATA1(4), Z => n8324);
   U556 : NAND2_X1 port map( A1 => n8152, A2 => n8324, ZN => n8088);
   U557 : NAND2_X1 port map( A1 => n8762, A2 => n9192, ZN => n7384);
   U558 : OAI211_X1 port map( C1 => n7978, C2 => n8585, A => n8088, B => n7384,
                           ZN => n7385);
   U559 : AOI211_X1 port map( C1 => n7832, C2 => DATA1(3), A => n7544, B => 
                           n7385, ZN => n7391);
   U560 : OAI222_X1 port map( A1 => n7986, A2 => n7802, B1 => n8186, B2 => 
                           n7392, C1 => n7898, C2 => n7391, ZN => n8041);
   U561 : NOR2_X1 port map( A1 => n7893, A2 => n7526, ZN => n7387);
   U562 : NAND2_X1 port map( A1 => n7896, A2 => n8324, ZN => n7580);
   U563 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(3), ZN => n8327);
   U564 : OAI211_X1 port map( C1 => n7680, C2 => n8585, A => n7580, B => n8327,
                           ZN => n7386);
   U565 : AOI211_X1 port map( C1 => DATA1(1), C2 => n7776, A => n7387, B => 
                           n7386, ZN => n7527);
   U566 : AND2_X1 port map( A1 => n8762, A2 => DATA1(4), ZN => n7389);
   U567 : INV_X1 port map( A => DATA1(1), ZN => n8314);
   U568 : NAND2_X1 port map( A1 => n8153, A2 => n9191, ZN => n8089);
   U569 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(2), ZN => n8766);
   U570 : OAI211_X1 port map( C1 => n7680, C2 => n8314, A => n8089, B => n8766,
                           ZN => n7388);
   U571 : AOI211_X1 port map( C1 => DATA1(0), C2 => n8087, A => n7389, B => 
                           n7388, ZN => n7538);
   U572 : OAI222_X1 port map( A1 => n7986, A2 => n7391, B1 => n8186, B2 => 
                           n7527, C1 => n7898, C2 => n7538, ZN => n8039);
   U573 : AOI22_X1 port map( A1 => n8230, A2 => n8041, B1 => n8335, B2 => n8039
                           , ZN => n7390);
   U574 : OAI21_X1 port map( B1 => n8777, B2 => n8045, A => n7390, ZN => n7394)
                           ;
   U575 : OAI222_X1 port map( A1 => n7986, A2 => n7392, B1 => n8186, B2 => 
                           n7391, C1 => n7898, C2 => n7527, ZN => n8040);
   U576 : NAND2_X1 port map( A1 => n8857, A2 => n7393, ZN => n8547);
   U577 : INV_X1 port map( A => n8547, ZN => n8479);
   U578 : OAI221_X1 port map( B1 => n7394, B2 => n8229, C1 => n7394, C2 => 
                           n8040, A => n8479, ZN => n7397);
   U579 : NAND2_X1 port map( A1 => FUNC(3), A2 => n7395, ZN => n8574);
   U580 : NAND2_X1 port map( A1 => n8857, A2 => n8567, ZN => n8527);
   U581 : NAND2_X1 port map( A1 => n8574, A2 => n8527, ZN => n8505);
   U582 : NAND3_X1 port map( A1 => DATA2(9), A2 => DATA1(9), A3 => n8505, ZN =>
                           n7396);
   U583 : NAND4_X1 port map( A1 => n7399, A2 => n7398, A3 => n7397, A4 => n7396
                           , ZN => OUTALU(9));
   U584 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => DATA1(8), A => n7400, 
                           ZN => n7622);
   U585 : INV_X1 port map( A => n7622, ZN => n7428);
   U586 : OAI22_X1 port map( A1 => n7487, A2 => n8821, B1 => n8552, B2 => n8817
                           , ZN => n7426);
   U587 : INV_X1 port map( A => n8230, ZN => n8778);
   U588 : OAI22_X1 port map( A1 => n8774, A2 => n7473, B1 => n8778, B2 => n7508
                           , ZN => n7407);
   U589 : NOR2_X1 port map( A1 => n8130, A2 => n8599, ZN => n7683);
   U590 : INV_X1 port map( A => n8504, ZN => n8602);
   U591 : NAND2_X1 port map( A1 => n7896, A2 => DATA1(9), ZN => n7726);
   U592 : OAI211_X1 port map( C1 => n7978, C2 => n8602, A => n7401, B => n7726,
                           ZN => n7402);
   U593 : AOI211_X1 port map( C1 => DATA1(11), C2 => n8763, A => n7683, B => 
                           n7402, ZN => n7403);
   U594 : INV_X1 port map( A => n7403, ZN => n7472);
   U595 : AOI222_X1 port map( A1 => n8770, A2 => n7472, B1 => n8768, B2 => 
                           n7444, C1 => n7586, C2 => n7404, ZN => n7548);
   U596 : OAI22_X1 port map( A1 => n8331, A2 => n7405, B1 => n8777, B2 => n7548
                           , ZN => n7406);
   U597 : AOI211_X1 port map( C1 => n7408, C2 => n8335, A => n7407, B => n7406,
                           ZN => n7551);
   U598 : INV_X1 port map( A => n7551, ZN => n7514);
   U599 : AOI22_X1 port map( A1 => n8522, A2 => n7514, B1 => n8524, B2 => n7480
                           , ZN => n7412);
   U600 : AOI22_X1 port map( A1 => n8496, A2 => n7410, B1 => n8339, B2 => n7409
                           , ZN => n7411);
   U601 : OAI211_X1 port map( C1 => n7413, C2 => n8477, A => n7412, B => n7411,
                           ZN => n7469);
   U602 : AOI222_X1 port map( A1 => n7943, A2 => n7451, B1 => n8456, B2 => 
                           n7469, C1 => n7414, C2 => n8051, ZN => n7520);
   U603 : OAI22_X1 port map( A1 => n8463, A2 => n7520, B1 => n7415, B2 => n8814
                           , ZN => n7418);
   U604 : AOI22_X1 port map( A1 => n8809, A2 => n8497, B1 => n7483, B2 => n8807
                           , ZN => n7416);
   U605 : INV_X1 port map( A => n7416, ZN => n7417);
   U606 : AOI211_X1 port map( C1 => n8811, C2 => n7516, A => n7418, B => n7417,
                           ZN => n7559);
   U607 : NAND3_X1 port map( A1 => n8889, A2 => n7420, A3 => n7419, ZN => n8823
                           );
   U608 : OAI22_X1 port map( A1 => n8553, A2 => n7559, B1 => n8551, B2 => n8823
                           , ZN => n7425);
   U609 : AOI222_X1 port map( A1 => n8041, A2 => n8231, B1 => n8040, B2 => 
                           n8230, C1 => n8039, C2 => n8229, ZN => n7423);
   U610 : INV_X1 port map( A => DATA2(8), ZN => n8882);
   U611 : OAI22_X1 port map( A1 => n8654, A2 => n8882, B1 => DATA2(8), B2 => 
                           DATA1(8), ZN => n8739);
   U612 : INV_X1 port map( A => n8739, ZN => n8650);
   U613 : AOI22_X1 port map( A1 => dataout_mul_8_port, A2 => n8575, B1 => n8567
                           , B2 => n8650, ZN => n7422);
   U614 : NAND3_X1 port map( A1 => DATA2(8), A2 => DATA1(8), A3 => n8505, ZN =>
                           n7421);
   U615 : OAI211_X1 port map( C1 => n7423, C2 => n8547, A => n7422, B => n7421,
                           ZN => n7424);
   U616 : AOI221_X1 port map( B1 => n7426, B2 => n8848, C1 => n7425, C2 => 
                           n8848, A => n7424, ZN => n7427);
   U617 : OAI221_X1 port map( B1 => n7622, B2 => n8451, C1 => n7428, C2 => 
                           n8543, A => n7427, ZN => OUTALU(8));
   U618 : INV_X1 port map( A => n7463, ZN => n7465);
   U619 : NOR2_X1 port map( A1 => n9190, A2 => cin, ZN => n8084);
   U620 : INV_X1 port map( A => n8319, ZN => n8315);
   U621 : INV_X1 port map( A => n7429, ZN => n7430);
   U622 : AOI21_X1 port map( B1 => n8316, B2 => n8315, A => n7430, ZN => n8083)
                           ;
   U623 : OAI21_X1 port map( B1 => n8083, B2 => n8125, A => n7431, ZN => n7578)
                           ;
   U624 : AOI21_X1 port map( B1 => n7611, B2 => n7578, A => n7432, ZN => n7567)
                           ;
   U625 : OAI21_X1 port map( B1 => n7567, B2 => n7572, A => n7433, ZN => n7501)
                           ;
   U626 : INV_X1 port map( A => n7535, ZN => n7537);
   U627 : AOI21_X1 port map( B1 => n7501, B2 => n7537, A => n7434, ZN => n7468)
                           ;
   U628 : INV_X1 port map( A => n7499, ZN => n7497);
   U629 : OAI21_X1 port map( B1 => n7468, B2 => n7497, A => n7435, ZN => n7437)
                           ;
   U630 : NAND2_X1 port map( A1 => n8858, A2 => cin, ZN => n8317);
   U631 : INV_X1 port map( A => n8317, ZN => n8572);
   U632 : NOR2_X1 port map( A1 => n7430, A2 => n8318, ZN => n8082);
   U633 : OAI21_X1 port map( B1 => n8082, B2 => n8125, A => n7431, ZN => n7577)
                           ;
   U634 : AOI21_X1 port map( B1 => n7611, B2 => n7577, A => n7432, ZN => n7566)
                           ;
   U635 : OAI21_X1 port map( B1 => n7566, B2 => n7572, A => n7433, ZN => n7500)
                           ;
   U636 : AOI21_X1 port map( B1 => n7500, B2 => n7537, A => n7434, ZN => n7467)
                           ;
   U637 : OAI21_X1 port map( B1 => n7467, B2 => n7497, A => n7435, ZN => n7436)
                           ;
   U638 : AOI22_X1 port map( A1 => n8084, A2 => n7437, B1 => n8572, B2 => n7436
                           , ZN => n7464);
   U639 : INV_X1 port map( A => n8084, ZN => n8568);
   U640 : OAI22_X1 port map( A1 => n8568, A2 => n7437, B1 => n8317, B2 => n7436
                           , ZN => n7438);
   U641 : INV_X1 port map( A => n7438, ZN => n7462);
   U642 : CLKBUF_X1 port map( A => n8514, Z => n8530);
   U643 : INV_X1 port map( A => n8817, ZN => n8239);
   U644 : INV_X1 port map( A => n7520, ZN => n7556);
   U645 : AOI22_X1 port map( A1 => n8500, A2 => n7483, B1 => n8809, B2 => n7440
                           , ZN => n7453);
   U646 : AOI22_X1 port map( A1 => n9193, A2 => n8323, B1 => DATA1(11), B2 => 
                           n8087, ZN => n7443);
   U647 : INV_X1 port map( A => n7441, ZN => n7442);
   U648 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(9), ZN => n7686);
   U649 : NAND2_X1 port map( A1 => n7832, A2 => DATA1(10), ZN => n7675);
   U650 : NAND4_X1 port map( A1 => n7443, A2 => n7442, A3 => n7686, A4 => n7675
                           , ZN => n7507);
   U651 : AOI222_X1 port map( A1 => n7444, A2 => n8772, B1 => n7507, B2 => 
                           n8770, C1 => n7472, C2 => n8768, ZN => n7547);
   U652 : INV_X1 port map( A => n7547, ZN => n7590);
   U653 : OAI22_X1 port map( A1 => n7473, A2 => n8780, B1 => n7548, B2 => n8044
                           , ZN => n7447);
   U654 : OAI22_X1 port map( A1 => n7445, A2 => n8331, B1 => n7508, B2 => n8774
                           , ZN => n7446);
   U655 : AOI211_X1 port map( C1 => n8203, C2 => n7590, A => n7447, B => n7446,
                           ZN => n7591);
   U656 : INV_X1 port map( A => n7591, ZN => n7554);
   U657 : AOI22_X1 port map( A1 => n8522, A2 => n7554, B1 => n8524, B2 => n7514
                           , ZN => n7450);
   U658 : AOI22_X1 port map( A1 => n8496, A2 => n7480, B1 => n7995, B2 => n7448
                           , ZN => n7449);
   U659 : OAI211_X1 port map( C1 => n7477, C2 => n8477, A => n7450, B => n7449,
                           ZN => n7481);
   U660 : AOI222_X1 port map( A1 => n7451, A2 => n8051, B1 => n7469, B2 => 
                           n7943, C1 => n7481, C2 => n8456, ZN => n7597);
   U661 : INV_X1 port map( A => n7597, ZN => n7517);
   U662 : AOI22_X1 port map( A1 => n8807, A2 => n7516, B1 => n8485, B2 => n7517
                           , ZN => n7452);
   U663 : NAND2_X1 port map( A1 => n7453, A2 => n7452, ZN => n7601);
   U664 : AOI21_X1 port map( B1 => n8811, B2 => n7556, A => n7601, ZN => n7560)
                           ;
   U665 : OAI22_X1 port map( A1 => n8553, A2 => n7560, B1 => n7559, B2 => n8821
                           , ZN => n7455);
   U666 : OAI22_X1 port map( A1 => n8552, A2 => n8823, B1 => n8551, B2 => n8819
                           , ZN => n7454);
   U667 : AOI211_X1 port map( C1 => n8239, C2 => n7523, A => n7455, B => n7454,
                           ZN => n7524);
   U668 : NOR3_X1 port map( A1 => n8832, A2 => n7524, A3 => n8536, ZN => n7460)
                           ;
   U669 : AOI22_X1 port map( A1 => n7919, A2 => n8039, B1 => n8203, B2 => n8040
                           , ZN => n7458);
   U670 : INV_X1 port map( A => DATA1(7), ZN => n7581);
   U671 : NOR2_X1 port map( A1 => DATA2(7), A2 => n7581, ZN => n8651);
   U672 : INV_X1 port map( A => DATA2(7), ZN => n8885);
   U673 : NOR2_X1 port map( A1 => DATA1(7), A2 => n8885, ZN => n8633);
   U674 : OAI21_X1 port map( B1 => n8651, B2 => n8633, A => n8567, ZN => n7457)
                           ;
   U675 : NAND3_X1 port map( A1 => DATA2(7), A2 => n9193, A3 => n8505, ZN => 
                           n7456);
   U676 : OAI211_X1 port map( C1 => n7458, C2 => n8547, A => n7457, B => n7456,
                           ZN => n7459);
   U677 : AOI211_X1 port map( C1 => n8530, C2 => dataout_mul_7_port, A => n7460
                           , B => n7459, ZN => n7461);
   U678 : OAI221_X1 port map( B1 => n7465, B2 => n7464, C1 => n7463, C2 => 
                           n7462, A => n7461, ZN => OUTALU(7));
   U679 : OAI22_X1 port map( A1 => n8568, A2 => n7468, B1 => n8317, B2 => n7467
                           , ZN => n7466);
   U680 : INV_X1 port map( A => n7466, ZN => n7498);
   U681 : AOI22_X1 port map( A1 => n8084, A2 => n7468, B1 => n8572, B2 => n7467
                           , ZN => n7496);
   U682 : INV_X1 port map( A => n8103, ZN => n8383);
   U683 : INV_X1 port map( A => n7469, ZN => n7482);
   U684 : INV_X1 port map( A => n7508, ZN => n7476);
   U685 : AOI22_X1 port map( A1 => n7832, A2 => DATA1(9), B1 => n8762, B2 => 
                           DATA1(6), ZN => n7471);
   U686 : NAND2_X1 port map( A1 => n8152, A2 => DATA1(8), ZN => n7725);
   U687 : NAND2_X1 port map( A1 => DATA1(10), A2 => n8087, ZN => n7689);
   U688 : NAND4_X1 port map( A1 => n7471, A2 => n7470, A3 => n7725, A4 => n7689
                           , ZN => n7546);
   U689 : AOI222_X1 port map( A1 => n7472, A2 => n8772, B1 => n7546, B2 => 
                           n8770, C1 => n7507, C2 => n8768, ZN => n7587);
   U690 : OAI22_X1 port map( A1 => n8777, A2 => n7587, B1 => n7548, B2 => n8774
                           , ZN => n7475);
   U691 : OAI22_X1 port map( A1 => n7473, A2 => n8331, B1 => n7547, B2 => n8778
                           , ZN => n7474);
   U692 : AOI211_X1 port map( C1 => n8335, C2 => n7476, A => n7475, B => n7474,
                           ZN => n8097);
   U693 : OAI22_X1 port map( A1 => n7591, A2 => n8790, B1 => n8097, B2 => n8786
                           , ZN => n7479);
   U694 : OAI22_X1 port map( A1 => n7551, A2 => n8788, B1 => n8793, B2 => n7477
                           , ZN => n7478);
   U695 : AOI211_X1 port map( C1 => n8100, C2 => n7480, A => n7479, B => n7478,
                           ZN => n7555);
   U696 : INV_X1 port map( A => n7481, ZN => n7515);
   U697 : OAI222_X1 port map( A1 => n7482, A2 => n8101, B1 => n7555, B2 => 
                           n7862, C1 => n7515, C2 => n8803, ZN => n8104);
   U698 : AOI22_X1 port map( A1 => n8811, A2 => n7517, B1 => n8805, B2 => n8104
                           , ZN => n7485);
   U699 : AOI22_X1 port map( A1 => n8500, A2 => n7516, B1 => n8809, B2 => n7483
                           , ZN => n7484);
   U700 : OAI211_X1 port map( C1 => n7520, C2 => n8383, A => n7485, B => n7484,
                           ZN => n8110);
   U701 : OAI22_X1 port map( A1 => n7560, A2 => n8821, B1 => n7486, B2 => n8819
                           , ZN => n7489);
   U702 : OAI22_X1 port map( A1 => n7487, A2 => n8823, B1 => n7559, B2 => n8817
                           , ZN => n7488);
   U703 : AOI211_X1 port map( C1 => n8828, C2 => n8110, A => n7489, B => n7488,
                           ZN => n7564);
   U704 : OAI211_X1 port map( C1 => DATA2(2), C2 => DATA2(1), A => DATA2(3), B 
                           => DATA2(4), ZN => n8829);
   U705 : NAND2_X1 port map( A1 => n8829, A2 => n8832, ZN => n8834);
   U706 : OAI22_X1 port map( A1 => n8832, A2 => n7564, B1 => n7524, B2 => n8834
                           , ZN => n7494);
   U707 : INV_X1 port map( A => DATA2(6), ZN => n8886);
   U708 : INV_X1 port map( A => n9192, ZN => n8634);
   U709 : AOI22_X1 port map( A1 => n9192, A2 => n8886, B1 => DATA2(6), B2 => 
                           n8634, ZN => n8649);
   U710 : OAI21_X1 port map( B1 => n8574, B2 => n8634, A => n8527, ZN => n7490)
                           ;
   U711 : AOI22_X1 port map( A1 => DATA2(6), A2 => n7490, B1 => n8530, B2 => 
                           dataout_mul_6_port, ZN => n7492);
   U712 : NAND3_X1 port map( A1 => n8479, A2 => n8203, A3 => n8039, ZN => n7491
                           );
   U713 : OAI211_X1 port map( C1 => n8649, C2 => n8525, A => n7492, B => n7491,
                           ZN => n7493);
   U714 : AOI21_X1 port map( B1 => n8848, B2 => n7494, A => n7493, ZN => n7495)
                           ;
   U715 : OAI221_X1 port map( B1 => n7499, B2 => n7498, C1 => n7497, C2 => 
                           n7496, A => n7495, ZN => OUTALU(6));
   U716 : AOI22_X1 port map( A1 => n8084, A2 => n7501, B1 => n8572, B2 => n7500
                           , ZN => n7536);
   U717 : OAI22_X1 port map( A1 => n8568, A2 => n7501, B1 => n8317, B2 => n7500
                           , ZN => n7502);
   U718 : INV_X1 port map( A => n7502, ZN => n7534);
   U719 : OAI21_X1 port map( B1 => n8574, B2 => n7526, A => n8527, ZN => n7532)
                           ;
   U720 : INV_X1 port map( A => n7587, ZN => n8096);
   U721 : AOI22_X1 port map( A1 => n7832, A2 => DATA1(8), B1 => n8762, B2 => 
                           DATA1(5), ZN => n7505);
   U722 : NAND2_X1 port map( A1 => DATA1(9), A2 => n8087, ZN => n7674);
   U723 : NAND4_X1 port map( A1 => n7505, A2 => n7504, A3 => n7503, A4 => n7674
                           , ZN => n7585);
   U724 : AOI222_X1 port map( A1 => n7507, A2 => n8772, B1 => n7585, B2 => 
                           n8770, C1 => n7546, C2 => n7506, ZN => n8332);
   U725 : OAI22_X1 port map( A1 => n8777, A2 => n8332, B1 => n7547, B2 => n8330
                           , ZN => n7510);
   U726 : OAI22_X1 port map( A1 => n7508, A2 => n8331, B1 => n7548, B2 => n8780
                           , ZN => n7509);
   U727 : AOI211_X1 port map( C1 => n7919, C2 => n8096, A => n7510, B => n7509,
                           ZN => n8086);
   U728 : OAI22_X1 port map( A1 => n8097, A2 => n8790, B1 => n8086, B2 => n8786
                           , ZN => n7513);
   U729 : OAI22_X1 port map( A1 => n8793, A2 => n7511, B1 => n7591, B2 => n8788
                           , ZN => n7512);
   U730 : AOI211_X1 port map( C1 => n8100, C2 => n7514, A => n7513, B => n7512,
                           ZN => n7595);
   U731 : OAI222_X1 port map( A1 => n7515, A2 => n8101, B1 => n7555, B2 => 
                           n8803, C1 => n7595, C2 => n8801, ZN => n8342);
   U732 : AOI22_X1 port map( A1 => n8811, A2 => n8104, B1 => n8805, B2 => n8342
                           , ZN => n7519);
   U733 : AOI22_X1 port map( A1 => n8807, A2 => n7517, B1 => n8809, B2 => n7516
                           , ZN => n7518);
   U734 : OAI211_X1 port map( C1 => n7520, C2 => n8814, A => n7519, B => n7518,
                           ZN => n8108);
   U735 : INV_X1 port map( A => n8108, ZN => n8348);
   U736 : OAI22_X1 port map( A1 => n8553, A2 => n8348, B1 => n7560, B2 => n8817
                           , ZN => n7522);
   U737 : INV_X1 port map( A => n8110, ZN => n7561);
   U738 : OAI22_X1 port map( A1 => n7561, A2 => n8821, B1 => n7559, B2 => n8823
                           , ZN => n7521);
   U739 : AOI211_X1 port map( C1 => n8111, C2 => n7523, A => n7522, B => n7521,
                           ZN => n7605);
   U740 : CLKBUF_X1 port map( A => n8829, Z => n8060);
   U741 : OAI222_X1 port map( A1 => n8834, A2 => n7564, B1 => n8832, B2 => 
                           n7605, C1 => n7524, C2 => n8060, ZN => n8353);
   U742 : OAI21_X1 port map( B1 => n8888, B2 => n7525, A => n8021, ZN => n8064)
                           ;
   U743 : INV_X1 port map( A => n8064, ZN => n8838);
   U744 : AND3_X1 port map( A1 => n8353, A2 => n8848, A3 => n8838, ZN => n7531)
                           ;
   U745 : INV_X1 port map( A => DATA2(5), ZN => n8887);
   U746 : NAND2_X1 port map( A1 => n8887, A2 => DATA1(5), ZN => n8648);
   U747 : NAND2_X1 port map( A1 => DATA2(5), A2 => n7526, ZN => n8644);
   U748 : AND2_X1 port map( A1 => n8648, A2 => n8644, ZN => n8746);
   U749 : OAI22_X1 port map( A1 => n7527, A2 => n7986, B1 => n7538, B2 => n7984
                           , ZN => n7528);
   U750 : AOI22_X1 port map( A1 => n8575, A2 => dataout_mul_5_port, B1 => n8479
                           , B2 => n7528, ZN => n7529);
   U751 : OAI21_X1 port map( B1 => n8746, B2 => n8525, A => n7529, ZN => n7530)
                           ;
   U752 : AOI211_X1 port map( C1 => DATA2(5), C2 => n7532, A => n7531, B => 
                           n7530, ZN => n7533);
   U753 : OAI221_X1 port map( B1 => n7537, B2 => n7536, C1 => n7535, C2 => 
                           n7534, A => n7533, ZN => OUTALU(5));
   U754 : AOI22_X1 port map( A1 => n8084, A2 => n7567, B1 => n8572, B2 => n7566
                           , ZN => n7573);
   U755 : NOR3_X1 port map( A1 => n7538, A2 => n8547, A3 => n7224, ZN => n7541)
                           ;
   U756 : NOR2_X1 port map( A1 => n8888, A2 => n8324, ZN => n8589);
   U757 : INV_X1 port map( A => n8589, ZN => n8645);
   U758 : NAND2_X1 port map( A1 => n8324, A2 => n8888, ZN => n8642);
   U759 : NAND3_X1 port map( A1 => n8324, A2 => DATA2(4), A3 => n8505, ZN => 
                           n7539);
   U760 : OAI221_X1 port map( B1 => n8525, B2 => n8645, C1 => n8525, C2 => 
                           n8642, A => n7539, ZN => n7540);
   U761 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n8530, A => n7541
                           , B => n7540, ZN => n7571);
   U762 : INV_X1 port map( A => n8342, ZN => n7596);
   U763 : NAND2_X1 port map( A1 => n8763, A2 => n9193, ZN => n7724);
   U764 : OAI211_X1 port map( C1 => n7978, C2 => n8654, A => n7542, B => n7724,
                           ZN => n7543);
   U765 : AOI211_X1 port map( C1 => n8323, C2 => n8324, A => n7544, B => n7543,
                           ZN => n7545);
   U766 : INV_X1 port map( A => n7545, ZN => n8092);
   U767 : AOI222_X1 port map( A1 => n8770, A2 => n8092, B1 => n8768, B2 => 
                           n7585, C1 => n7586, C2 => n7546, ZN => n8093);
   U768 : INV_X1 port map( A => n8093, ZN => n8784);
   U769 : OAI22_X1 port map( A1 => n7547, A2 => n8780, B1 => n8332, B2 => n8778
                           , ZN => n7550);
   U770 : OAI22_X1 port map( A1 => n7548, A2 => n8331, B1 => n7587, B2 => n8774
                           , ZN => n7549);
   U771 : AOI211_X1 port map( C1 => n8203, C2 => n8784, A => n7550, B => n7549,
                           ZN => n8792);
   U772 : OAI22_X1 port map( A1 => n8792, A2 => n8786, B1 => n8086, B2 => n8790
                           , ZN => n7553);
   U773 : OAI22_X1 port map( A1 => n8793, A2 => n7551, B1 => n8097, B2 => n8788
                           , ZN => n7552);
   U774 : AOI211_X1 port map( C1 => n8100, C2 => n7554, A => n7553, B => n7552,
                           ZN => n8102);
   U775 : OAI222_X1 port map( A1 => n8803, A2 => n7595, B1 => n7862, B2 => 
                           n8102, C1 => n7555, C2 => n8798, ZN => n8808);
   U776 : AOI22_X1 port map( A1 => n8807, A2 => n8104, B1 => n8809, B2 => n7556
                           , ZN => n7557);
   U777 : OAI21_X1 port map( B1 => n7597, B2 => n8814, A => n7557, ZN => n7558)
                           ;
   U778 : AOI21_X1 port map( B1 => n8485, B2 => n8808, A => n7558, ZN => n8820)
                           ;
   U779 : OAI21_X1 port map( B1 => n7596, B2 => n8461, A => n8820, ZN => n8107)
                           ;
   U780 : INV_X1 port map( A => n8107, ZN => n8347);
   U781 : OAI22_X1 port map( A1 => n8553, A2 => n8347, B1 => n7559, B2 => n8819
                           , ZN => n7563);
   U782 : OAI22_X1 port map( A1 => n7561, A2 => n8817, B1 => n7560, B2 => n8823
                           , ZN => n7562);
   U783 : AOI211_X1 port map( C1 => n8351, C2 => n8108, A => n7563, B => n7562,
                           ZN => n8115);
   U784 : OAI222_X1 port map( A1 => n8834, A2 => n7605, B1 => n8832, B2 => 
                           n8115, C1 => n7564, C2 => n8060, ZN => n8841);
   U785 : NAND2_X1 port map( A1 => n8021, A2 => n8064, ZN => n8845);
   U786 : INV_X1 port map( A => n8845, ZN => n8167);
   U787 : AOI22_X1 port map( A1 => n8841, A2 => n8838, B1 => n8353, B2 => n8167
                           , ZN => n7565);
   U788 : INV_X1 port map( A => n7565, ZN => n7569);
   U789 : OAI22_X1 port map( A1 => n7567, A2 => n8568, B1 => n7566, B2 => n8317
                           , ZN => n7568);
   U790 : AOI22_X1 port map( A1 => n8848, A2 => n7569, B1 => n7572, B2 => n7568
                           , ZN => n7570);
   U791 : OAI211_X1 port map( C1 => n7573, C2 => n7572, A => n7571, B => n7570,
                           ZN => OUTALU(4));
   U792 : AOI22_X1 port map( A1 => n8152, A2 => DATA1(1), B1 => n8763, B2 => 
                           DATA1(0), ZN => n7574);
   U793 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(2), ZN => n8326);
   U794 : OAI211_X1 port map( C1 => n7575, C2 => n7893, A => n7574, B => n8326,
                           ZN => n7576);
   U795 : AOI22_X1 port map( A1 => n8530, A2 => dataout_mul_3_port, B1 => n8479
                           , B2 => n7576, ZN => n7615);
   U796 : OAI22_X1 port map( A1 => n8568, A2 => n7578, B1 => n8317, B2 => n7577
                           , ZN => n7610);
   U797 : AOI22_X1 port map( A1 => n8084, A2 => n7578, B1 => n8572, B2 => n7577
                           , ZN => n7608);
   U798 : INV_X1 port map( A => n8792, ZN => n7594);
   U799 : OAI211_X1 port map( C1 => n7978, C2 => n7581, A => n7580, B => n7579,
                           ZN => n7582);
   U800 : AOI211_X1 port map( C1 => n8323, C2 => DATA1(3), A => n7583, B => 
                           n7582, ZN => n7584);
   U801 : INV_X1 port map( A => n7584, ZN => n8329);
   U802 : AOI222_X1 port map( A1 => n8770, A2 => n8329, B1 => n8768, B2 => 
                           n8092, C1 => n7586, C2 => n7585, ZN => n8781);
   U803 : OAI22_X1 port map( A1 => n8330, A2 => n8332, B1 => n8777, B2 => n8781
                           , ZN => n7589);
   U804 : OAI22_X1 port map( A1 => n8778, A2 => n8093, B1 => n8780, B2 => n7587
                           , ZN => n7588);
   U805 : AOI211_X1 port map( C1 => n7590, C2 => n8785, A => n7589, B => n7588,
                           ZN => n8761);
   U806 : OAI22_X1 port map( A1 => n8477, A2 => n8097, B1 => n8786, B2 => n8761
                           , ZN => n7593);
   U807 : OAI22_X1 port map( A1 => n8788, A2 => n8086, B1 => n8793, B2 => n7591
                           , ZN => n7592);
   U808 : AOI211_X1 port map( C1 => n7594, C2 => n8524, A => n7593, B => n7592,
                           ZN => n8340);
   U809 : OAI222_X1 port map( A1 => n7595, A2 => n8101, B1 => n8102, B2 => 
                           n8803, C1 => n8340, C2 => n8801, ZN => n8341);
   U810 : INV_X1 port map( A => n8341, ZN => n8815);
   U811 : OAI22_X1 port map( A1 => n7596, A2 => n8383, B1 => n8463, B2 => n8815
                           , ZN => n7600);
   U812 : INV_X1 port map( A => n8104, ZN => n7598);
   U813 : OAI22_X1 port map( A1 => n7598, A2 => n8814, B1 => n8052, B2 => n7597
                           , ZN => n7599);
   U814 : AOI211_X1 port map( C1 => n8811, C2 => n8808, A => n7600, B => n7599,
                           ZN => n8824);
   U815 : AOI22_X1 port map( A1 => n8111, A2 => n7601, B1 => n8351, B2 => n8107
                           , ZN => n7603);
   U816 : INV_X1 port map( A => n8823, ZN => n8109);
   U817 : AOI22_X1 port map( A1 => n8109, A2 => n8110, B1 => n8239, B2 => n8108
                           , ZN => n7602);
   U818 : OAI211_X1 port map( C1 => n8553, C2 => n8824, A => n7603, B => n7602,
                           ZN => n7604);
   U819 : INV_X1 port map( A => n7604, ZN => n8352);
   U820 : OAI222_X1 port map( A1 => n8834, A2 => n8115, B1 => n8352, B2 => 
                           n8832, C1 => n7605, C2 => n8829, ZN => n8839);
   U821 : NOR2_X1 port map( A1 => n8021, A2 => n7606, ZN => n8836);
   U822 : AOI222_X1 port map( A1 => n8839, A2 => n8838, B1 => n8841, B2 => 
                           n8167, C1 => n8353, C2 => n8836, ZN => n7607);
   U823 : OAI22_X1 port map( A1 => n7611, A2 => n7608, B1 => n7607, B2 => n8536
                           , ZN => n7609);
   U824 : AOI21_X1 port map( B1 => n7611, B2 => n7610, A => n7609, ZN => n7614)
                           ;
   U825 : NAND3_X1 port map( A1 => n9191, A2 => DATA2(3), A3 => n8505, ZN => 
                           n7613);
   U826 : NAND2_X1 port map( A1 => n8889, A2 => DATA1(3), ZN => n8643);
   U827 : INV_X1 port map( A => n8643, ZN => n8586);
   U828 : NOR2_X1 port map( A1 => n8889, A2 => DATA1(3), ZN => n8639);
   U829 : OAI21_X1 port map( B1 => n8586, B2 => n8639, A => n8567, ZN => n7612)
                           ;
   U830 : NAND4_X1 port map( A1 => n7615, A2 => n7614, A3 => n7613, A4 => n7612
                           , ZN => OUTALU(3));
   U831 : NAND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => 
                           n8071);
   U832 : INV_X1 port map( A => n8071, ZN => n7616);
   U833 : XOR2_X1 port map( A => DATA2_I_30_port, B => DATA1(30), Z => n8080);
   U834 : AOI22_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, B1 => 
                           n7616, B2 => n8080, ZN => n7632);
   U835 : XOR2_X1 port map( A => DATA2_I_23_port, B => DATA1(23), Z => n8250);
   U836 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n8255);
   U837 : OAI21_X1 port map( B1 => DATA1(22), B2 => DATA2_I_22_port, A => n8255
                           , ZN => n8264);
   U838 : XOR2_X1 port map( A => DATA2_I_21_port, B => n8286, Z => n8297);
   U839 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n7617);
   U840 : INV_X1 port map( A => n7617, ZN => n8245);
   U841 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n8401);
   U842 : INV_X1 port map( A => n8401, ZN => n8421);
   U843 : XOR2_X1 port map( A => DATA2_I_17_port, B => n8403, Z => n8413);
   U844 : AOI22_X1 port map( A1 => n8403, A2 => DATA2_I_17_port, B1 => n8421, 
                           B2 => n8413, ZN => n8381);
   U845 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n8243);
   U846 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => n8243
                           , ZN => n8397);
   U847 : OAI21_X1 port map( B1 => n8381, B2 => n8397, A => n8243, ZN => n8362)
                           ;
   U848 : OAI22_X1 port map( A1 => n8365, A2 => DATA2_I_19_port, B1 => n8245, 
                           B2 => n8362, ZN => n8299);
   U849 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n8246);
   U850 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => n8246
                           , ZN => n8309);
   U851 : OAI21_X1 port map( B1 => n8299, B2 => n8309, A => n8246, ZN => n8282)
                           ;
   U852 : AOI22_X1 port map( A1 => n8286, A2 => DATA2_I_21_port, B1 => n8297, 
                           B2 => n8282, ZN => n8251);
   U853 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => n8420
                           );
   U854 : INV_X1 port map( A => n8413, ZN => n8411);
   U855 : NOR2_X1 port map( A1 => n8420, A2 => n8411, ZN => n8241);
   U856 : INV_X1 port map( A => n8297, ZN => n8295);
   U857 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => n7617
                           , ZN => n8374);
   U858 : NOR4_X1 port map( A1 => n8397, A2 => n8309, A3 => n8295, A4 => n8374,
                           ZN => n7625);
   U859 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n7623);
   U860 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => n7623
                           , ZN => n8446);
   U861 : XOR2_X1 port map( A => DATA2_I_14_port, B => n9195, Z => n8473);
   U862 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n8467);
   U863 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => n8467
                           , ZN => n8492);
   U864 : NAND2_X1 port map( A1 => n8504, A2 => DATA2_I_12_port, ZN => n8493);
   U865 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => n8493
                           , ZN => n8508);
   U866 : NOR2_X1 port map( A1 => n8492, A2 => n8508, ZN => n8444);
   U867 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => n8442
                           );
   U868 : AND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n8561);
   U869 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n8440);
   U870 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => n8440
                           , ZN => n7619);
   U871 : INV_X1 port map( A => n7619, ZN => n8560);
   U872 : OAI21_X1 port map( B1 => n8561, B2 => n8545, A => n8560, ZN => n7618)
                           ;
   U873 : INV_X1 port map( A => n7618, ZN => n8544);
   U874 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => DATA1(10), A => n8544
                           , ZN => n8535);
   U875 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n8441);
   U876 : OAI21_X1 port map( B1 => n8442, B2 => n8535, A => n8441, ZN => n8507)
                           ;
   U877 : NOR2_X1 port map( A1 => n8493, A2 => n8492, ZN => n8443);
   U878 : AOI21_X1 port map( B1 => n8444, B2 => n8507, A => n8443, ZN => n8465)
                           ;
   U879 : NAND2_X1 port map( A1 => n8465, A2 => n8467, ZN => n8452);
   U880 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n8473, B2 => n8452, ZN => n8433);
   U881 : INV_X1 port map( A => n8473, ZN => n8466);
   U882 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => n8441
                           , ZN => n8534);
   U883 : NOR4_X1 port map( A1 => n8466, A2 => n7620, A3 => n7619, A4 => n8534,
                           ZN => n7621);
   U884 : NAND4_X1 port map( A1 => n8444, A2 => n7622, A3 => n7621, A4 => n8486
                           , ZN => n7624);
   U885 : OAI221_X1 port map( B1 => n8446, B2 => n8433, C1 => n8446, C2 => 
                           n7624, A => n7623, ZN => n8248);
   U886 : NAND3_X1 port map( A1 => n8241, A2 => n7625, A3 => n8248, ZN => n7626
                           );
   U887 : OAI221_X1 port map( B1 => n8264, B2 => n8251, C1 => n8264, C2 => 
                           n7626, A => n8255, ZN => n7627);
   U888 : AOI22_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, B1 => 
                           n8250, B2 => n7627, ZN => n7628);
   U889 : NOR2_X1 port map( A1 => n7628, A2 => n9190, ZN => n8224);
   U890 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n8136);
   U891 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n8151);
   U892 : INV_X1 port map( A => n8151, ZN => n8161);
   U893 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n8183);
   U894 : INV_X1 port map( A => n8183, ZN => n7629);
   U895 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => n8225
                           );
   U896 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => n8183
                           , ZN => n8201);
   U897 : NOR2_X1 port map( A1 => n8225, A2 => n8201, ZN => n8182);
   U898 : NOR2_X1 port map( A1 => n7629, A2 => n8182, ZN => n8185);
   U899 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n7630);
   U900 : OAI21_X1 port map( B1 => DATA1(26), B2 => DATA2_I_26_port, A => n7630
                           , ZN => n8197);
   U901 : OAI21_X1 port map( B1 => n8185, B2 => n8197, A => n7630, ZN => n8170)
                           ;
   U902 : NOR2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => n8160
                           );
   U903 : OAI21_X1 port map( B1 => DATA1(28), B2 => DATA2_I_28_port, A => n8136
                           , ZN => n8163);
   U904 : NOR2_X1 port map( A1 => n8160, A2 => n8163, ZN => n7631);
   U905 : OAI21_X1 port map( B1 => n8161, B2 => n8170, A => n7631, ZN => n8149)
                           ;
   U906 : OAI21_X1 port map( B1 => DATA1(29), B2 => DATA2_I_29_port, A => n8071
                           , ZN => n8143);
   U907 : AOI21_X1 port map( B1 => n8136, B2 => n8149, A => n8143, ZN => n7634)
                           ;
   U908 : NAND2_X1 port map( A1 => n8858, A2 => n7628, ZN => n8199);
   U909 : INV_X1 port map( A => n8199, ZN => n8218);
   U910 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n8216);
   U911 : NOR2_X1 port map( A1 => n8201, A2 => n8216, ZN => n8200);
   U912 : NOR2_X1 port map( A1 => n7629, A2 => n8200, ZN => n8184);
   U913 : OAI21_X1 port map( B1 => n8184, B2 => n8197, A => n7630, ZN => n8169)
                           ;
   U914 : OAI21_X1 port map( B1 => n8161, B2 => n8169, A => n7631, ZN => n8148)
                           ;
   U915 : AOI21_X1 port map( B1 => n8136, B2 => n8148, A => n8143, ZN => n7633)
                           ;
   U916 : AOI22_X1 port map( A1 => n8224, A2 => n7634, B1 => n8218, B2 => n7633
                           , ZN => n8079);
   U917 : INV_X1 port map( A => n8080, ZN => n8070);
   U918 : OAI22_X1 port map( A1 => n7632, A2 => n9190, B1 => n8079, B2 => n8070
                           , ZN => n8027);
   U919 : INV_X1 port map( A => n8224, ZN => n8202);
   U920 : OAI22_X1 port map( A1 => n7634, A2 => n8202, B1 => n7633, B2 => n8199
                           , ZN => n8134);
   U921 : AOI22_X1 port map( A1 => n8858, A2 => n8070, B1 => n8071, B2 => n8134
                           , ZN => n8069);
   U922 : AND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => n7635
                           );
   U923 : AOI211_X1 port map( C1 => DATA1(31), C2 => DATA2_I_31_port, A => 
                           n8069, B => n7635, ZN => n8029);
   U924 : INV_X1 port map( A => DATA2(31), ZN => n8859);
   U925 : NAND2_X1 port map( A1 => n8323, A2 => n8848, ZN => n8147);
   U926 : OAI21_X1 port map( B1 => n8574, B2 => n8859, A => n8147, ZN => n7636)
                           ;
   U927 : AOI211_X1 port map( C1 => DATA2_I_31_port, C2 => n8027, A => n8029, B
                           => n7636, ZN => n8068);
   U928 : AOI22_X1 port map( A1 => n7832, A2 => n9195, B1 => n9194, B2 => n7776
                           , ZN => n7640);
   U929 : NAND2_X1 port map( A1 => n8762, A2 => DATA1(17), ZN => n7637);
   U930 : AND4_X1 port map( A1 => n7640, A2 => n7639, A3 => n7638, A4 => n7637,
                           ZN => n7660);
   U931 : NAND4_X1 port map( A1 => n7644, A2 => n7643, A3 => n7642, A4 => n7641
                           , ZN => n7645);
   U932 : AOI21_X1 port map( B1 => n8762, B2 => n8365, A => n7645, ZN => n7671)
                           ;
   U933 : AND3_X1 port map( A1 => n7648, A2 => n7647, A3 => n7646, ZN => n7650)
                           ;
   U934 : OAI211_X1 port map( C1 => n7978, C2 => n8454, A => n7650, B => n7649,
                           ZN => n7651);
   U935 : INV_X1 port map( A => n7651, ZN => n7665);
   U936 : OAI222_X1 port map( A1 => n7660, A2 => n7898, B1 => n7671, B2 => 
                           n7224, C1 => n7665, C2 => n7984, ZN => n7746);
   U937 : INV_X1 port map( A => n7746, ZN => n7718);
   U938 : NAND2_X1 port map( A1 => n8504, A2 => n7776, ZN => n7652);
   U939 : OAI211_X1 port map( C1 => n8474, C2 => n7680, A => n7653, B => n7652,
                           ZN => n7654);
   U940 : AOI211_X1 port map( C1 => n8762, C2 => DATA1(16), A => n7655, B => 
                           n7654, ZN => n7696);
   U941 : NOR2_X1 port map( A1 => n8434, A2 => n7893, ZN => n7659);
   U942 : OAI211_X1 port map( C1 => n7978, C2 => n8526, A => n7657, B => n7656,
                           ZN => n7658);
   U943 : AOI211_X1 port map( C1 => DATA1(12), C2 => n7832, A => n7659, B => 
                           n7658, ZN => n7695);
   U944 : OAI222_X1 port map( A1 => n7986, A2 => n7660, B1 => n8186, B2 => 
                           n7696, C1 => n7898, C2 => n7695, ZN => n7694);
   U945 : OAI222_X1 port map( A1 => n7986, A2 => n7665, B1 => n8186, B2 => 
                           n7660, C1 => n7982, C2 => n7696, ZN => n7701);
   U946 : AOI22_X1 port map( A1 => n8785, A2 => n7694, B1 => n8335, B2 => n7701
                           , ZN => n7673);
   U947 : INV_X1 port map( A => DATA1(16), ZN => n8671);
   U948 : NOR2_X1 port map( A1 => n7978, A2 => n8671, ZN => n7664);
   U949 : OAI211_X1 port map( C1 => n7893, C2 => n8681, A => n7662, B => n7661,
                           ZN => n7663);
   U950 : AOI211_X1 port map( C1 => DATA1(17), C2 => n7832, A => n7664, B => 
                           n7663, ZN => n7716);
   U951 : OAI222_X1 port map( A1 => n7986, A2 => n7716, B1 => n7984, B2 => 
                           n7671, C1 => n7898, C2 => n7665, ZN => n7761);
   U952 : NAND2_X1 port map( A1 => n8403, A2 => n8087, ZN => n7669);
   U953 : NAND4_X1 port map( A1 => n7669, A2 => n7668, A3 => n7667, A4 => n7666
                           , ZN => n7670);
   U954 : AOI21_X1 port map( B1 => n8323, B2 => DATA1(21), A => n7670, ZN => 
                           n7752);
   U955 : OAI222_X1 port map( A1 => n7986, A2 => n7752, B1 => n7984, B2 => 
                           n7716, C1 => n7982, C2 => n7671, ZN => n7783);
   U956 : AOI22_X1 port map( A1 => n7919, A2 => n7761, B1 => n8203, B2 => n7783
                           , ZN => n7672);
   U957 : OAI211_X1 port map( C1 => n7718, C2 => n8330, A => n7673, B => n7672,
                           ZN => n7771);
   U958 : NAND4_X1 port map( A1 => n7677, A2 => n7676, A3 => n7675, A4 => n7674
                           , ZN => n7678);
   U959 : AOI21_X1 port map( B1 => n8762, B2 => DATA1(13), A => n7678, ZN => 
                           n7693);
   U960 : NOR2_X1 port map( A1 => n7680, A2 => n7679, ZN => n7682);
   U961 : OAI22_X1 port map( A1 => n7978, A2 => n8654, B1 => n8602, B2 => n7893
                           , ZN => n7681);
   U962 : NOR4_X1 port map( A1 => n7684, A2 => n7683, A3 => n7682, A4 => n7681,
                           ZN => n7730);
   U963 : NAND2_X1 port map( A1 => n9193, A2 => n7776, ZN => n7685);
   U964 : OAI211_X1 port map( C1 => n8526, C2 => n7893, A => n7686, B => n7685,
                           ZN => n7687);
   U965 : AOI211_X1 port map( C1 => n8763, C2 => DATA1(8), A => n7688, B => 
                           n7687, ZN => n7738);
   U966 : OAI222_X1 port map( A1 => n7986, A2 => n7693, B1 => n7984, B2 => 
                           n7730, C1 => n7898, C2 => n7738, ZN => n7920);
   U967 : AOI22_X1 port map( A1 => DATA1(14), A2 => n8762, B1 => n8763, B2 => 
                           DATA1(11), ZN => n7692);
   U968 : AND4_X1 port map( A1 => n7692, A2 => n7691, A3 => n7690, A4 => n7689,
                           ZN => n7697);
   U969 : OAI222_X1 port map( A1 => n7693, A2 => n7898, B1 => n7695, B2 => 
                           n7224, C1 => n7697, C2 => n8186, ZN => n7739);
   U970 : INV_X1 port map( A => n7739, ZN => n7732);
   U971 : OAI222_X1 port map( A1 => n7730, A2 => n7898, B1 => n7697, B2 => 
                           n7224, C1 => n7693, C2 => n8186, ZN => n7803);
   U972 : INV_X1 port map( A => n7803, ZN => n7731);
   U973 : OAI22_X1 port map( A1 => n7732, A2 => n8330, B1 => n7731, B2 => n8780
                           , ZN => n7700);
   U974 : INV_X1 port map( A => n7694, ZN => n7706);
   U975 : OAI222_X1 port map( A1 => n7697, A2 => n7898, B1 => n7696, B2 => 
                           n7224, C1 => n7695, C2 => n7984, ZN => n7698);
   U976 : INV_X1 port map( A => n7698, ZN => n7733);
   U977 : OAI22_X1 port map( A1 => n8777, A2 => n7706, B1 => n7733, B2 => n8778
                           , ZN => n7699);
   U978 : AOI211_X1 port map( C1 => n8785, C2 => n7920, A => n7700, B => n7699,
                           ZN => n7723);
   U979 : OAI22_X1 port map( A1 => n7733, A2 => n8780, B1 => n7732, B2 => n8331
                           , ZN => n7703);
   U980 : INV_X1 port map( A => n7701, ZN => n7717);
   U981 : OAI22_X1 port map( A1 => n7717, A2 => n8044, B1 => n7706, B2 => n8330
                           , ZN => n7702);
   U982 : AOI211_X1 port map( C1 => n8231, C2 => n7746, A => n7703, B => n7702,
                           ZN => n7742);
   U983 : OAI22_X1 port map( A1 => n8793, A2 => n7723, B1 => n7742, B2 => n8788
                           , ZN => n7710);
   U984 : OAI22_X1 port map( A1 => n7718, A2 => n8044, B1 => n7733, B2 => n8331
                           , ZN => n7705);
   U985 : OAI22_X1 port map( A1 => n7717, A2 => n8774, B1 => n7706, B2 => n8780
                           , ZN => n7704);
   U986 : AOI211_X1 port map( C1 => n8203, C2 => n7761, A => n7705, B => n7704,
                           ZN => n7773);
   U987 : OAI22_X1 port map( A1 => n7733, A2 => n8330, B1 => n7731, B2 => n8331
                           , ZN => n7708);
   U988 : OAI22_X1 port map( A1 => n8777, A2 => n7717, B1 => n7706, B2 => n8778
                           , ZN => n7707);
   U989 : AOI211_X1 port map( C1 => n8335, C2 => n7739, A => n7708, B => n7707,
                           ZN => n7928);
   U990 : OAI22_X1 port map( A1 => n7773, A2 => n8790, B1 => n7928, B2 => n8477
                           , ZN => n7709);
   U991 : AOI211_X1 port map( C1 => n8522, C2 => n7771, A => n7710, B => n7709,
                           ZN => n7760);
   U992 : INV_X1 port map( A => n7742, ZN => n7756);
   U993 : AOI21_X1 port map( B1 => n8762, B2 => DATA1(22), A => n7711, ZN => 
                           n7715);
   U994 : AND4_X1 port map( A1 => n7715, A2 => n7714, A3 => n7713, A4 => n7712,
                           ZN => n7767);
   U995 : OAI222_X1 port map( A1 => n7716, A2 => n7898, B1 => n7767, B2 => 
                           n7224, C1 => n7752, C2 => n8186, ZN => n7819);
   U996 : INV_X1 port map( A => n7819, ZN => n7768);
   U997 : OAI22_X1 port map( A1 => n8777, A2 => n7768, B1 => n7717, B2 => n8331
                           , ZN => n7720);
   U998 : INV_X1 port map( A => n7761, ZN => n7755);
   U999 : OAI22_X1 port map( A1 => n7755, A2 => n8774, B1 => n7718, B2 => n8780
                           , ZN => n7719);
   U1000 : AOI211_X1 port map( C1 => n7919, C2 => n7783, A => n7720, B => n7719
                           , ZN => n7824);
   U1001 : OAI22_X1 port map( A1 => n8793, A2 => n7928, B1 => n7824, B2 => 
                           n8786, ZN => n7722);
   U1002 : INV_X1 port map( A => n7771, ZN => n7790);
   U1003 : OAI22_X1 port map( A1 => n7790, A2 => n8790, B1 => n7773, B2 => 
                           n8788, ZN => n7721);
   U1004 : AOI211_X1 port map( C1 => n8100, C2 => n7756, A => n7722, B => n7721
                           , ZN => n7794);
   U1005 : INV_X1 port map( A => n7723, ZN => n7923);
   U1006 : AND3_X1 port map( A1 => n7726, A2 => n7725, A3 => n7724, ZN => n7728
                           );
   U1007 : OAI211_X1 port map( C1 => n7978, C2 => n8634, A => n7728, B => n7727
                           , ZN => n7729);
   U1008 : INV_X1 port map( A => n7729, ZN => n7801);
   U1009 : OAI222_X1 port map( A1 => n7801, A2 => n7898, B1 => n7730, B2 => 
                           n7224, C1 => n7738, C2 => n8186, ZN => n7935);
   U1010 : INV_X1 port map( A => n7935, ZN => n7799);
   U1011 : OAI22_X1 port map( A1 => n7731, A2 => n8330, B1 => n7799, B2 => 
                           n8331, ZN => n7735);
   U1012 : OAI22_X1 port map( A1 => n8777, A2 => n7733, B1 => n7732, B2 => 
                           n8778, ZN => n7734);
   U1013 : AOI211_X1 port map( C1 => n8335, C2 => n7920, A => n7735, B => n7734
                           , ZN => n7963);
   U1014 : OAI22_X1 port map( A1 => n8793, A2 => n7963, B1 => n7928, B2 => 
                           n8788, ZN => n7737);
   U1015 : OAI22_X1 port map( A1 => n7773, A2 => n8786, B1 => n7742, B2 => 
                           n8790, ZN => n7736);
   U1016 : AOI211_X1 port map( C1 => n8797, C2 => n7923, A => n7737, B => n7736
                           , ZN => n7809);
   U1017 : OAI222_X1 port map( A1 => n8803, A2 => n7760, B1 => n7862, B2 => 
                           n7794, C1 => n7809, C2 => n8798, ZN => n7970);
   U1018 : INV_X1 port map( A => n7970, ZN => n7797);
   U1019 : OAI222_X1 port map( A1 => n7986, A2 => n7738, B1 => n7984, B2 => 
                           n7801, C1 => n7898, C2 => n7800, ZN => n7798);
   U1020 : AOI22_X1 port map( A1 => n8272, A2 => n7920, B1 => n8785, B2 => 
                           n7798, ZN => n7741);
   U1021 : AOI22_X1 port map( A1 => n8230, A2 => n7803, B1 => n8203, B2 => 
                           n7739, ZN => n7740);
   U1022 : OAI211_X1 port map( C1 => n7799, C2 => n8780, A => n7741, B => n7740
                           , ZN => n7959);
   U1023 : AOI22_X1 port map( A1 => n8496, A2 => n7923, B1 => n7995, B2 => 
                           n7959, ZN => n7745);
   U1024 : OAI22_X1 port map( A1 => n8790, A2 => n7928, B1 => n8786, B2 => 
                           n7742, ZN => n7743);
   U1025 : INV_X1 port map( A => n7743, ZN => n7744);
   U1026 : OAI211_X1 port map( C1 => n7963, C2 => n8477, A => n7745, B => n7744
                           , ZN => n7929);
   U1027 : INV_X1 port map( A => n7929, ZN => n7810);
   U1028 : OAI222_X1 port map( A1 => n7810, A2 => n8798, B1 => n7809, B2 => 
                           n8803, C1 => n7760, C2 => n8801, ZN => n7968);
   U1029 : AOI22_X1 port map( A1 => n8785, A2 => n7746, B1 => n8230, B2 => 
                           n7819, ZN => n7754);
   U1030 : NAND2_X1 port map( A1 => n8365, A2 => n8087, ZN => n7750);
   U1031 : NAND4_X1 port map( A1 => n7750, A2 => n7749, A3 => n7748, A4 => 
                           n7747, ZN => n7751);
   U1032 : AOI21_X1 port map( B1 => n8323, B2 => DATA1(23), A => n7751, ZN => 
                           n7782);
   U1033 : OAI222_X1 port map( A1 => n7986, A2 => n7782, B1 => n7984, B2 => 
                           n7767, C1 => n7982, C2 => n7752, ZN => n7835);
   U1034 : AOI22_X1 port map( A1 => n8272, A2 => n7783, B1 => n8203, B2 => 
                           n7835, ZN => n7753);
   U1035 : OAI211_X1 port map( C1 => n7755, C2 => n8780, A => n7754, B => n7753
                           , ZN => n7838);
   U1036 : AOI22_X1 port map( A1 => n8522, A2 => n7838, B1 => n7995, B2 => 
                           n7756, ZN => n7758);
   U1037 : INV_X1 port map( A => n7824, ZN => n7786);
   U1038 : AOI22_X1 port map( A1 => n8496, A2 => n7771, B1 => n8524, B2 => 
                           n7786, ZN => n7757);
   U1039 : OAI211_X1 port map( C1 => n7773, C2 => n8477, A => n7758, B => n7757
                           , ZN => n7759);
   U1040 : INV_X1 port map( A => n7759, ZN => n7793);
   U1041 : OAI222_X1 port map( A1 => n7760, A2 => n8798, B1 => n7794, B2 => 
                           n8803, C1 => n7793, C2 => n8801, ZN => n7931);
   U1042 : AOI22_X1 port map( A1 => n8809, A2 => n7968, B1 => n7931, B2 => 
                           n8807, ZN => n7796);
   U1043 : AOI22_X1 port map( A1 => n7835, A2 => n8230, B1 => n7761, B2 => 
                           n8785, ZN => n7762);
   U1044 : INV_X1 port map( A => n7762, ZN => n7770);
   U1045 : AOI22_X1 port map( A1 => DATA1(21), A2 => n8763, B1 => DATA1(20), B2
                           => n7776, ZN => n7766);
   U1046 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(24), ZN => n7763);
   U1047 : AND4_X1 port map( A1 => n7766, A2 => n7765, A3 => n7764, A4 => n7763
                           , ZN => n7818);
   U1048 : OAI222_X1 port map( A1 => n7767, A2 => n7982, B1 => n7818, B2 => 
                           n7224, C1 => n7782, C2 => n8186, ZN => n7834);
   U1049 : INV_X1 port map( A => n7834, ZN => n7853);
   U1050 : OAI22_X1 port map( A1 => n8777, A2 => n7853, B1 => n7768, B2 => 
                           n8330, ZN => n7769);
   U1051 : AOI211_X1 port map( C1 => n8335, C2 => n7783, A => n7770, B => n7769
                           , ZN => n7787);
   U1052 : AOI22_X1 port map( A1 => n8100, A2 => n7771, B1 => n8496, B2 => 
                           n7786, ZN => n7772);
   U1053 : OAI21_X1 port map( B1 => n8793, B2 => n7773, A => n7772, ZN => n7774
                           );
   U1054 : AOI21_X1 port map( B1 => n8524, B2 => n7838, A => n7774, ZN => n7826
                           );
   U1055 : OAI21_X1 port map( B1 => n7787, B2 => n8786, A => n7826, ZN => n7775
                           );
   U1056 : INV_X1 port map( A => n7775, ZN => n7792);
   U1057 : NAND2_X1 port map( A1 => n8286, A2 => n7776, ZN => n7780);
   U1058 : NAND4_X1 port map( A1 => n7780, A2 => n7779, A3 => n7778, A4 => 
                           n7777, ZN => n7781);
   U1059 : AOI21_X1 port map( B1 => n8323, B2 => DATA1(25), A => n7781, ZN => 
                           n7833);
   U1060 : OAI222_X1 port map( A1 => n7986, A2 => n7833, B1 => n7984, B2 => 
                           n7818, C1 => n7982, C2 => n7782, ZN => n7877);
   U1061 : AOI22_X1 port map( A1 => n8335, A2 => n7819, B1 => n8203, B2 => 
                           n7877, ZN => n7785);
   U1062 : AOI22_X1 port map( A1 => n8272, A2 => n7835, B1 => n8785, B2 => 
                           n7783, ZN => n7784);
   U1063 : OAI211_X1 port map( C1 => n7853, C2 => n8044, A => n7785, B => n7784
                           , ZN => n7880);
   U1064 : AOI22_X1 port map( A1 => n8100, A2 => n7786, B1 => n8522, B2 => 
                           n7880, ZN => n7789);
   U1065 : INV_X1 port map( A => n7787, ZN => n7857);
   U1066 : AOI22_X1 port map( A1 => n8496, A2 => n7838, B1 => n8524, B2 => 
                           n7857, ZN => n7788);
   U1067 : OAI211_X1 port map( C1 => n8793, C2 => n7790, A => n7789, B => n7788
                           , ZN => n7791);
   U1068 : INV_X1 port map( A => n7791, ZN => n7841);
   U1069 : OAI222_X1 port map( A1 => n7793, A2 => n8798, B1 => n7792, B2 => 
                           n8803, C1 => n7841, C2 => n8801, ZN => n7886);
   U1070 : OAI222_X1 port map( A1 => n7794, A2 => n8101, B1 => n7793, B2 => 
                           n8803, C1 => n7792, C2 => n8801, ZN => n7864);
   U1071 : AOI22_X1 port map( A1 => n8485, A2 => n7886, B1 => n7864, B2 => 
                           n8811, ZN => n7795);
   U1072 : OAI211_X1 port map( C1 => n8814, C2 => n7797, A => n7796, B => n7795
                           , ZN => n7974);
   U1073 : INV_X1 port map( A => n7974, ZN => n7950);
   U1074 : INV_X1 port map( A => n7968, ZN => n7930);
   U1075 : INV_X1 port map( A => n7798, ZN => n7958);
   U1076 : OAI22_X1 port map( A1 => n7799, A2 => n8330, B1 => n7958, B2 => 
                           n8780, ZN => n7806);
   U1077 : OAI222_X1 port map( A1 => n7802, A2 => n7898, B1 => n7801, B2 => 
                           n7224, C1 => n7800, C2 => n8186, ZN => n8038);
   U1078 : AOI22_X1 port map( A1 => n8231, A2 => n7803, B1 => n8038, B2 => 
                           n8785, ZN => n7804);
   U1079 : INV_X1 port map( A => n7804, ZN => n7805);
   U1080 : AOI211_X1 port map( C1 => n8230, C2 => n7920, A => n7806, B => n7805
                           , ZN => n7938);
   U1081 : INV_X1 port map( A => n7963, ZN => n7924);
   U1082 : AOI22_X1 port map( A1 => n8496, A2 => n7924, B1 => n8524, B2 => 
                           n7923, ZN => n7807);
   U1083 : OAI21_X1 port map( B1 => n8793, B2 => n7938, A => n7807, ZN => n7808
                           );
   U1084 : AOI21_X1 port map( B1 => n8100, B2 => n7959, A => n7808, ZN => n7927
                           );
   U1085 : OAI222_X1 port map( A1 => n8803, A2 => n7810, B1 => n7862, B2 => 
                           n7809, C1 => n7927, C2 => n8798, ZN => n7965);
   U1086 : AOI22_X1 port map( A1 => n8807, A2 => n7970, B1 => n8809, B2 => 
                           n7965, ZN => n7812);
   U1087 : AOI22_X1 port map( A1 => n8811, A2 => n7931, B1 => n8805, B2 => 
                           n7864, ZN => n7811);
   U1088 : OAI211_X1 port map( C1 => n7930, C2 => n8814, A => n7812, B => n7811
                           , ZN => n8059);
   U1089 : NOR2_X1 port map( A1 => n7978, A2 => n8618, ZN => n7817);
   U1090 : NAND3_X1 port map( A1 => n7815, A2 => n7814, A3 => n7813, ZN => 
                           n7816);
   U1091 : AOI211_X1 port map( C1 => n7832, C2 => DATA1(23), A => n7817, B => 
                           n7816, ZN => n7852);
   U1092 : OAI222_X1 port map( A1 => n7986, A2 => n7852, B1 => n7984, B2 => 
                           n7833, C1 => n7982, C2 => n7818, ZN => n7900);
   U1093 : AOI22_X1 port map( A1 => n8785, A2 => n7819, B1 => n8203, B2 => 
                           n7900, ZN => n7821);
   U1094 : AOI22_X1 port map( A1 => n7919, A2 => n7877, B1 => n8335, B2 => 
                           n7835, ZN => n7820);
   U1095 : OAI211_X1 port map( C1 => n7853, C2 => n8330, A => n7821, B => n7820
                           , ZN => n7904);
   U1096 : AOI22_X1 port map( A1 => n8797, A2 => n7838, B1 => n8522, B2 => 
                           n7904, ZN => n7823);
   U1097 : AOI22_X1 port map( A1 => n8496, A2 => n7857, B1 => n8524, B2 => 
                           n7880, ZN => n7822);
   U1098 : OAI211_X1 port map( C1 => n8793, C2 => n7824, A => n7823, B => n7822
                           , ZN => n7825);
   U1099 : INV_X1 port map( A => n7825, ZN => n7861);
   U1100 : OAI222_X1 port map( A1 => n7826, A2 => n8101, B1 => n7841, B2 => 
                           n8803, C1 => n7861, C2 => n8801, ZN => n7885);
   U1101 : INV_X1 port map( A => n7885, ZN => n7909);
   U1102 : AOI22_X1 port map( A1 => n8500, A2 => n7864, B1 => n8809, B2 => 
                           n7931, ZN => n7843);
   U1103 : AOI22_X1 port map( A1 => n8100, A2 => n7857, B1 => n8524, B2 => 
                           n7904, ZN => n7840);
   U1104 : INV_X1 port map( A => n7900, ZN => n7846);
   U1105 : INV_X1 port map( A => DATA1(23), ZN => n8233);
   U1106 : NOR2_X1 port map( A1 => n7978, A2 => n8233, ZN => n7831);
   U1107 : NAND3_X1 port map( A1 => n7829, A2 => n7828, A3 => n7827, ZN => 
                           n7830);
   U1108 : AOI211_X1 port map( C1 => n7832, C2 => n8692, A => n7831, B => n7830
                           , ZN => n7876);
   U1109 : OAI222_X1 port map( A1 => n7986, A2 => n7876, B1 => n7984, B2 => 
                           n7852, C1 => n7898, C2 => n7833, ZN => n7990);
   U1110 : AOI22_X1 port map( A1 => n8272, A2 => n7877, B1 => n8203, B2 => 
                           n7990, ZN => n7837);
   U1111 : AOI22_X1 port map( A1 => n8785, A2 => n7835, B1 => n8335, B2 => 
                           n7834, ZN => n7836);
   U1112 : OAI211_X1 port map( C1 => n7846, C2 => n8778, A => n7837, B => n7836
                           , ZN => n7994);
   U1113 : AOI22_X1 port map( A1 => n8522, A2 => n7994, B1 => n8339, B2 => 
                           n7838, ZN => n7839);
   U1114 : NAND2_X1 port map( A1 => n7840, A2 => n7839, ZN => n7883);
   U1115 : AOI21_X1 port map( B1 => n8496, B2 => n7880, A => n7883, ZN => n7863
                           );
   U1116 : OAI222_X1 port map( A1 => n8803, A2 => n7861, B1 => n7862, B2 => 
                           n7863, C1 => n7841, C2 => n8798, ZN => n8009);
   U1117 : AOI22_X1 port map( A1 => n8807, A2 => n7886, B1 => n8805, B2 => 
                           n8009, ZN => n7842);
   U1118 : OAI211_X1 port map( C1 => n7909, C2 => n8461, A => n7843, B => n7842
                           , ZN => n7954);
   U1119 : AOI22_X1 port map( A1 => n8111, A2 => n8059, B1 => n8351, B2 => 
                           n7954, ZN => n7868);
   U1120 : AOI22_X1 port map( A1 => n8103, A2 => n7864, B1 => n8809, B2 => 
                           n7970, ZN => n7845);
   U1121 : AOI22_X1 port map( A1 => n8811, A2 => n7886, B1 => n8500, B2 => 
                           n7931, ZN => n7844);
   U1122 : OAI211_X1 port map( C1 => n8463, C2 => n7909, A => n7845, B => n7844
                           , ZN => n7914);
   U1123 : INV_X1 port map( A => n7904, ZN => n7856);
   U1124 : INV_X1 port map( A => n7990, ZN => n7903);
   U1125 : OAI22_X1 port map( A1 => n7846, A2 => n8774, B1 => n7903, B2 => 
                           n8778, ZN => n7855);
   U1126 : NAND2_X1 port map( A1 => n8763, A2 => DATA1(25), ZN => n7849);
   U1127 : NAND4_X1 port map( A1 => n7850, A2 => n7849, A3 => n7848, A4 => 
                           n7847, ZN => n7851);
   U1128 : AOI21_X1 port map( B1 => n8323, B2 => DATA1(28), A => n7851, ZN => 
                           n7897);
   U1129 : OAI222_X1 port map( A1 => n7852, A2 => n7982, B1 => n7897, B2 => 
                           n7224, C1 => n7876, C2 => n8186, ZN => n7899);
   U1130 : INV_X1 port map( A => n7899, ZN => n7993);
   U1131 : OAI22_X1 port map( A1 => n8777, A2 => n7993, B1 => n7853, B2 => 
                           n8331, ZN => n7854);
   U1132 : AOI211_X1 port map( C1 => n8335, C2 => n7877, A => n7855, B => n7854
                           , ZN => n7999);
   U1133 : OAI22_X1 port map( A1 => n7856, A2 => n8788, B1 => n7999, B2 => 
                           n8786, ZN => n7860);
   U1134 : AOI22_X1 port map( A1 => n8339, A2 => n7857, B1 => n7994, B2 => 
                           n8524, ZN => n7858);
   U1135 : INV_X1 port map( A => n7858, ZN => n7859);
   U1136 : AOI211_X1 port map( C1 => n8100, C2 => n7880, A => n7860, B => n7859
                           , ZN => n7870);
   U1137 : OAI222_X1 port map( A1 => n8803, A2 => n7863, B1 => n7862, B2 => 
                           n7870, C1 => n7861, C2 => n8798, ZN => n7912);
   U1138 : AOI22_X1 port map( A1 => n8811, A2 => n8009, B1 => n8805, B2 => 
                           n7912, ZN => n7866);
   U1139 : AOI22_X1 port map( A1 => n8500, A2 => n7886, B1 => n8809, B2 => 
                           n7864, ZN => n7865);
   U1140 : OAI211_X1 port map( C1 => n7909, C2 => n8383, A => n7866, B => n7865
                           , ZN => n7913);
   U1141 : AOI22_X1 port map( A1 => n8239, A2 => n7914, B1 => n8828, B2 => 
                           n7913, ZN => n7867);
   U1142 : OAI211_X1 port map( C1 => n7950, C2 => n8823, A => n7868, B => n7867
                           , ZN => n7869);
   U1143 : INV_X1 port map( A => n7869, ZN => n8022);
   U1144 : INV_X1 port map( A => n7912, ZN => n8006);
   U1145 : INV_X1 port map( A => n7870, ZN => n7907);
   U1146 : NAND4_X1 port map( A1 => n7874, A2 => n7873, A3 => n7872, A4 => 
                           n7871, ZN => n7875);
   U1147 : AOI21_X1 port map( B1 => n8762, B2 => DATA1(29), A => n7875, ZN => 
                           n7981);
   U1148 : OAI222_X1 port map( A1 => n7986, A2 => n7981, B1 => n7984, B2 => 
                           n7897, C1 => n7982, C2 => n7876, ZN => n7988);
   U1149 : AOI22_X1 port map( A1 => n8229, A2 => n7990, B1 => n8203, B2 => 
                           n7988, ZN => n7879);
   U1150 : AOI22_X1 port map( A1 => n8785, A2 => n7877, B1 => n8335, B2 => 
                           n7900, ZN => n7878);
   U1151 : OAI211_X1 port map( C1 => n7993, C2 => n8044, A => n7879, B => n7878
                           , ZN => n7976);
   U1152 : AOI22_X1 port map( A1 => n8496, A2 => n7994, B1 => n8522, B2 => 
                           n7976, ZN => n7882);
   U1153 : AOI22_X1 port map( A1 => n8100, A2 => n7904, B1 => n7995, B2 => 
                           n7880, ZN => n7881);
   U1154 : OAI211_X1 port map( C1 => n7999, C2 => n8790, A => n7882, B => n7881
                           , ZN => n8002);
   U1155 : AOI222_X1 port map( A1 => n7883, A2 => n8051, B1 => n7907, B2 => 
                           n8431, C1 => n8002, C2 => n8456, ZN => n8003);
   U1156 : INV_X1 port map( A => n8009, ZN => n7908);
   U1157 : OAI22_X1 port map( A1 => n8463, A2 => n8003, B1 => n7908, B2 => 
                           n8383, ZN => n7884);
   U1158 : INV_X1 port map( A => n7884, ZN => n7888);
   U1159 : AOI22_X1 port map( A1 => n8809, A2 => n7886, B1 => n7885, B2 => 
                           n8500, ZN => n7887);
   U1160 : OAI211_X1 port map( C1 => n8461, C2 => n8006, A => n7888, B => n7887
                           , ZN => n8016);
   U1161 : INV_X1 port map( A => n7954, ZN => n8010);
   U1162 : OAI22_X1 port map( A1 => n8819, A2 => n7950, B1 => n8817, B2 => 
                           n8010, ZN => n7890);
   U1163 : INV_X1 port map( A => n7914, ZN => n7951);
   U1164 : INV_X1 port map( A => n7913, ZN => n8012);
   U1165 : OAI22_X1 port map( A1 => n8823, A2 => n7951, B1 => n8821, B2 => 
                           n8012, ZN => n7889);
   U1166 : AOI211_X1 port map( C1 => n8828, C2 => n8016, A => n7890, B => n7889
                           , ZN => n8017);
   U1167 : OAI211_X1 port map( C1 => n7893, C2 => n8577, A => n7892, B => n7891
                           , ZN => n7894);
   U1168 : AOI211_X1 port map( C1 => DATA1(29), C2 => n7896, A => n7895, B => 
                           n7894, ZN => n7983);
   U1169 : OAI222_X1 port map( A1 => n7986, A2 => n7983, B1 => n7984, B2 => 
                           n7981, C1 => n7898, C2 => n7897, ZN => n7989);
   U1170 : AOI22_X1 port map( A1 => n8229, A2 => n7899, B1 => n8231, B2 => 
                           n7989, ZN => n7902);
   U1171 : AOI22_X1 port map( A1 => n8785, A2 => n7900, B1 => n8230, B2 => 
                           n7988, ZN => n7901);
   U1172 : OAI211_X1 port map( C1 => n7903, C2 => n8780, A => n7902, B => n7901
                           , ZN => n7975);
   U1173 : AOI22_X1 port map( A1 => n8797, A2 => n7994, B1 => n8522, B2 => 
                           n7975, ZN => n7906);
   U1174 : AOI22_X1 port map( A1 => n8524, A2 => n7976, B1 => n7995, B2 => 
                           n7904, ZN => n7905);
   U1175 : OAI211_X1 port map( C1 => n7999, C2 => n8788, A => n7906, B => n7905
                           , ZN => n8001);
   U1176 : AOI222_X1 port map( A1 => n7907, A2 => n8051, B1 => n8002, B2 => 
                           n8431, C1 => n8001, C2 => n8456, ZN => n8005);
   U1177 : OAI22_X1 port map( A1 => n8463, A2 => n8005, B1 => n7908, B2 => 
                           n8814, ZN => n7911);
   U1178 : OAI22_X1 port map( A1 => n8052, A2 => n7909, B1 => n8003, B2 => 
                           n8461, ZN => n7910);
   U1179 : AOI211_X1 port map( C1 => n8807, C2 => n7912, A => n7911, B => n7910
                           , ZN => n8013);
   U1180 : AOI22_X1 port map( A1 => n8109, A2 => n7954, B1 => n8351, B2 => 
                           n8016, ZN => n7916);
   U1181 : AOI22_X1 port map( A1 => n8111, A2 => n7914, B1 => n8239, B2 => 
                           n7913, ZN => n7915);
   U1182 : OAI211_X1 port map( C1 => n8553, C2 => n8013, A => n7916, B => n7915
                           , ZN => n7917);
   U1183 : INV_X1 port map( A => n7917, ZN => n8019);
   U1184 : OAI222_X1 port map( A1 => n8060, A2 => n8022, B1 => n8017, B2 => 
                           n8834, C1 => n8019, C2 => n8832, ZN => n7918);
   U1185 : INV_X1 port map( A => n7918, ZN => n8065);
   U1186 : AOI22_X1 port map( A1 => n7919, A2 => n7935, B1 => n8335, B2 => 
                           n8038, ZN => n7922);
   U1187 : AOI22_X1 port map( A1 => n8785, A2 => n7955, B1 => n8231, B2 => 
                           n7920, ZN => n7921);
   U1188 : OAI211_X1 port map( C1 => n7958, C2 => n8330, A => n7922, B => n7921
                           , ZN => n8047);
   U1189 : AOI22_X1 port map( A1 => n8496, A2 => n7959, B1 => n7995, B2 => 
                           n8047, ZN => n7926);
   U1190 : AOI22_X1 port map( A1 => n8524, A2 => n7924, B1 => n8522, B2 => 
                           n7923, ZN => n7925);
   U1191 : OAI211_X1 port map( C1 => n7938, C2 => n8477, A => n7926, B => n7925
                           , ZN => n7964);
   U1192 : OAI21_X1 port map( B1 => n7928, B2 => n8786, A => n7927, ZN => n7942
                           );
   U1193 : AOI222_X1 port map( A1 => n7964, A2 => n8051, B1 => n7942, B2 => 
                           n7943, C1 => n7929, C2 => n8456, ZN => n8364);
   U1194 : OAI22_X1 port map( A1 => n8052, A2 => n8364, B1 => n7930, B2 => 
                           n8383, ZN => n7934);
   U1195 : AOI22_X1 port map( A1 => n8485, A2 => n7931, B1 => n7970, B2 => 
                           n8811, ZN => n7932);
   U1196 : INV_X1 port map( A => n7932, ZN => n7933);
   U1197 : AOI211_X1 port map( C1 => n8500, C2 => n7965, A => n7934, B => n7933
                           , ZN => n8236);
   U1198 : AOI22_X1 port map( A1 => n8229, A2 => n8038, B1 => n8231, B2 => 
                           n7935, ZN => n7937);
   U1199 : AOI22_X1 port map( A1 => n8785, A2 => n8041, B1 => n8335, B2 => 
                           n7955, ZN => n7936);
   U1200 : OAI211_X1 port map( C1 => n7958, C2 => n8044, A => n7937, B => n7936
                           , ZN => n8495);
   U1201 : INV_X1 port map( A => n8047, ZN => n8476);
   U1202 : INV_X1 port map( A => n7938, ZN => n8046);
   U1203 : AOI22_X1 port map( A1 => n8496, A2 => n8046, B1 => n8524, B2 => 
                           n7959, ZN => n7939);
   U1204 : OAI21_X1 port map( B1 => n8476, B2 => n8477, A => n7939, ZN => n7940
                           );
   U1205 : AOI21_X1 port map( B1 => n8339, B2 => n8495, A => n7940, ZN => n7962
                           );
   U1206 : INV_X1 port map( A => n7962, ZN => n7941);
   U1207 : AOI222_X1 port map( A1 => n7943, A2 => n7964, B1 => n8456, B2 => 
                           n7942, C1 => n7941, C2 => n8051, ZN => n8382);
   U1208 : AOI22_X1 port map( A1 => n8811, A2 => n7968, B1 => n8807, B2 => 
                           n7965, ZN => n7944);
   U1209 : OAI21_X1 port map( B1 => n8364, B2 => n8814, A => n7944, ZN => n7945
                           );
   U1210 : INV_X1 port map( A => n7945, ZN => n7946);
   U1211 : OAI21_X1 port map( B1 => n8052, B2 => n8382, A => n7946, ZN => n7969
                           );
   U1212 : INV_X1 port map( A => n7969, ZN => n7947);
   U1213 : OAI22_X1 port map( A1 => n8236, A2 => n8823, B1 => n7947, B2 => 
                           n8819, ZN => n7949);
   U1214 : OAI22_X1 port map( A1 => n8553, A2 => n7951, B1 => n7950, B2 => 
                           n8821, ZN => n7948);
   U1215 : AOI211_X1 port map( C1 => n8239, C2 => n8059, A => n7949, B => n7948
                           , ZN => n8061);
   U1216 : OAI22_X1 port map( A1 => n7950, A2 => n8817, B1 => n8236, B2 => 
                           n8819, ZN => n7953);
   U1217 : INV_X1 port map( A => n8059, ZN => n7971);
   U1218 : OAI22_X1 port map( A1 => n7951, A2 => n8821, B1 => n7971, B2 => 
                           n8823, ZN => n7952);
   U1219 : AOI211_X1 port map( C1 => n8828, C2 => n7954, A => n7953, B => n7952
                           , ZN => n8023);
   U1220 : INV_X1 port map( A => n8495, ZN => n8475);
   U1221 : AOI22_X1 port map( A1 => n8229, A2 => n7955, B1 => n8230, B2 => 
                           n8038, ZN => n7957);
   U1222 : AOI22_X1 port map( A1 => n8785, A2 => n8040, B1 => n8335, B2 => 
                           n8041, ZN => n7956);
   U1223 : OAI211_X1 port map( C1 => n8777, C2 => n7958, A => n7957, B => n7956
                           , ZN => n8521);
   U1224 : AOI22_X1 port map( A1 => n8496, A2 => n8047, B1 => n8339, B2 => 
                           n8521, ZN => n7961);
   U1225 : AOI22_X1 port map( A1 => n8524, A2 => n8046, B1 => n8522, B2 => 
                           n7959, ZN => n7960);
   U1226 : OAI211_X1 port map( C1 => n8475, C2 => n8477, A => n7961, B => n7960
                           , ZN => n8432);
   U1227 : OAI21_X1 port map( B1 => n7963, B2 => n8786, A => n7962, ZN => n8050
                           );
   U1228 : AOI222_X1 port map( A1 => n8432, A2 => n8051, B1 => n8050, B2 => 
                           n8431, C1 => n7964, C2 => n8456, ZN => n8402);
   U1229 : OAI22_X1 port map( A1 => n8052, A2 => n8402, B1 => n8364, B2 => 
                           n8383, ZN => n7967);
   U1230 : INV_X1 port map( A => n7965, ZN => n8053);
   U1231 : OAI22_X1 port map( A1 => n8053, A2 => n8461, B1 => n8382, B2 => 
                           n8814, ZN => n7966);
   U1232 : AOI211_X1 port map( C1 => n8485, C2 => n7968, A => n7967, B => n7966
                           , ZN => n8285);
   U1233 : OAI22_X1 port map( A1 => n8236, A2 => n8817, B1 => n8285, B2 => 
                           n8819, ZN => n7973);
   U1234 : AOI21_X1 port map( B1 => n8485, B2 => n7970, A => n7969, ZN => n8263
                           );
   U1235 : OAI22_X1 port map( A1 => n7971, A2 => n8821, B1 => n8263, B2 => 
                           n8823, ZN => n7972);
   U1236 : AOI211_X1 port map( C1 => n8828, C2 => n7974, A => n7973, B => n7972
                           , ZN => n8208);
   U1237 : OAI222_X1 port map( A1 => n8834, A2 => n8061, B1 => n8832, B2 => 
                           n8023, C1 => n8208, C2 => n8060, ZN => n8168);
   U1238 : OAI222_X1 port map( A1 => n8834, A2 => n8022, B1 => n8832, B2 => 
                           n8017, C1 => n8023, C2 => n8060, ZN => n8137);
   U1239 : AOI22_X1 port map( A1 => n8842, A2 => n8168, B1 => n8836, B2 => 
                           n8137, ZN => n8026);
   U1240 : AOI22_X1 port map( A1 => n8496, A2 => n7976, B1 => n8524, B2 => 
                           n7975, ZN => n7998);
   U1241 : INV_X1 port map( A => DATA1(27), ZN => n8171);
   U1242 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(30), ZN => n8129);
   U1243 : OAI211_X1 port map( C1 => n7978, C2 => n8171, A => n8129, B => n7977
                           , ZN => n7979);
   U1244 : AOI211_X1 port map( C1 => n8323, C2 => DATA1(31), A => n7980, B => 
                           n7979, ZN => n7985);
   U1245 : OAI222_X1 port map( A1 => n7986, A2 => n7985, B1 => n7984, B2 => 
                           n7983, C1 => n7982, C2 => n7981, ZN => n7987);
   U1246 : AOI22_X1 port map( A1 => n8229, A2 => n7988, B1 => n8231, B2 => 
                           n7987, ZN => n7992);
   U1247 : AOI22_X1 port map( A1 => n8785, A2 => n7990, B1 => n8230, B2 => 
                           n7989, ZN => n7991);
   U1248 : OAI211_X1 port map( C1 => n7993, C2 => n8780, A => n7992, B => n7991
                           , ZN => n7996);
   U1249 : AOI22_X1 port map( A1 => n8522, A2 => n7996, B1 => n7995, B2 => 
                           n7994, ZN => n7997);
   U1250 : OAI211_X1 port map( C1 => n7999, C2 => n8477, A => n7998, B => n7997
                           , ZN => n8000);
   U1251 : AOI222_X1 port map( A1 => n8002, A2 => n8051, B1 => n8001, B2 => 
                           n8431, C1 => n8000, C2 => n8456, ZN => n8004);
   U1252 : OAI22_X1 port map( A1 => n8463, A2 => n8004, B1 => n8003, B2 => 
                           n8383, ZN => n8008);
   U1253 : OAI22_X1 port map( A1 => n8006, A2 => n8814, B1 => n8005, B2 => 
                           n8461, ZN => n8007);
   U1254 : AOI211_X1 port map( C1 => n8809, C2 => n8009, A => n8008, B => n8007
                           , ZN => n8011);
   U1255 : OAI22_X1 port map( A1 => n8553, A2 => n8011, B1 => n8010, B2 => 
                           n8819, ZN => n8015);
   U1256 : OAI22_X1 port map( A1 => n8013, A2 => n8821, B1 => n8012, B2 => 
                           n8823, ZN => n8014);
   U1257 : AOI211_X1 port map( C1 => n8239, C2 => n8016, A => n8015, B => n8014
                           , ZN => n8018);
   U1258 : OAI222_X1 port map( A1 => n8834, A2 => n8019, B1 => n8832, B2 => 
                           n8018, C1 => n8017, C2 => n8060, ZN => n8024);
   U1259 : NOR2_X1 port map( A1 => n8021, A2 => n8020, ZN => n8840);
   U1260 : OAI222_X1 port map( A1 => n8834, A2 => n8023, B1 => n8832, B2 => 
                           n8022, C1 => n8061, C2 => n8829, ZN => n8146);
   U1261 : AOI22_X1 port map( A1 => n8838, A2 => n8024, B1 => n8840, B2 => 
                           n8146, ZN => n8025);
   U1262 : OAI211_X1 port map( C1 => n8065, C2 => n8845, A => n8026, B => n8025
                           , ZN => n8035);
   U1263 : INV_X1 port map( A => n8027, ZN => n8028);
   U1264 : NOR3_X1 port map( A1 => DATA1(31), A2 => DATA2_I_31_port, A3 => 
                           n8028, ZN => n8034);
   U1265 : AOI22_X1 port map( A1 => n8530, A2 => dataout_mul_31_port, B1 => 
                           DATA2_I_31_port, B2 => n8029, ZN => n8032);
   U1266 : NOR2_X1 port map( A1 => DATA2(31), A2 => n8128, ZN => n8705);
   U1267 : NAND2_X1 port map( A1 => n8128, A2 => DATA2(31), ZN => n8707);
   U1268 : INV_X1 port map( A => n8707, ZN => n8030);
   U1269 : OAI21_X1 port map( B1 => n8705, B2 => n8030, A => n8567, ZN => n8031
                           );
   U1270 : OAI211_X1 port map( C1 => n8527, C2 => n8859, A => n8032, B => n8031
                           , ZN => n8033);
   U1271 : AOI211_X1 port map( C1 => n8479, C2 => n8035, A => n8034, B => n8033
                           , ZN => n8067);
   U1272 : NAND2_X1 port map( A1 => DATA2(0), A2 => n8842, ZN => n8037);
   U1273 : NOR2_X1 port map( A1 => n8037, A2 => n8036, ZN => n8852);
   U1274 : AOI22_X1 port map( A1 => n8167, A2 => n8137, B1 => n8840, B2 => 
                           n8168, ZN => n8063);
   U1275 : INV_X1 port map( A => n8402, ZN => n8056);
   U1276 : INV_X1 port map( A => n8521, ZN => n8478);
   U1277 : AOI22_X1 port map( A1 => n8785, A2 => n8039, B1 => n8231, B2 => 
                           n8038, ZN => n8043);
   U1278 : AOI22_X1 port map( A1 => n8229, A2 => n8041, B1 => n8335, B2 => 
                           n8040, ZN => n8042);
   U1279 : OAI211_X1 port map( C1 => n8045, C2 => n8044, A => n8043, B => n8042
                           , ZN => n8523);
   U1280 : AOI22_X1 port map( A1 => n8496, A2 => n8495, B1 => n8339, B2 => 
                           n8523, ZN => n8049);
   U1281 : AOI22_X1 port map( A1 => n8524, A2 => n8047, B1 => n8522, B2 => 
                           n8046, ZN => n8048);
   U1282 : OAI211_X1 port map( C1 => n8478, C2 => n8477, A => n8049, B => n8048
                           , ZN => n8455);
   U1283 : AOI222_X1 port map( A1 => n8455, A2 => n8051, B1 => n8432, B2 => 
                           n8431, C1 => n8050, C2 => n8456, ZN => n8422);
   U1284 : OAI22_X1 port map( A1 => n8052, A2 => n8422, B1 => n8382, B2 => 
                           n8383, ZN => n8055);
   U1285 : OAI22_X1 port map( A1 => n8463, A2 => n8053, B1 => n8364, B2 => 
                           n8461, ZN => n8054);
   U1286 : AOI211_X1 port map( C1 => n8500, C2 => n8056, A => n8055, B => n8054
                           , ZN => n8301);
   U1287 : OAI22_X1 port map( A1 => n8263, A2 => n8817, B1 => n8301, B2 => 
                           n8819, ZN => n8058);
   U1288 : OAI22_X1 port map( A1 => n8236, A2 => n8821, B1 => n8285, B2 => 
                           n8823, ZN => n8057);
   U1289 : AOI211_X1 port map( C1 => n8828, C2 => n8059, A => n8058, B => n8057
                           , ZN => n8215);
   U1290 : OAI222_X1 port map( A1 => n8834, A2 => n8208, B1 => n8832, B2 => 
                           n8061, C1 => n8215, C2 => n8060, ZN => n8194);
   U1291 : AOI22_X1 port map( A1 => n8842, A2 => n8194, B1 => n8836, B2 => 
                           n8146, ZN => n8062);
   U1292 : OAI211_X1 port map( C1 => n8065, C2 => n8064, A => n8063, B => n8062
                           , ZN => n8077);
   U1293 : NAND3_X1 port map( A1 => n8852, A2 => n8857, A3 => n8077, ZN => 
                           n8066);
   U1294 : OAI211_X1 port map( C1 => n8068, C2 => n8128, A => n8067, B => n8066
                           , ZN => OUTALU(31));
   U1295 : AOI21_X1 port map( B1 => n8071, B2 => n8070, A => n8069, ZN => n8076
                           );
   U1296 : INV_X1 port map( A => DATA2(30), ZN => n8860);
   U1297 : OAI22_X1 port map( A1 => n8577, A2 => DATA2(30), B1 => n8860, B2 => 
                           DATA1(30), ZN => n8701);
   U1298 : INV_X1 port map( A => n8701, ZN => n8626);
   U1299 : INV_X1 port map( A => n8505, ZN => n8546);
   U1300 : OAI21_X1 port map( B1 => n8546, B2 => n8860, A => n8147, ZN => n8072
                           );
   U1301 : AOI22_X1 port map( A1 => DATA1(30), A2 => n8072, B1 => n8575, B2 => 
                           dataout_mul_30_port, ZN => n8074);
   U1302 : NAND3_X1 port map( A1 => n8153, A2 => n8848, A3 => DATA1(31), ZN => 
                           n8073);
   U1303 : OAI211_X1 port map( C1 => n8626, C2 => n8525, A => n8074, B => n8073
                           , ZN => n8075);
   U1304 : AOI211_X1 port map( C1 => n8479, C2 => n8077, A => n8076, B => n8075
                           , ZN => n8078);
   U1305 : OAI21_X1 port map( B1 => n8080, B2 => n8079, A => n8078, ZN => 
                           OUTALU(30));
   U1306 : INV_X1 port map( A => n8125, ZN => n8127);
   U1307 : OAI22_X1 port map( A1 => n8568, A2 => n8083, B1 => n8317, B2 => 
                           n8082, ZN => n8081);
   U1308 : INV_X1 port map( A => n8081, ZN => n8126);
   U1309 : AOI22_X1 port map( A1 => n8084, A2 => n8083, B1 => n8572, B2 => 
                           n8082, ZN => n8124);
   U1310 : INV_X1 port map( A => DATA1(0), ZN => n8635);
   U1311 : NAND2_X1 port map( A1 => n8323, A2 => DATA1(2), ZN => n8085);
   U1312 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(1), ZN => n8765);
   U1313 : OAI211_X1 port map( C1 => n8130, C2 => n8635, A => n8085, B => n8765
                           , ZN => n8122);
   U1314 : AOI22_X1 port map( A1 => n8167, A2 => n8839, B1 => n8836, B2 => 
                           n8841, ZN => n8117);
   U1315 : INV_X1 port map( A => n8086, ZN => n8338);
   U1316 : AOI22_X1 port map( A1 => DATA1(2), A2 => n8323, B1 => n9192, B2 => 
                           n8087, ZN => n8091);
   U1317 : NAND4_X1 port map( A1 => n8091, A2 => n8090, A3 => n8089, A4 => 
                           n8088, ZN => n8773);
   U1318 : AOI222_X1 port map( A1 => n8092, A2 => n8772, B1 => n8773, B2 => 
                           n8770, C1 => n8329, C2 => n8768, ZN => n8775);
   U1319 : OAI22_X1 port map( A1 => n8777, A2 => n8775, B1 => n8332, B2 => 
                           n8780, ZN => n8095);
   U1320 : OAI22_X1 port map( A1 => n8093, A2 => n8774, B1 => n8781, B2 => 
                           n8778, ZN => n8094);
   U1321 : AOI211_X1 port map( C1 => n8785, C2 => n8096, A => n8095, B => n8094
                           , ZN => n8789);
   U1322 : OAI22_X1 port map( A1 => n8792, A2 => n8788, B1 => n8789, B2 => 
                           n8786, ZN => n8099);
   U1323 : OAI22_X1 port map( A1 => n8793, A2 => n8097, B1 => n8761, B2 => 
                           n8790, ZN => n8098);
   U1324 : AOI211_X1 port map( C1 => n8100, C2 => n8338, A => n8099, B => n8098
                           , ZN => n8799);
   U1325 : OAI222_X1 port map( A1 => n8803, A2 => n8340, B1 => n8801, B2 => 
                           n8799, C1 => n8102, C2 => n8101, ZN => n8806);
   U1326 : AOI22_X1 port map( A1 => n8103, A2 => n8808, B1 => n8805, B2 => 
                           n8806, ZN => n8106);
   U1327 : AOI22_X1 port map( A1 => n8500, A2 => n8342, B1 => n8809, B2 => 
                           n8104, ZN => n8105);
   U1328 : OAI211_X1 port map( C1 => n8815, C2 => n8461, A => n8106, B => n8105
                           , ZN => n8816);
   U1329 : AOI22_X1 port map( A1 => n8239, A2 => n8107, B1 => n8828, B2 => 
                           n8816, ZN => n8113);
   U1330 : AOI22_X1 port map( A1 => n8111, A2 => n8110, B1 => n8109, B2 => 
                           n8108, ZN => n8112);
   U1331 : OAI211_X1 port map( C1 => n8824, C2 => n8821, A => n8113, B => n8112
                           , ZN => n8114);
   U1332 : INV_X1 port map( A => n8114, ZN => n8830);
   U1333 : OAI222_X1 port map( A1 => n8834, A2 => n8352, B1 => n8829, B2 => 
                           n8115, C1 => n8830, C2 => n8832, ZN => n8835);
   U1334 : AOI22_X1 port map( A1 => n8838, A2 => n8835, B1 => n8840, B2 => 
                           n8353, ZN => n8116);
   U1335 : AOI21_X1 port map( B1 => n8117, B2 => n8116, A => n8536, ZN => n8121
                           );
   U1336 : AOI22_X1 port map( A1 => DATA2(2), A2 => n8585, B1 => DATA1(2), B2 
                           => n8890, ZN => n8742);
   U1337 : NOR3_X1 port map( A1 => n8546, A2 => n8585, A3 => n8890, ZN => n8118
                           );
   U1338 : AOI21_X1 port map( B1 => dataout_mul_2_port, B2 => n8530, A => n8118
                           , ZN => n8119);
   U1339 : OAI21_X1 port map( B1 => n8742, B2 => n8525, A => n8119, ZN => n8120
                           );
   U1340 : AOI211_X1 port map( C1 => n8479, C2 => n8122, A => n8121, B => n8120
                           , ZN => n8123);
   U1341 : OAI221_X1 port map( B1 => n8127, B2 => n8126, C1 => n8125, C2 => 
                           n8124, A => n8123, ZN => OUTALU(2));
   U1342 : NOR2_X1 port map( A1 => DATA2(29), A2 => n8131, ZN => n8702);
   U1343 : INV_X1 port map( A => DATA2(29), ZN => n8861);
   U1344 : NOR2_X1 port map( A1 => n8861, A2 => DATA1(29), ZN => n8625);
   U1345 : NOR2_X1 port map( A1 => n8702, A2 => n8625, ZN => n8745);
   U1346 : AOI221_X1 port map( B1 => n8130, B2 => n8129, C1 => n8128, C2 => 
                           n8129, A => n8536, ZN => n8133);
   U1347 : AOI221_X1 port map( B1 => n8546, B2 => n8147, C1 => n8861, C2 => 
                           n8147, A => n8131, ZN => n8132);
   U1348 : AOI211_X1 port map( C1 => dataout_mul_29_port, C2 => n8530, A => 
                           n8133, B => n8132, ZN => n8145);
   U1349 : OAI22_X1 port map( A1 => n8202, A2 => n8149, B1 => n8199, B2 => 
                           n8148, ZN => n8142);
   U1350 : INV_X1 port map( A => n8134, ZN => n8135);
   U1351 : AOI21_X1 port map( B1 => n8136, B2 => n8143, A => n8135, ZN => n8141
                           );
   U1352 : AOI22_X1 port map( A1 => n8838, A2 => n8137, B1 => n8836, B2 => 
                           n8168, ZN => n8139);
   U1353 : AOI22_X1 port map( A1 => n8167, A2 => n8146, B1 => n8840, B2 => 
                           n8194, ZN => n8138);
   U1354 : AOI21_X1 port map( B1 => n8139, B2 => n8138, A => n8547, ZN => n8140
                           );
   U1355 : AOI211_X1 port map( C1 => n8143, C2 => n8142, A => n8141, B => n8140
                           , ZN => n8144);
   U1356 : OAI211_X1 port map( C1 => n8745, C2 => n8525, A => n8145, B => n8144
                           , ZN => OUTALU(29));
   U1357 : AOI222_X1 port map( A1 => n8146, A2 => n8838, B1 => n8168, B2 => 
                           n8167, C1 => n8194, C2 => n8836, ZN => n8166);
   U1358 : INV_X1 port map( A => DATA2(28), ZN => n8862);
   U1359 : OAI21_X1 port map( B1 => n8546, B2 => n8862, A => n8147, ZN => n8159
                           );
   U1360 : AOI22_X1 port map( A1 => n8224, A2 => n8149, B1 => n8218, B2 => 
                           n8148, ZN => n8150);
   U1361 : AOI21_X1 port map( B1 => n8151, B2 => n8163, A => n8150, ZN => n8158
                           );
   U1362 : AOI22_X1 port map( A1 => n8152, A2 => DATA1(30), B1 => n8763, B2 => 
                           DATA1(31), ZN => n8156);
   U1363 : NAND2_X1 port map( A1 => n8153, A2 => DATA1(29), ZN => n8155);
   U1364 : AOI22_X1 port map( A1 => DATA1(28), A2 => DATA2(28), B1 => n8862, B2
                           => n8700, ZN => n8717);
   U1365 : AOI22_X1 port map( A1 => dataout_mul_28_port, A2 => n8575, B1 => 
                           n8567, B2 => n8717, ZN => n8154);
   U1366 : OAI221_X1 port map( B1 => n8536, B2 => n8156, C1 => n8536, C2 => 
                           n8155, A => n8154, ZN => n8157);
   U1367 : AOI211_X1 port map( C1 => DATA1(28), C2 => n8159, A => n8158, B => 
                           n8157, ZN => n8165);
   U1368 : NOR2_X1 port map( A1 => n8161, A2 => n8160, ZN => n8179);
   U1369 : AOI22_X1 port map( A1 => n8170, A2 => n8224, B1 => n8169, B2 => 
                           n8218, ZN => n8162);
   U1370 : INV_X1 port map( A => n8162, ZN => n8176);
   U1371 : NAND3_X1 port map( A1 => n8179, A2 => n8163, A3 => n8176, ZN => 
                           n8164);
   U1372 : OAI211_X1 port map( C1 => n8166, C2 => n8547, A => n8165, B => n8164
                           , ZN => OUTALU(28));
   U1373 : AOI22_X1 port map( A1 => n8838, A2 => n8168, B1 => n8167, B2 => 
                           n8194, ZN => n8181);
   U1374 : OAI22_X1 port map( A1 => n8202, A2 => n8170, B1 => n8199, B2 => 
                           n8169, ZN => n8178);
   U1375 : INV_X1 port map( A => n8179, ZN => n8177);
   U1376 : NOR2_X1 port map( A1 => n8171, A2 => DATA2(27), ZN => n8696);
   U1377 : INV_X1 port map( A => n8696, ZN => n8578);
   U1378 : NAND2_X1 port map( A1 => DATA2(27), A2 => n8171, ZN => n8630);
   U1379 : INV_X1 port map( A => DATA2(27), ZN => n8863);
   U1380 : AOI211_X1 port map( C1 => n8527, C2 => n8574, A => n8171, B => n8863
                           , ZN => n8173);
   U1381 : NOR3_X1 port map( A1 => n8187, A2 => n8536, A3 => n7224, ZN => n8172
                           );
   U1382 : AOI211_X1 port map( C1 => n8530, C2 => dataout_mul_27_port, A => 
                           n8173, B => n8172, ZN => n8174);
   U1383 : OAI221_X1 port map( B1 => n8525, B2 => n8578, C1 => n8525, C2 => 
                           n8630, A => n8174, ZN => n8175);
   U1384 : AOI221_X1 port map( B1 => n8179, B2 => n8178, C1 => n8177, C2 => 
                           n8176, A => n8175, ZN => n8180);
   U1385 : OAI21_X1 port map( B1 => n8181, B2 => n8547, A => n8180, ZN => 
                           OUTALU(27));
   U1386 : OAI22_X1 port map( A1 => n8182, A2 => n8202, B1 => n8200, B2 => 
                           n8199, ZN => n8209);
   U1387 : NAND2_X1 port map( A1 => n8183, A2 => n8209, ZN => n8198);
   U1388 : OAI22_X1 port map( A1 => n8185, A2 => n8202, B1 => n8184, B2 => 
                           n8199, ZN => n8193);
   U1389 : INV_X1 port map( A => DATA2(26), ZN => n8864);
   U1390 : INV_X1 port map( A => DATA1(26), ZN => n8579);
   U1391 : AOI22_X1 port map( A1 => DATA1(26), A2 => n8864, B1 => DATA2(26), B2
                           => n8579, ZN => n8695);
   U1392 : OAI22_X1 port map( A1 => n8188, A2 => n7986, B1 => n8187, B2 => 
                           n8186, ZN => n8189);
   U1393 : AOI22_X1 port map( A1 => n8848, A2 => n8189, B1 => n8530, B2 => 
                           dataout_mul_26_port, ZN => n8191);
   U1394 : NAND3_X1 port map( A1 => DATA2(26), A2 => DATA1(26), A3 => n8505, ZN
                           => n8190);
   U1395 : OAI211_X1 port map( C1 => n8695, C2 => n8525, A => n8191, B => n8190
                           , ZN => n8192);
   U1396 : AOI21_X1 port map( B1 => n8197, B2 => n8193, A => n8192, ZN => n8196
                           );
   U1397 : NAND3_X1 port map( A1 => n8479, A2 => n8838, A3 => n8194, ZN => 
                           n8195);
   U1398 : OAI211_X1 port map( C1 => n8198, C2 => n8197, A => n8196, B => n8195
                           , ZN => OUTALU(26));
   U1399 : OR2_X1 port map( A1 => n8200, A2 => n8199, ZN => n8214);
   U1400 : INV_X1 port map( A => n8201, ZN => n8210);
   U1401 : NOR3_X1 port map( A1 => n8225, A2 => n8210, A3 => n8202, ZN => n8207
                           );
   U1402 : INV_X1 port map( A => DATA2(25), ZN => n8865);
   U1403 : NAND2_X1 port map( A1 => DATA1(25), A2 => n8865, ZN => n8694);
   U1404 : NOR2_X1 port map( A1 => DATA1(25), A2 => n8865, ZN => n8622);
   U1405 : INV_X1 port map( A => n8622, ZN => n8690);
   U1406 : AND2_X1 port map( A1 => n8694, A2 => n8690, ZN => n8744);
   U1407 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n8505, ZN
                           => n8205);
   U1408 : NAND3_X1 port map( A1 => n8848, A2 => n8203, A3 => n8271, ZN => 
                           n8204);
   U1409 : OAI211_X1 port map( C1 => n8744, C2 => n8525, A => n8205, B => n8204
                           , ZN => n8206);
   U1410 : AOI211_X1 port map( C1 => dataout_mul_25_port, C2 => n8530, A => 
                           n8207, B => n8206, ZN => n8213);
   U1411 : OAI22_X1 port map( A1 => n8832, A2 => n8208, B1 => n8215, B2 => 
                           n8834, ZN => n8211);
   U1412 : AOI22_X1 port map( A1 => n8479, A2 => n8211, B1 => n8210, B2 => 
                           n8209, ZN => n8212);
   U1413 : OAI211_X1 port map( C1 => n8216, C2 => n8214, A => n8213, B => n8212
                           , ZN => OUTALU(25));
   U1414 : INV_X1 port map( A => DATA1(24), ZN => n8228);
   U1415 : INV_X1 port map( A => n8574, ZN => n8415);
   U1416 : AOI22_X1 port map( A1 => DATA2(24), A2 => n8415, B1 => n8224, B2 => 
                           DATA2_I_24_port, ZN => n8227);
   U1417 : NOR3_X1 port map( A1 => n8832, A2 => n8215, A3 => n8547, ZN => n8223
                           );
   U1418 : AOI22_X1 port map( A1 => n8230, A2 => n8271, B1 => n8231, B2 => 
                           n8273, ZN => n8221);
   U1419 : INV_X1 port map( A => DATA2(24), ZN => n8866);
   U1420 : OAI22_X1 port map( A1 => n8228, A2 => DATA2(24), B1 => n8866, B2 => 
                           n8692, ZN => n8719);
   U1421 : AOI22_X1 port map( A1 => dataout_mul_24_port, A2 => n8575, B1 => 
                           n8567, B2 => n8719, ZN => n8220);
   U1422 : INV_X1 port map( A => n8225, ZN => n8217);
   U1423 : NAND3_X1 port map( A1 => n8218, A2 => n8217, A3 => n8216, ZN => 
                           n8219);
   U1424 : OAI211_X1 port map( C1 => n8221, C2 => n8536, A => n8220, B => n8219
                           , ZN => n8222);
   U1425 : AOI211_X1 port map( C1 => n8225, C2 => n8224, A => n8223, B => n8222
                           , ZN => n8226);
   U1426 : OAI221_X1 port map( B1 => n8228, B2 => n8227, C1 => n8228, C2 => 
                           n8527, A => n8226, ZN => OUTALU(24));
   U1427 : AOI222_X1 port map( A1 => n8232, A2 => n8231, B1 => n8273, B2 => 
                           n8230, C1 => n8271, C2 => n8229, ZN => n8262);
   U1428 : INV_X1 port map( A => DATA2(23), ZN => n8867);
   U1429 : NAND2_X1 port map( A1 => DATA1(23), A2 => n8867, ZN => n8687);
   U1430 : NAND2_X1 port map( A1 => DATA2(23), A2 => n8233, ZN => n8686);
   U1431 : AOI21_X1 port map( B1 => n8687, B2 => n8686, A => n8525, ZN => n8235
                           );
   U1432 : NOR3_X1 port map( A1 => n8546, A2 => n8867, A3 => n8233, ZN => n8234
                           );
   U1433 : AOI211_X1 port map( C1 => dataout_mul_23_port, C2 => n8530, A => 
                           n8235, B => n8234, ZN => n8261);
   U1434 : INV_X1 port map( A => n8285, ZN => n8238);
   U1435 : OAI22_X1 port map( A1 => n8553, A2 => n8236, B1 => n8263, B2 => 
                           n8821, ZN => n8237);
   U1436 : AOI21_X1 port map( B1 => n8239, B2 => n8238, A => n8237, ZN => n8240
                           );
   U1437 : OAI21_X1 port map( B1 => n8301, B2 => n8823, A => n8240, ZN => n8259
                           );
   U1438 : NAND2_X1 port map( A1 => n8248, A2 => n8858, ZN => n8378);
   U1439 : INV_X1 port map( A => n8378, ZN => n8427);
   U1440 : AND2_X1 port map( A1 => n8403, A2 => DATA2_I_17_port, ZN => n8242);
   U1441 : NOR2_X1 port map( A1 => n8242, A2 => n8241, ZN => n8380);
   U1442 : OAI21_X1 port map( B1 => n8397, B2 => n8380, A => n8243, ZN => n8361
                           );
   U1443 : OR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => n8244
                           );
   U1444 : OAI21_X1 port map( B1 => n8361, B2 => n8245, A => n8244, ZN => n8300
                           );
   U1445 : OAI21_X1 port map( B1 => n8309, B2 => n8300, A => n8246, ZN => n8281
                           );
   U1446 : INV_X1 port map( A => n8281, ZN => n8283);
   U1447 : NAND2_X1 port map( A1 => n8286, A2 => DATA2_I_21_port, ZN => n8247);
   U1448 : OAI21_X1 port map( B1 => n8283, B2 => n8295, A => n8247, ZN => n8253
                           );
   U1449 : NOR2_X1 port map( A1 => n9190, A2 => n8248, ZN => n8425);
   U1450 : INV_X1 port map( A => n8251, ZN => n8249);
   U1451 : AOI22_X1 port map( A1 => n8427, A2 => n8253, B1 => n8425, B2 => 
                           n8249, ZN => n8265);
   U1452 : NOR3_X1 port map( A1 => n8250, A2 => n8265, A3 => n8264, ZN => n8258
                           );
   U1453 : INV_X1 port map( A => n8250, ZN => n8256);
   U1454 : AOI21_X1 port map( B1 => n8251, B2 => n8425, A => n8264, ZN => n8252
                           );
   U1455 : OAI21_X1 port map( B1 => n8378, B2 => n8253, A => n8252, ZN => n8267
                           );
   U1456 : AOI21_X1 port map( B1 => n8267, B2 => n8255, A => n8256, ZN => n8254
                           );
   U1457 : AOI211_X1 port map( C1 => n8256, C2 => n8255, A => n9190, B => n8254
                           , ZN => n8257);
   U1458 : AOI211_X1 port map( C1 => n8479, C2 => n8259, A => n8258, B => n8257
                           , ZN => n8260);
   U1459 : OAI211_X1 port map( C1 => n8262, C2 => n8536, A => n8261, B => n8260
                           , ZN => OUTALU(23));
   U1460 : INV_X1 port map( A => DATA2(22), ZN => n8868);
   U1461 : AOI22_X1 port map( A1 => DATA1(22), A2 => DATA2(22), B1 => n8868, B2
                           => n8618, ZN => n8682);
   U1462 : AOI22_X1 port map( A1 => dataout_mul_22_port, A2 => n8575, B1 => 
                           n8567, B2 => n8682, ZN => n8280);
   U1463 : OAI222_X1 port map( A1 => n8821, A2 => n8285, B1 => n8817, B2 => 
                           n8301, C1 => n8263, C2 => n8553, ZN => n8268);
   U1464 : NAND2_X1 port map( A1 => n8265, A2 => n8264, ZN => n8266);
   U1465 : AOI22_X1 port map( A1 => n8479, A2 => n8268, B1 => n8267, B2 => 
                           n8266, ZN => n8279);
   U1466 : OAI22_X1 port map( A1 => n8777, A2 => n8270, B1 => n8269, B2 => 
                           n8778, ZN => n8276);
   U1467 : AOI22_X1 port map( A1 => n8273, A2 => n8272, B1 => n8271, B2 => 
                           n8335, ZN => n8274);
   U1468 : INV_X1 port map( A => n8274, ZN => n8275);
   U1469 : OAI21_X1 port map( B1 => n8276, B2 => n8275, A => n8848, ZN => n8278
                           );
   U1470 : NAND3_X1 port map( A1 => DATA2(22), A2 => DATA1(22), A3 => n8505, ZN
                           => n8277);
   U1471 : NAND4_X1 port map( A1 => n8280, A2 => n8279, A3 => n8278, A4 => 
                           n8277, ZN => OUTALU(22));
   U1472 : AOI22_X1 port map( A1 => n8427, A2 => n8281, B1 => n8425, B2 => 
                           n8282, ZN => n8296);
   U1473 : INV_X1 port map( A => n8282, ZN => n8284);
   U1474 : AOI22_X1 port map( A1 => n8284, A2 => n8425, B1 => n8427, B2 => 
                           n8283, ZN => n8294);
   U1475 : OAI22_X1 port map( A1 => n8553, A2 => n8285, B1 => n8301, B2 => 
                           n8821, ZN => n8292);
   U1476 : INV_X1 port map( A => n8527, ZN => n8414);
   U1477 : AOI21_X1 port map( B1 => n8415, B2 => DATA2(21), A => n8414, ZN => 
                           n8290);
   U1478 : INV_X1 port map( A => n8286, ZN => n8289);
   U1479 : NOR2_X1 port map( A1 => DATA2(21), A2 => n8289, ZN => n8683);
   U1480 : NAND2_X1 port map( A1 => n8289, A2 => DATA2(21), ZN => n8684);
   U1481 : INV_X1 port map( A => n8684, ZN => n8616);
   U1482 : OR2_X1 port map( A1 => n8683, A2 => n8616, ZN => n8723);
   U1483 : AOI22_X1 port map( A1 => dataout_mul_21_port, A2 => n8575, B1 => 
                           n8567, B2 => n8723, ZN => n8288);
   U1484 : NAND3_X1 port map( A1 => n8848, A2 => n8522, A3 => n8387, ZN => 
                           n8287);
   U1485 : OAI211_X1 port map( C1 => n8290, C2 => n8289, A => n8288, B => n8287
                           , ZN => n8291);
   U1486 : AOI21_X1 port map( B1 => n8479, B2 => n8292, A => n8291, ZN => n8293
                           );
   U1487 : OAI221_X1 port map( B1 => n8297, B2 => n8296, C1 => n8295, C2 => 
                           n8294, A => n8293, ZN => OUTALU(21));
   U1488 : INV_X1 port map( A => n8309, ZN => n8311);
   U1489 : INV_X1 port map( A => n8425, ZN => n8377);
   U1490 : OAI22_X1 port map( A1 => n8299, A2 => n8377, B1 => n8378, B2 => 
                           n8300, ZN => n8298);
   U1491 : INV_X1 port map( A => n8298, ZN => n8310);
   U1492 : AOI22_X1 port map( A1 => n8427, A2 => n8300, B1 => n8425, B2 => 
                           n8299, ZN => n8308);
   U1493 : INV_X1 port map( A => DATA2(20), ZN => n8870);
   U1494 : OAI21_X1 port map( B1 => n8574, B2 => n8870, A => n8527, ZN => n8306
                           );
   U1495 : NOR3_X1 port map( A1 => n8553, A2 => n8301, A3 => n8547, ZN => n8305
                           );
   U1496 : AOI22_X1 port map( A1 => n8524, A2 => n8387, B1 => n8522, B2 => 
                           n8386, ZN => n8303);
   U1497 : NAND2_X1 port map( A1 => n8870, A2 => DATA1(20), ZN => n8613);
   U1498 : OAI21_X1 port map( B1 => DATA1(20), B2 => n8870, A => n8613, ZN => 
                           n8721);
   U1499 : AOI22_X1 port map( A1 => dataout_mul_20_port, A2 => n8575, B1 => 
                           n8567, B2 => n8721, ZN => n8302);
   U1500 : OAI21_X1 port map( B1 => n8303, B2 => n8536, A => n8302, ZN => n8304
                           );
   U1501 : AOI211_X1 port map( C1 => DATA1(20), C2 => n8306, A => n8305, B => 
                           n8304, ZN => n8307);
   U1502 : OAI221_X1 port map( B1 => n8311, B2 => n8310, C1 => n8309, C2 => 
                           n8308, A => n8307, ZN => OUTALU(20));
   U1503 : NOR2_X1 port map( A1 => n8312, A2 => n8635, ZN => n8313);
   U1504 : AOI22_X1 port map( A1 => n8575, A2 => dataout_mul_1_port, B1 => 
                           n8479, B2 => n8313, ZN => n8360);
   U1505 : NOR2_X1 port map( A1 => n8314, A2 => DATA2(1), ZN => n8638);
   U1506 : INV_X1 port map( A => n8638, ZN => n8582);
   U1507 : NAND2_X1 port map( A1 => n8314, A2 => DATA2(1), ZN => n8636);
   U1508 : NAND2_X1 port map( A1 => n8582, A2 => n8636, ZN => n8726);
   U1509 : AOI221_X1 port map( B1 => n8316, B2 => n8315, C1 => n8566, C2 => 
                           n8319, A => n8568, ZN => n8322);
   U1510 : AOI211_X1 port map( C1 => n8320, C2 => n8319, A => n8318, B => n8317
                           , ZN => n8321);
   U1511 : AOI211_X1 port map( C1 => n8567, C2 => n8726, A => n8322, B => n8321
                           , ZN => n8359);
   U1512 : AOI21_X1 port map( B1 => n8479, B2 => n8323, A => n8414, ZN => n8573
                           );
   U1513 : OAI21_X1 port map( B1 => n8891, B2 => n8574, A => n8573, ZN => n8357
                           );
   U1514 : INV_X1 port map( A => n8835, ZN => n8356);
   U1515 : INV_X1 port map( A => n8806, ZN => n8345);
   U1516 : AOI22_X1 port map( A1 => n8763, A2 => n8324, B1 => n8762, B2 => 
                           DATA1(1), ZN => n8328);
   U1517 : NAND4_X1 port map( A1 => n8328, A2 => n8327, A3 => n8326, A4 => 
                           n8325, ZN => n8769);
   U1518 : AOI222_X1 port map( A1 => n8329, A2 => n8772, B1 => n8769, B2 => 
                           n8770, C1 => n8773, C2 => n8768, ZN => n8779);
   U1519 : OAI22_X1 port map( A1 => n8777, A2 => n8779, B1 => n8781, B2 => 
                           n8330, ZN => n8334);
   U1520 : OAI22_X1 port map( A1 => n8332, A2 => n8331, B1 => n8775, B2 => 
                           n8778, ZN => n8333);
   U1521 : AOI211_X1 port map( C1 => n8335, C2 => n8784, A => n8334, B => n8333
                           , ZN => n8791);
   U1522 : OAI22_X1 port map( A1 => n8761, A2 => n8788, B1 => n8791, B2 => 
                           n8786, ZN => n8337);
   U1523 : OAI22_X1 port map( A1 => n8792, A2 => n8477, B1 => n8789, B2 => 
                           n8790, ZN => n8336);
   U1524 : AOI211_X1 port map( C1 => n8339, C2 => n8338, A => n8337, B => n8336
                           , ZN => n8802);
   U1525 : OAI222_X1 port map( A1 => n8803, A2 => n8799, B1 => n8801, B2 => 
                           n8802, C1 => n8340, C2 => n8798, ZN => n8810);
   U1526 : AOI22_X1 port map( A1 => n8807, A2 => n8341, B1 => n8805, B2 => 
                           n8810, ZN => n8344);
   U1527 : AOI22_X1 port map( A1 => n8500, A2 => n8808, B1 => n8809, B2 => 
                           n8342, ZN => n8343);
   U1528 : OAI211_X1 port map( C1 => n8345, C2 => n8461, A => n8344, B => n8343
                           , ZN => n8346);
   U1529 : INV_X1 port map( A => n8346, ZN => n8822);
   U1530 : OAI22_X1 port map( A1 => n8817, A2 => n8824, B1 => n8553, B2 => 
                           n8822, ZN => n8350);
   U1531 : OAI22_X1 port map( A1 => n8819, A2 => n8348, B1 => n8823, B2 => 
                           n8347, ZN => n8349);
   U1532 : AOI211_X1 port map( C1 => n8816, C2 => n8351, A => n8350, B => n8349
                           , ZN => n8833);
   U1533 : OAI222_X1 port map( A1 => n8829, A2 => n8352, B1 => n8830, B2 => 
                           n8834, C1 => n8833, C2 => n8832, ZN => n8760);
   U1534 : AOI22_X1 port map( A1 => n8840, A2 => n8841, B1 => n8838, B2 => 
                           n8760, ZN => n8355);
   U1535 : AOI22_X1 port map( A1 => n8842, A2 => n8353, B1 => n8836, B2 => 
                           n8839, ZN => n8354);
   U1536 : OAI211_X1 port map( C1 => n8356, C2 => n8845, A => n8355, B => n8354
                           , ZN => n8851);
   U1537 : AOI22_X1 port map( A1 => DATA1(1), A2 => n8357, B1 => n8848, B2 => 
                           n8851, ZN => n8358);
   U1538 : NAND3_X1 port map( A1 => n8360, A2 => n8359, A3 => n8358, ZN => 
                           OUTALU(1));
   U1539 : INV_X1 port map( A => n8374, ZN => n8376);
   U1540 : AOI22_X1 port map( A1 => n8427, A2 => n8361, B1 => n8425, B2 => 
                           n8362, ZN => n8375);
   U1541 : OAI22_X1 port map( A1 => n8362, A2 => n8377, B1 => n8378, B2 => 
                           n8361, ZN => n8363);
   U1542 : INV_X1 port map( A => n8363, ZN => n8373);
   U1543 : OAI22_X1 port map( A1 => n8463, A2 => n8364, B1 => n8382, B2 => 
                           n8461, ZN => n8371);
   U1544 : OAI22_X1 port map( A1 => n8402, A2 => n8383, B1 => n8422, B2 => 
                           n8814, ZN => n8370);
   U1545 : AOI222_X1 port map( A1 => n8387, A2 => n8496, B1 => n8386, B2 => 
                           n8524, C1 => n8385, C2 => n8522, ZN => n8368);
   U1546 : INV_X1 port map( A => DATA2(19), ZN => n8871);
   U1547 : AND2_X1 port map( A1 => n8871, A2 => DATA1(19), ZN => n8677);
   U1548 : NOR2_X1 port map( A1 => n8365, A2 => n8871, ZN => n8676);
   U1549 : OR2_X1 port map( A1 => n8677, A2 => n8676, ZN => n8731);
   U1550 : AOI22_X1 port map( A1 => dataout_mul_19_port, A2 => n8575, B1 => 
                           n8567, B2 => n8731, ZN => n8367);
   U1551 : OAI211_X1 port map( C1 => n8414, C2 => n8415, A => DATA2(19), B => 
                           DATA1(19), ZN => n8366);
   U1552 : OAI211_X1 port map( C1 => n8368, C2 => n8536, A => n8367, B => n8366
                           , ZN => n8369);
   U1553 : AOI221_X1 port map( B1 => n8371, B2 => n8479, C1 => n8370, C2 => 
                           n8479, A => n8369, ZN => n8372);
   U1554 : OAI221_X1 port map( B1 => n8376, B2 => n8375, C1 => n8374, C2 => 
                           n8373, A => n8372, ZN => OUTALU(19));
   U1555 : INV_X1 port map( A => n8397, ZN => n8399);
   U1556 : OAI22_X1 port map( A1 => n8378, A2 => n8380, B1 => n8377, B2 => 
                           n8381, ZN => n8379);
   U1557 : INV_X1 port map( A => n8379, ZN => n8398);
   U1558 : AOI22_X1 port map( A1 => n8381, A2 => n8425, B1 => n8427, B2 => 
                           n8380, ZN => n8396);
   U1559 : OAI222_X1 port map( A1 => n8383, A2 => n8422, B1 => n8461, B2 => 
                           n8402, C1 => n8382, C2 => n8463, ZN => n8394);
   U1560 : AOI22_X1 port map( A1 => n8524, A2 => n8385, B1 => n8522, B2 => 
                           n8384, ZN => n8389);
   U1561 : AOI22_X1 port map( A1 => n8797, A2 => n8387, B1 => n8496, B2 => 
                           n8386, ZN => n8388);
   U1562 : AOI21_X1 port map( B1 => n8389, B2 => n8388, A => n8536, ZN => n8393
                           );
   U1563 : INV_X1 port map( A => DATA2(18), ZN => n8872);
   U1564 : NOR2_X1 port map( A1 => DATA1(18), A2 => n8872, ZN => n8612);
   U1565 : INV_X1 port map( A => n8612, ZN => n8727);
   U1566 : NAND2_X1 port map( A1 => n8872, A2 => DATA1(18), ZN => n8580);
   U1567 : OAI21_X1 port map( B1 => n8574, B2 => n8872, A => n8527, ZN => n8390
                           );
   U1568 : AOI22_X1 port map( A1 => DATA1(18), A2 => n8390, B1 => n8514, B2 => 
                           dataout_mul_18_port, ZN => n8391);
   U1569 : OAI221_X1 port map( B1 => n8525, B2 => n8727, C1 => n8525, C2 => 
                           n8580, A => n8391, ZN => n8392);
   U1570 : AOI211_X1 port map( C1 => n8479, C2 => n8394, A => n8393, B => n8392
                           , ZN => n8395);
   U1571 : OAI221_X1 port map( B1 => n8399, B2 => n8398, C1 => n8397, C2 => 
                           n8396, A => n8395, ZN => OUTALU(18));
   U1572 : INV_X1 port map( A => n8420, ZN => n8400);
   U1573 : AOI22_X1 port map( A1 => n8421, A2 => n8425, B1 => n8427, B2 => 
                           n8400, ZN => n8412);
   U1574 : AOI22_X1 port map( A1 => n8427, A2 => n8420, B1 => n8425, B2 => 
                           n8401, ZN => n8410);
   U1575 : OAI22_X1 port map( A1 => n8463, A2 => n8402, B1 => n8422, B2 => 
                           n8461, ZN => n8408);
   U1576 : INV_X1 port map( A => DATA2(17), ZN => n8873);
   U1577 : NAND2_X1 port map( A1 => n8873, A2 => n8403, ZN => n8608);
   U1578 : OR2_X1 port map( A1 => n8873, A2 => DATA1(17), ZN => n8673);
   U1579 : NAND2_X1 port map( A1 => n8608, A2 => n8673, ZN => n8724);
   U1580 : AOI22_X1 port map( A1 => dataout_mul_17_port, A2 => n8575, B1 => 
                           n8567, B2 => n8724, ZN => n8406);
   U1581 : NAND3_X1 port map( A1 => n8848, A2 => n8456, A3 => n8416, ZN => 
                           n8405);
   U1582 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n8505, ZN
                           => n8404);
   U1583 : NAND3_X1 port map( A1 => n8406, A2 => n8405, A3 => n8404, ZN => 
                           n8407);
   U1584 : AOI21_X1 port map( B1 => n8479, B2 => n8408, A => n8407, ZN => n8409
                           );
   U1585 : OAI221_X1 port map( B1 => n8413, B2 => n8412, C1 => n8411, C2 => 
                           n8410, A => n8409, ZN => OUTALU(17));
   U1586 : AOI21_X1 port map( B1 => n8415, B2 => DATA2(16), A => n8414, ZN => 
                           n8430);
   U1587 : NOR2_X1 port map( A1 => DATA2(16), A2 => n8671, ZN => n8668);
   U1588 : AOI21_X1 port map( B1 => n8671, B2 => DATA2(16), A => n8668, ZN => 
                           n8735);
   U1589 : AOI22_X1 port map( A1 => n8456, A2 => n8417, B1 => n8431, B2 => 
                           n8416, ZN => n8418);
   U1590 : OAI22_X1 port map( A1 => n8735, A2 => n8525, B1 => n8418, B2 => 
                           n8536, ZN => n8419);
   U1591 : AOI21_X1 port map( B1 => n8514, B2 => dataout_mul_16_port, A => 
                           n8419, ZN => n8429);
   U1592 : NOR2_X1 port map( A1 => n8421, A2 => n8420, ZN => n8424);
   U1593 : INV_X1 port map( A => n8424, ZN => n8426);
   U1594 : NOR3_X1 port map( A1 => n8463, A2 => n8422, A3 => n8547, ZN => n8423
                           );
   U1595 : AOI221_X1 port map( B1 => n8427, B2 => n8426, C1 => n8425, C2 => 
                           n8424, A => n8423, ZN => n8428);
   U1596 : OAI211_X1 port map( C1 => n8430, C2 => n8671, A => n8429, B => n8428
                           , ZN => OUTALU(16));
   U1597 : AOI22_X1 port map( A1 => n8456, A2 => n8432, B1 => n8431, B2 => 
                           n8455, ZN => n8450);
   U1598 : NOR3_X1 port map( A1 => n8463, A2 => n8484, A3 => n8536, ZN => n8439
                           );
   U1599 : XNOR2_X1 port map( A => n8433, B => n8446, ZN => n8437);
   U1600 : NOR2_X1 port map( A1 => DATA2(15), A2 => n8434, ZN => n8667);
   U1601 : INV_X1 port map( A => DATA2(15), ZN => n8875);
   U1602 : NOR2_X1 port map( A1 => DATA1(15), A2 => n8875, ZN => n8631);
   U1603 : OAI21_X1 port map( B1 => n8667, B2 => n8631, A => n8567, ZN => n8436
                           );
   U1604 : NAND3_X1 port map( A1 => DATA2(15), A2 => DATA1(15), A3 => n8505, ZN
                           => n8435);
   U1605 : OAI211_X1 port map( C1 => n8543, C2 => n8437, A => n8436, B => n8435
                           , ZN => n8438);
   U1606 : AOI211_X1 port map( C1 => n8514, C2 => dataout_mul_15_port, A => 
                           n8439, B => n8438, ZN => n8449);
   U1607 : OAI21_X1 port map( B1 => n8561, B2 => n8556, A => n8560, ZN => n8555
                           );
   U1608 : AND2_X1 port map( A1 => n8440, A2 => n8555, ZN => n8531);
   U1609 : OAI21_X1 port map( B1 => n8442, B2 => n8531, A => n8441, ZN => n8516
                           );
   U1610 : AOI21_X1 port map( B1 => n8444, B2 => n8516, A => n8443, ZN => n8464
                           );
   U1611 : NAND2_X1 port map( A1 => n8464, A2 => n8467, ZN => n8453);
   U1612 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n8473, B2 => n8453, ZN => n8447);
   U1613 : AOI21_X1 port map( B1 => n8447, B2 => n8446, A => n8451, ZN => n8445
                           );
   U1614 : OAI21_X1 port map( B1 => n8447, B2 => n8446, A => n8445, ZN => n8448
                           );
   U1615 : OAI211_X1 port map( C1 => n8450, C2 => n8547, A => n8449, B => n8448
                           , ZN => OUTALU(15));
   U1616 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           ZN => n9122);
   U1617 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A => n9122, ZN => n9123);
   U1618 : NOR3_X1 port map( A1 => n5126, A2 => n5134, A3 => n9123, ZN => n3087
                           );
   U1619 : INV_X1 port map( A => n8451, ZN => n8554);
   U1620 : AOI22_X1 port map( A1 => n8554, A2 => n8453, B1 => n8506, B2 => 
                           n8452, ZN => n8472);
   U1621 : AOI221_X1 port map( B1 => n5134, B2 => n5126, C1 => n9123, C2 => 
                           n5126, A => n3087, ZN => n8460);
   U1622 : INV_X1 port map( A => DATA2(14), ZN => n8876);
   U1623 : NOR3_X1 port map( A1 => n8546, A2 => n8876, A3 => n8454, ZN => n8459
                           );
   U1624 : NOR2_X1 port map( A1 => n8876, A2 => DATA1(14), ZN => n8632);
   U1625 : INV_X1 port map( A => n8632, ZN => n8603);
   U1626 : NAND2_X1 port map( A1 => n8876, A2 => DATA1(14), ZN => n8665);
   U1627 : NAND3_X1 port map( A1 => n8479, A2 => n8456, A3 => n8455, ZN => 
                           n8457);
   U1628 : OAI221_X1 port map( B1 => n8525, B2 => n8603, C1 => n8525, C2 => 
                           n8665, A => n8457, ZN => n8458);
   U1629 : AOI211_X1 port map( C1 => n8460, C2 => n8530, A => n8459, B => n8458
                           , ZN => n8471);
   U1630 : OAI22_X1 port map( A1 => n8463, A2 => n8462, B1 => n8484, B2 => 
                           n8461, ZN => n8469);
   U1631 : AOI22_X1 port map( A1 => n8465, A2 => n8506, B1 => n8554, B2 => 
                           n8464, ZN => n8494);
   U1632 : NOR2_X1 port map( A1 => n8494, A2 => n8466, ZN => n8468);
   U1633 : AOI22_X1 port map( A1 => n8848, A2 => n8469, B1 => n8468, B2 => 
                           n8467, ZN => n8470);
   U1634 : OAI211_X1 port map( C1 => n8473, C2 => n8472, A => n8471, B => n8470
                           , ZN => OUTALU(14));
   U1635 : NAND2_X1 port map( A1 => n8877, A2 => n9194, ZN => n8666);
   U1636 : NAND2_X1 port map( A1 => DATA2(13), A2 => n8474, ZN => n8662);
   U1637 : AND2_X1 port map( A1 => n8666, A2 => n8662, ZN => n8743);
   U1638 : OAI22_X1 port map( A1 => n8476, A2 => n8786, B1 => n8475, B2 => 
                           n8790, ZN => n8481);
   U1639 : INV_X1 port map( A => n8523, ZN => n8548);
   U1640 : OAI22_X1 port map( A1 => n8478, A2 => n8788, B1 => n8548, B2 => 
                           n8477, ZN => n8480);
   U1641 : OAI21_X1 port map( B1 => n8481, B2 => n8480, A => n8479, ZN => n8483
                           );
   U1642 : NAND3_X1 port map( A1 => DATA2(13), A2 => n9194, A3 => n8505, ZN => 
                           n8482);
   U1643 : OAI211_X1 port map( C1 => n8743, C2 => n8525, A => n8483, B => n8482
                           , ZN => n8490);
   U1644 : INV_X1 port map( A => n8484, ZN => n8499);
   U1645 : AOI222_X1 port map( A1 => n8501, A2 => n8485, B1 => n8499, B2 => 
                           n8807, C1 => n8498, C2 => n8811, ZN => n8488);
   U1646 : INV_X1 port map( A => n8508, ZN => n8517);
   U1647 : NAND2_X1 port map( A1 => n8517, A2 => n8516, ZN => n8515);
   U1648 : OAI211_X1 port map( C1 => n8507, C2 => n8486, A => n8858, B => n8492
                           , ZN => n8487);
   U1649 : OAI22_X1 port map( A1 => n8488, A2 => n8536, B1 => n8515, B2 => 
                           n8487, ZN => n8489);
   U1650 : AOI211_X1 port map( C1 => n8530, C2 => dataout_mul_13_port, A => 
                           n8490, B => n8489, ZN => n8491);
   U1651 : OAI221_X1 port map( B1 => n8494, B2 => n8493, C1 => n8494, C2 => 
                           n8492, A => n8491, ZN => OUTALU(13));
   U1652 : AOI222_X1 port map( A1 => n8523, A2 => n8496, B1 => n8521, B2 => 
                           n8524, C1 => n8495, C2 => n8522, ZN => n8520);
   U1653 : AOI22_X1 port map( A1 => n8807, A2 => n8498, B1 => n8805, B2 => 
                           n8497, ZN => n8503);
   U1654 : AOI22_X1 port map( A1 => n8811, A2 => n8501, B1 => n8500, B2 => 
                           n8499, ZN => n8502);
   U1655 : AOI21_X1 port map( B1 => n8503, B2 => n8502, A => n8536, ZN => n8513
                           );
   U1656 : AOI22_X1 port map( A1 => n8504, A2 => n8878, B1 => DATA2(12), B2 => 
                           n8602, ZN => n8737);
   U1657 : NAND3_X1 port map( A1 => DATA2(12), A2 => DATA1(12), A3 => n8505, ZN
                           => n8511);
   U1658 : INV_X1 port map( A => n8507, ZN => n8509);
   U1659 : OAI221_X1 port map( B1 => n8509, B2 => n8508, C1 => n8507, C2 => 
                           n8517, A => n8506, ZN => n8510);
   U1660 : OAI211_X1 port map( C1 => n8737, C2 => n8525, A => n8511, B => n8510
                           , ZN => n8512);
   U1661 : AOI211_X1 port map( C1 => n8514, C2 => dataout_mul_12_port, A => 
                           n8513, B => n8512, ZN => n8519);
   U1662 : OAI211_X1 port map( C1 => n8517, C2 => n8516, A => n8554, B => n8515
                           , ZN => n8518);
   U1663 : OAI211_X1 port map( C1 => n8520, C2 => n8547, A => n8519, B => n8518
                           , ZN => OUTALU(12));
   U1664 : AOI22_X1 port map( A1 => n8524, A2 => n8523, B1 => n8522, B2 => 
                           n8521, ZN => n8542);
   U1665 : NAND2_X1 port map( A1 => DATA1(11), A2 => n8879, ZN => n8660);
   U1666 : NAND2_X1 port map( A1 => DATA2(11), A2 => n8526, ZN => n8659);
   U1667 : AOI21_X1 port map( B1 => n8660, B2 => n8659, A => n8525, ZN => n8529
                           );
   U1668 : AOI211_X1 port map( C1 => n8527, C2 => n8574, A => n8526, B => n8879
                           , ZN => n8528);
   U1669 : AOI211_X1 port map( C1 => dataout_mul_11_port, C2 => n8530, A => 
                           n8529, B => n8528, ZN => n8541);
   U1670 : INV_X1 port map( A => n8534, ZN => n8532);
   U1671 : XNOR2_X1 port map( A => n8531, B => n8532, ZN => n8539);
   U1672 : INV_X1 port map( A => n8535, ZN => n8533);
   U1673 : AOI221_X1 port map( B1 => n8535, B2 => n8534, C1 => n8533, C2 => 
                           n8532, A => n8543, ZN => n8538);
   U1674 : NOR3_X1 port map( A1 => n8553, A2 => n8551, A3 => n8536, ZN => n8537
                           );
   U1675 : AOI211_X1 port map( C1 => n8539, C2 => n8554, A => n8538, B => n8537
                           , ZN => n8540);
   U1676 : OAI211_X1 port map( C1 => n8542, C2 => n8547, A => n8541, B => n8540
                           , ZN => OUTALU(11));
   U1677 : NOR2_X1 port map( A1 => n8544, A2 => n8543, ZN => n8558);
   U1678 : AOI22_X1 port map( A1 => n8575, A2 => dataout_mul_10_port, B1 => 
                           n8545, B2 => n8558, ZN => n8565);
   U1679 : AOI22_X1 port map( A1 => DATA1(10), A2 => DATA2(10), B1 => n8880, B2
                           => n8599, ZN => n8655);
   U1680 : NOR3_X1 port map( A1 => n8546, A2 => n8880, A3 => n8599, ZN => n8550
                           );
   U1681 : NOR3_X1 port map( A1 => n8548, A2 => n8547, A3 => n8786, ZN => n8549
                           );
   U1682 : AOI211_X1 port map( C1 => n8567, C2 => n8655, A => n8550, B => n8549
                           , ZN => n8564);
   U1683 : OAI22_X1 port map( A1 => n8553, A2 => n8552, B1 => n8551, B2 => 
                           n8821, ZN => n8557);
   U1684 : AND2_X1 port map( A1 => n8555, A2 => n8554, ZN => n8559);
   U1685 : AOI22_X1 port map( A1 => n8848, A2 => n8557, B1 => n8556, B2 => 
                           n8559, ZN => n8563);
   U1686 : OAI22_X1 port map( A1 => n8561, A2 => n8560, B1 => n8559, B2 => 
                           n8558, ZN => n8562);
   U1687 : NAND4_X1 port map( A1 => n8565, A2 => n8564, A3 => n8563, A4 => 
                           n8562, ZN => OUTALU(10));
   U1688 : OAI21_X1 port map( B1 => DATA1(0), B2 => DATA2_I_0_port, A => n8566,
                           ZN => n8571);
   U1689 : OAI22_X1 port map( A1 => n8892, A2 => DATA1(0), B1 => n8635, B2 => 
                           DATA2(0), ZN => n8732);
   U1690 : AND2_X1 port map( A1 => n8732, A2 => n8567, ZN => n8570);
   U1691 : NOR2_X1 port map( A1 => n8568, A2 => n8571, ZN => n8569);
   U1692 : AOI211_X1 port map( C1 => n8572, C2 => n8571, A => n8570, B => n8569
                           , ZN => n8856);
   U1693 : OAI21_X1 port map( B1 => n8892, B2 => n8574, A => n8573, ZN => n8576
                           );
   U1694 : AOI22_X1 port map( A1 => DATA1(0), A2 => n8576, B1 => n8575, B2 => 
                           dataout_mul_0_port, ZN => n8855);
   U1695 : OAI21_X1 port map( B1 => n8577, B2 => DATA2(30), A => n8707, ZN => 
                           n8716);
   U1696 : INV_X1 port map( A => n8716, ZN => n8629);
   U1697 : OAI21_X1 port map( B1 => DATA2(26), B2 => n8579, A => n8578, ZN => 
                           n8718);
   U1698 : NAND2_X1 port map( A1 => n8692, A2 => n8866, ZN => n8621);
   U1699 : INV_X1 port map( A => n8580, ZN => n8733);
   U1700 : NOR2_X1 port map( A1 => n8733, A2 => n8677, ZN => n8611);
   U1701 : INV_X1 port map( A => n8665, ZN => n8581);
   U1702 : NOR2_X1 port map( A1 => n8581, A2 => n8667, ZN => n8736);
   U1703 : INV_X1 port map( A => n8666, ZN => n8605);
   U1704 : NOR2_X1 port map( A1 => DATA2(8), A2 => n8654, ZN => n8596);
   U1705 : AOI21_X1 port map( B1 => DATA1(6), B2 => n8886, A => n8651, ZN => 
                           n8740);
   U1706 : INV_X1 port map( A => n8648, ZN => n8593);
   U1707 : INV_X1 port map( A => n8636, ZN => n8584);
   U1708 : NAND2_X1 port map( A1 => DATA1(0), A2 => n8892, ZN => n8583);
   U1709 : OAI21_X1 port map( B1 => n8584, B2 => n8583, A => n8582, ZN => n8588
                           );
   U1710 : NOR2_X1 port map( A1 => DATA2(2), A2 => n8585, ZN => n8587);
   U1711 : AOI211_X1 port map( C1 => n8742, C2 => n8588, A => n8587, B => n8586
                           , ZN => n8591);
   U1712 : NOR2_X1 port map( A1 => n8639, A2 => n8589, ZN => n8741);
   U1713 : INV_X1 port map( A => n8741, ZN => n8590);
   U1714 : OAI21_X1 port map( B1 => n8591, B2 => n8590, A => n8642, ZN => n8592
                           );
   U1715 : OAI211_X1 port map( C1 => n8593, C2 => n8592, A => n8649, B => n8644
                           , ZN => n8594);
   U1716 : AOI211_X1 port map( C1 => n8740, C2 => n8594, A => n8633, B => n8650
                           , ZN => n8595);
   U1717 : OAI21_X1 port map( B1 => n8596, B2 => n8595, A => n8657, ZN => n8597
                           );
   U1718 : AOI21_X1 port map( B1 => n8598, B2 => n8597, A => n8655, ZN => n8600
                           );
   U1719 : OAI21_X1 port map( B1 => DATA2(10), B2 => n8599, A => n8660, ZN => 
                           n8734);
   U1720 : OAI211_X1 port map( C1 => n8600, C2 => n8734, A => n8737, B => n8659
                           , ZN => n8601);
   U1721 : OAI21_X1 port map( B1 => DATA2(12), B2 => n8602, A => n8601, ZN => 
                           n8604);
   U1722 : OAI211_X1 port map( C1 => n8605, C2 => n8604, A => n8603, B => n8662
                           , ZN => n8607);
   U1723 : INV_X1 port map( A => n8735, ZN => n8606);
   U1724 : AOI211_X1 port map( C1 => n8736, C2 => n8607, A => n8631, B => n8606
                           , ZN => n8609);
   U1725 : INV_X1 port map( A => n8608, ZN => n8672);
   U1726 : AOI221_X1 port map( B1 => n8668, B2 => n8673, C1 => n8609, C2 => 
                           n8673, A => n8672, ZN => n8610);
   U1727 : AOI221_X1 port map( B1 => n8612, B2 => n8611, C1 => n8610, C2 => 
                           n8611, A => n8676, ZN => n8615);
   U1728 : NAND2_X1 port map( A1 => DATA2(20), A2 => n8681, ZN => n8614);
   U1729 : INV_X1 port map( A => n8613, ZN => n8678);
   U1730 : AOI211_X1 port map( C1 => n8615, C2 => n8614, A => n8678, B => n8683
                           , ZN => n8617);
   U1731 : NOR3_X1 port map( A1 => n8617, A2 => n8616, A3 => n8682, ZN => n8619
                           );
   U1732 : OAI21_X1 port map( B1 => DATA2(22), B2 => n8618, A => n8687, ZN => 
                           n8720);
   U1733 : INV_X1 port map( A => n8719, ZN => n8688);
   U1734 : OAI211_X1 port map( C1 => n8619, C2 => n8720, A => n8688, B => n8686
                           , ZN => n8620);
   U1735 : OAI221_X1 port map( B1 => n8622, B2 => n8621, C1 => n8622, C2 => 
                           n8620, A => n8694, ZN => n8623);
   U1736 : OAI221_X1 port map( B1 => n8718, B2 => n8695, C1 => n8718, C2 => 
                           n8623, A => n8630, ZN => n8624);
   U1737 : OAI22_X1 port map( A1 => DATA2(28), A2 => n8700, B1 => n8717, B2 => 
                           n8624, ZN => n8627);
   U1738 : INV_X1 port map( A => n8625, ZN => n8703);
   U1739 : OAI211_X1 port map( C1 => n8702, C2 => n8627, A => n8626, B => n8703
                           , ZN => n8628);
   U1740 : AOI21_X1 port map( B1 => n8629, B2 => n8628, A => n8705, ZN => n8712
                           );
   U1741 : OAI21_X1 port map( B1 => n8864, B2 => DATA1(26), A => n8630, ZN => 
                           n8749);
   U1742 : INV_X1 port map( A => n8749, ZN => n8698);
   U1743 : NOR2_X1 port map( A1 => n8632, A2 => n8631, ZN => n8747);
   U1744 : AOI21_X1 port map( B1 => DATA2(6), B2 => n8634, A => n8633, ZN => 
                           n8713);
   U1745 : NAND2_X1 port map( A1 => DATA2(0), A2 => n8635, ZN => n8637);
   U1746 : OAI21_X1 port map( B1 => n8638, B2 => n8637, A => n8636, ZN => n8641
                           );
   U1747 : NOR2_X1 port map( A1 => DATA1(2), A2 => n8890, ZN => n8640);
   U1748 : AOI211_X1 port map( C1 => n8742, C2 => n8641, A => n8640, B => n8639
                           , ZN => n8646);
   U1749 : NAND2_X1 port map( A1 => n8643, A2 => n8642, ZN => n8722);
   U1750 : OAI211_X1 port map( C1 => n8646, C2 => n8722, A => n8645, B => n8644
                           , ZN => n8647);
   U1751 : NAND3_X1 port map( A1 => n8649, A2 => n8648, A3 => n8647, ZN => 
                           n8652);
   U1752 : AOI211_X1 port map( C1 => n8713, C2 => n8652, A => n8651, B => n8650
                           , ZN => n8653);
   U1753 : AOI21_X1 port map( B1 => DATA2(8), B2 => n8654, A => n8653, ZN => 
                           n8658);
   U1754 : AOI211_X1 port map( C1 => n8658, C2 => n8657, A => n8656, B => n8655
                           , ZN => n8661);
   U1755 : OAI21_X1 port map( B1 => DATA1(10), B2 => n8880, A => n8659, ZN => 
                           n8714);
   U1756 : OAI211_X1 port map( C1 => n8661, C2 => n8714, A => n8737, B => n8660
                           , ZN => n8663);
   U1757 : OAI211_X1 port map( C1 => DATA1(12), C2 => n8878, A => n8663, B => 
                           n8662, ZN => n8664);
   U1758 : NAND3_X1 port map( A1 => n8666, A2 => n8665, A3 => n8664, ZN => 
                           n8669);
   U1759 : AOI211_X1 port map( C1 => n8747, C2 => n8669, A => n8668, B => n8667
                           , ZN => n8670);
   U1760 : AOI21_X1 port map( B1 => DATA2(16), B2 => n8671, A => n8670, ZN => 
                           n8674);
   U1761 : AOI211_X1 port map( C1 => n8674, C2 => n8673, A => n8672, B => n8733
                           , ZN => n8675);
   U1762 : NOR2_X1 port map( A1 => n8676, A2 => n8675, ZN => n8679);
   U1763 : AOI211_X1 port map( C1 => n8679, C2 => n8727, A => n8678, B => n8677
                           , ZN => n8680);
   U1764 : AOI21_X1 port map( B1 => DATA2(20), B2 => n8681, A => n8680, ZN => 
                           n8685);
   U1765 : AOI211_X1 port map( C1 => n8685, C2 => n8684, A => n8683, B => n8682
                           , ZN => n8689);
   U1766 : OAI21_X1 port map( B1 => DATA1(22), B2 => n8868, A => n8686, ZN => 
                           n8750);
   U1767 : OAI211_X1 port map( C1 => n8689, C2 => n8750, A => n8688, B => n8687
                           , ZN => n8691);
   U1768 : OAI211_X1 port map( C1 => n8692, C2 => n8866, A => n8691, B => n8690
                           , ZN => n8693);
   U1769 : NAND3_X1 port map( A1 => n8695, A2 => n8694, A3 => n8693, ZN => 
                           n8697);
   U1770 : AOI211_X1 port map( C1 => n8698, C2 => n8697, A => n8696, B => n8717
                           , ZN => n8699);
   U1771 : AOI21_X1 port map( B1 => DATA2(28), B2 => n8700, A => n8699, ZN => 
                           n8704);
   U1772 : AOI211_X1 port map( C1 => n8704, C2 => n8703, A => n8702, B => n8701
                           , ZN => n8708);
   U1773 : INV_X1 port map( A => n8705, ZN => n8706);
   U1774 : OAI21_X1 port map( B1 => DATA1(30), B2 => n8860, A => n8706, ZN => 
                           n8748);
   U1775 : OAI211_X1 port map( C1 => n8708, C2 => n8748, A => n8857, B => n8707
                           , ZN => n8710);
   U1776 : OAI211_X1 port map( C1 => FUNC(2), C2 => n8710, A => FUNC(0), B => 
                           n8709, ZN => n8711);
   U1777 : AOI221_X1 port map( B1 => FUNC(2), B2 => FUNC(3), C1 => n8712, C2 =>
                           FUNC(3), A => n8711, ZN => n8850);
   U1778 : INV_X1 port map( A => n8713, ZN => n8715);
   U1779 : NOR4_X1 port map( A1 => n8717, A2 => n8716, A3 => n8715, A4 => n8714
                           , ZN => n8759);
   U1780 : NOR4_X1 port map( A1 => n8721, A2 => n8720, A3 => n8719, A4 => n8718
                           , ZN => n8758);
   U1781 : INV_X1 port map( A => n8722, ZN => n8729);
   U1782 : NOR4_X1 port map( A1 => n8726, A2 => n8725, A3 => n8724, A4 => n8723
                           , ZN => n8728);
   U1783 : NAND4_X1 port map( A1 => FUNC(2), A2 => n8729, A3 => n8728, A4 => 
                           n8727, ZN => n8730);
   U1784 : NOR4_X1 port map( A1 => n8733, A2 => n8732, A3 => n8731, A4 => n8730
                           , ZN => n8757);
   U1785 : INV_X1 port map( A => n8734, ZN => n8738);
   U1786 : NAND4_X1 port map( A1 => n8738, A2 => n8737, A3 => n8736, A4 => 
                           n8735, ZN => n8755);
   U1787 : NAND4_X1 port map( A1 => n8742, A2 => n8741, A3 => n8740, A4 => 
                           n8739, ZN => n8754);
   U1788 : NAND4_X1 port map( A1 => n8746, A2 => n8745, A3 => n8744, A4 => 
                           n8743, ZN => n8753);
   U1789 : INV_X1 port map( A => n8747, ZN => n8751);
   U1790 : OR4_X1 port map( A1 => n8751, A2 => n8750, A3 => n8749, A4 => n8748,
                           ZN => n8752);
   U1791 : NOR4_X1 port map( A1 => n8755, A2 => n8754, A3 => n8753, A4 => n8752
                           , ZN => n8756);
   U1792 : NAND4_X1 port map( A1 => n8759, A2 => n8758, A3 => n8757, A4 => 
                           n8756, ZN => n8849);
   U1793 : INV_X1 port map( A => n8760, ZN => n8846);
   U1794 : INV_X1 port map( A => n8761, ZN => n8796);
   U1795 : AOI22_X1 port map( A1 => n8763, A2 => DATA1(3), B1 => n8762, B2 => 
                           DATA1(0), ZN => n8767);
   U1796 : NAND4_X1 port map( A1 => n8767, A2 => n8766, A3 => n8765, A4 => 
                           n8764, ZN => n8771);
   U1797 : AOI222_X1 port map( A1 => n8773, A2 => n8772, B1 => n8771, B2 => 
                           n8770, C1 => n8769, C2 => n8768, ZN => n8776);
   U1798 : OAI22_X1 port map( A1 => n8777, A2 => n8776, B1 => n8775, B2 => 
                           n8774, ZN => n8783);
   U1799 : OAI22_X1 port map( A1 => n8781, A2 => n8780, B1 => n8779, B2 => 
                           n8778, ZN => n8782);
   U1800 : AOI211_X1 port map( C1 => n8785, C2 => n8784, A => n8783, B => n8782
                           , ZN => n8787);
   U1801 : OAI22_X1 port map( A1 => n8789, A2 => n8788, B1 => n8787, B2 => 
                           n8786, ZN => n8795);
   U1802 : OAI22_X1 port map( A1 => n8793, A2 => n8792, B1 => n8791, B2 => 
                           n8790, ZN => n8794);
   U1803 : AOI211_X1 port map( C1 => n8797, C2 => n8796, A => n8795, B => n8794
                           , ZN => n8800);
   U1804 : OAI222_X1 port map( A1 => n8803, A2 => n8802, B1 => n8801, B2 => 
                           n8800, C1 => n8799, C2 => n8798, ZN => n8804);
   U1805 : AOI22_X1 port map( A1 => n8807, A2 => n8806, B1 => n8805, B2 => 
                           n8804, ZN => n8813);
   U1806 : AOI22_X1 port map( A1 => n8811, A2 => n8810, B1 => n8809, B2 => 
                           n8808, ZN => n8812);
   U1807 : OAI211_X1 port map( C1 => n8815, C2 => n8814, A => n8813, B => n8812
                           , ZN => n8827);
   U1808 : INV_X1 port map( A => n8816, ZN => n8818);
   U1809 : OAI22_X1 port map( A1 => n8820, A2 => n8819, B1 => n8818, B2 => 
                           n8817, ZN => n8826);
   U1810 : OAI22_X1 port map( A1 => n8824, A2 => n8823, B1 => n8822, B2 => 
                           n8821, ZN => n8825);
   U1811 : AOI211_X1 port map( C1 => n8828, C2 => n8827, A => n8826, B => n8825
                           , ZN => n8831);
   U1812 : OAI222_X1 port map( A1 => n8834, A2 => n8833, B1 => n8832, B2 => 
                           n8831, C1 => n8830, C2 => n8829, ZN => n8837);
   U1813 : AOI22_X1 port map( A1 => n8838, A2 => n8837, B1 => n8836, B2 => 
                           n8835, ZN => n8844);
   U1814 : AOI22_X1 port map( A1 => n8842, A2 => n8841, B1 => n8840, B2 => 
                           n8839, ZN => n8843);
   U1815 : OAI211_X1 port map( C1 => n8846, C2 => n8845, A => n8844, B => n8843
                           , ZN => n8847);
   U1816 : AOI22_X1 port map( A1 => n8850, A2 => n8849, B1 => n8848, B2 => 
                           n8847, ZN => n8854);
   U1817 : NAND3_X1 port map( A1 => FUNC(3), A2 => n8852, A3 => n8851, ZN => 
                           n8853);
   U1818 : NAND4_X1 port map( A1 => n8856, A2 => n8855, A3 => n8854, A4 => 
                           n8853, ZN => OUTALU(0));
   U1819 : NAND2_X1 port map( A1 => n8858, A2 => n8857, ZN => n8894);
   U1820 : CLKBUF_X1 port map( A => n8894, Z => n8884);
   U1821 : NAND2_X1 port map( A1 => FUNC(3), A2 => n8858, ZN => n8893);
   U1822 : AOI22_X1 port map( A1 => DATA2(31), A2 => n8884, B1 => n8883, B2 => 
                           n8859, ZN => N2548);
   U1823 : AOI22_X1 port map( A1 => DATA2(30), A2 => n8894, B1 => n8893, B2 => 
                           n8860, ZN => N2547);
   U1824 : AOI22_X1 port map( A1 => DATA2(29), A2 => n8884, B1 => n8883, B2 => 
                           n8861, ZN => N2546);
   U1825 : AOI22_X1 port map( A1 => DATA2(28), A2 => n8894, B1 => n8893, B2 => 
                           n8862, ZN => N2545);
   U1826 : AOI22_X1 port map( A1 => DATA2(27), A2 => n8884, B1 => n8883, B2 => 
                           n8863, ZN => N2544);
   U1827 : AOI22_X1 port map( A1 => DATA2(26), A2 => n8894, B1 => n8893, B2 => 
                           n8864, ZN => N2543);
   U1828 : AOI22_X1 port map( A1 => DATA2(25), A2 => n8884, B1 => n8883, B2 => 
                           n8865, ZN => N2542);
   U1829 : AOI22_X1 port map( A1 => DATA2(24), A2 => n8894, B1 => n8893, B2 => 
                           n8866, ZN => N2541);
   U1830 : AOI22_X1 port map( A1 => DATA2(23), A2 => n8884, B1 => n8883, B2 => 
                           n8867, ZN => N2540);
   U1831 : AOI22_X1 port map( A1 => DATA2(22), A2 => n8894, B1 => n8893, B2 => 
                           n8868, ZN => N2539);
   U1832 : INV_X1 port map( A => DATA2(21), ZN => n8869);
   U1833 : AOI22_X1 port map( A1 => DATA2(21), A2 => n8894, B1 => n8893, B2 => 
                           n8869, ZN => N2538);
   U1834 : AOI22_X1 port map( A1 => DATA2(20), A2 => n8894, B1 => n8893, B2 => 
                           n8870, ZN => N2537);
   U1835 : AOI22_X1 port map( A1 => DATA2(19), A2 => n8884, B1 => n8883, B2 => 
                           n8871, ZN => N2536);
   U1836 : AOI22_X1 port map( A1 => DATA2(18), A2 => n8884, B1 => n8883, B2 => 
                           n8872, ZN => N2535);
   U1837 : AOI22_X1 port map( A1 => DATA2(17), A2 => n8884, B1 => n8883, B2 => 
                           n8873, ZN => N2534);
   U1838 : INV_X1 port map( A => DATA2(16), ZN => n8874);
   U1839 : AOI22_X1 port map( A1 => DATA2(16), A2 => n8884, B1 => n8883, B2 => 
                           n8874, ZN => N2533);
   U1840 : AOI22_X1 port map( A1 => DATA2(15), A2 => n8884, B1 => n8883, B2 => 
                           n8875, ZN => N2532);
   U1841 : AOI22_X1 port map( A1 => DATA2(14), A2 => n8884, B1 => n8883, B2 => 
                           n8876, ZN => N2531);
   U1842 : AOI22_X1 port map( A1 => DATA2(13), A2 => n8884, B1 => n8883, B2 => 
                           n8877, ZN => N2530);
   U1843 : AOI22_X1 port map( A1 => DATA2(12), A2 => n8884, B1 => n8883, B2 => 
                           n8878, ZN => N2529);
   U1844 : AOI22_X1 port map( A1 => DATA2(11), A2 => n8884, B1 => n8883, B2 => 
                           n8879, ZN => N2528);
   U1845 : AOI22_X1 port map( A1 => DATA2(10), A2 => n8884, B1 => n8883, B2 => 
                           n8880, ZN => N2527);
   U1846 : INV_X1 port map( A => DATA2(9), ZN => n8881);
   U1847 : AOI22_X1 port map( A1 => DATA2(9), A2 => n8884, B1 => n8883, B2 => 
                           n8881, ZN => N2526);
   U1848 : AOI22_X1 port map( A1 => DATA2(8), A2 => n8884, B1 => n8883, B2 => 
                           n8882, ZN => N2525);
   U1849 : AOI22_X1 port map( A1 => DATA2(7), A2 => n8894, B1 => n8893, B2 => 
                           n8885, ZN => N2524);
   U1850 : AOI22_X1 port map( A1 => DATA2(6), A2 => n8894, B1 => n8893, B2 => 
                           n8886, ZN => N2523);
   U1851 : AOI22_X1 port map( A1 => DATA2(5), A2 => n8894, B1 => n8893, B2 => 
                           n8887, ZN => N2522);
   U1852 : AOI22_X1 port map( A1 => DATA2(4), A2 => n8894, B1 => n8893, B2 => 
                           n8888, ZN => N2521);
   U1853 : AOI22_X1 port map( A1 => DATA2(3), A2 => n8894, B1 => n8893, B2 => 
                           n8889, ZN => N2520);
   U1854 : AOI22_X1 port map( A1 => DATA2(2), A2 => n8894, B1 => n8893, B2 => 
                           n8890, ZN => N2519);
   U1855 : AOI22_X1 port map( A1 => DATA2(1), A2 => n8894, B1 => n8893, B2 => 
                           n8891, ZN => N2518);
   U1856 : AOI22_X1 port map( A1 => DATA2(0), A2 => n8894, B1 => n8893, B2 => 
                           n8892, ZN => N2517);
   U1857 : NOR2_X1 port map( A1 => n8895, A2 => n1983, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1858 : NAND2_X1 port map( A1 => n8936, A2 => data2_mul_3_port, ZN => n8899)
                           ;
   U1859 : INV_X1 port map( A => data2_mul_3_port, ZN => n8932);
   U1860 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n8932, ZN => n8931);
   U1861 : INV_X1 port map( A => n8896, ZN => n8897);
   U1862 : NOR2_X1 port map( A1 => n8897, A2 => n8932, ZN => n8934);
   U1863 : NOR2_X1 port map( A1 => data2_mul_3_port, A2 => n8897, ZN => n8924);
   U1864 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n8934, B1 => data1_mul_1_port, B2 => n8924, ZN
                           => n8898);
   U1865 : OAI221_X1 port map( B1 => n1983, B2 => n8899, C1 => n1983, C2 => 
                           n8931, A => n8898, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1866 : INV_X1 port map( A => n8899, ZN => n8933);
   U1867 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n8924, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n8933, ZN => n8901);
   U1868 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n8934, ZN => n8900);
   U1869 : OAI211_X1 port map( C1 => n1982, C2 => n8931, A => n8901, B => n8900
                           , ZN => boothmul_pipelined_i_mux_out_1_4_port);
   U1870 : CLKBUF_X1 port map( A => n8924, Z => n8928);
   U1871 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n8933, B1 => n8928, B2 => data1_mul_3_port, ZN
                           => n8903);
   U1872 : CLKBUF_X1 port map( A => n8934, Z => n8925);
   U1873 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n8902);
   U1874 : OAI211_X1 port map( C1 => n8931, C2 => n1980, A => n8903, B => n8902
                           , ZN => boothmul_pipelined_i_mux_out_1_5_port);
   U1875 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n8928, B2 => data1_mul_4_port, ZN => n8905);
   U1876 : NAND2_X1 port map( A1 => n8934, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n8904);
   U1877 : OAI211_X1 port map( C1 => n1979, C2 => n8931, A => n8905, B => n8904
                           , ZN => boothmul_pipelined_i_mux_out_1_6_port);
   U1878 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n8928, B2 => data1_mul_5_port, ZN => n8907);
   U1879 : NAND2_X1 port map( A1 => n8934, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n8906);
   U1880 : OAI211_X1 port map( C1 => n1977, C2 => n8931, A => n8907, B => n8906
                           , ZN => boothmul_pipelined_i_mux_out_1_7_port);
   U1881 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n8928, B2 => data1_mul_6_port, ZN => n8909);
   U1882 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n8908);
   U1883 : OAI211_X1 port map( C1 => n1975, C2 => n8931, A => n8909, B => n8908
                           , ZN => boothmul_pipelined_i_mux_out_1_8_port);
   U1884 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n8924, B2 => data1_mul_7_port, ZN => n8911);
   U1885 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n8910);
   U1886 : OAI211_X1 port map( C1 => n1973, C2 => n8931, A => n8911, B => n8910
                           , ZN => boothmul_pipelined_i_mux_out_1_9_port);
   U1887 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n8924, B2 => data1_mul_8_port, ZN => n8913);
   U1888 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n8912);
   U1889 : OAI211_X1 port map( C1 => n1971, C2 => n8931, A => n8913, B => n8912
                           , ZN => boothmul_pipelined_i_mux_out_1_10_port);
   U1890 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n8928, B2 => data1_mul_9_port, ZN => n8915);
   U1891 : NAND2_X1 port map( A1 => n8934, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n8914);
   U1892 : OAI211_X1 port map( C1 => n1969, C2 => n8931, A => n8915, B => n8914
                           , ZN => boothmul_pipelined_i_mux_out_1_11_port);
   U1893 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n8924, B2 => data1_mul_10_port, ZN => n8917);
   U1894 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n8916);
   U1895 : OAI211_X1 port map( C1 => n1967, C2 => n8931, A => n8917, B => n8916
                           , ZN => boothmul_pipelined_i_mux_out_1_12_port);
   U1896 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n8928, B2 => data1_mul_11_port, ZN => n8919);
   U1897 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n8918);
   U1898 : OAI211_X1 port map( C1 => n1965, C2 => n8931, A => n8919, B => n8918
                           , ZN => boothmul_pipelined_i_mux_out_1_13_port);
   U1899 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n8928, B2 => data1_mul_12_port, ZN => n8921);
   U1900 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n8920);
   U1901 : OAI211_X1 port map( C1 => n1963, C2 => n8931, A => n8921, B => n8920
                           , ZN => boothmul_pipelined_i_mux_out_1_14_port);
   U1902 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n8924, B2 => data1_mul_13_port, ZN => n8923);
   U1903 : NAND2_X1 port map( A1 => n8934, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n8922);
   U1904 : OAI211_X1 port map( C1 => n1961, C2 => n8931, A => n8923, B => n8922
                           , ZN => boothmul_pipelined_i_mux_out_1_15_port);
   U1905 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n8924, B2 => data1_mul_14_port, ZN => n8927);
   U1906 : NAND2_X1 port map( A1 => n8925, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n8926);
   U1907 : OAI211_X1 port map( C1 => n1959, C2 => n8931, A => n8927, B => n8926
                           , ZN => boothmul_pipelined_i_mux_out_1_16_port);
   U1908 : AOI22_X1 port map( A1 => n8933, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n8928, B2 => data1_mul_15_port, ZN => n8930);
   U1909 : NAND2_X1 port map( A1 => n8934, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n8929);
   U1910 : OAI211_X1 port map( C1 => n1957, C2 => n8931, A => n8930, B => n8929
                           , ZN => boothmul_pipelined_i_mux_out_1_17_port);
   U1911 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n8932, ZN => n8937
                           );
   U1912 : AOI22_X1 port map( A1 => n8934, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n8933, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n8935);
   U1913 : OAI21_X1 port map( B1 => n8937, B2 => n8936, A => n8935, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1914 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n8976);
   U1915 : NAND2_X1 port map( A1 => n8976, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n8940);
   U1916 : NAND3_X1 port map( A1 => n3076, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n8972);
   U1917 : NOR2_X1 port map( A1 => n3076, A2 => n8938, ZN => n8953);
   U1918 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n8938, ZN => n8966);
   U1919 : CLKBUF_X1 port map( A => n8966, Z => n8969);
   U1920 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n8953, B1 => data1_mul_1_port, B2 => n8969, ZN
                           => n8939);
   U1921 : OAI221_X1 port map( B1 => n1983, B2 => n8940, C1 => n1983, C2 => 
                           n8972, A => n8939, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1922 : INV_X1 port map( A => n8940, ZN => n8974);
   U1923 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n8966, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n8974, ZN => n8942);
   U1924 : CLKBUF_X1 port map( A => n8953, Z => n8973);
   U1925 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n8973, ZN => n8941);
   U1926 : OAI211_X1 port map( C1 => n8972, C2 => n1982, A => n8942, B => n8941
                           , ZN => boothmul_pipelined_i_mux_out_2_6_port);
   U1927 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n8974, B1 => data1_mul_3_port, B2 => n8969, ZN
                           => n8944);
   U1928 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n8953, ZN => n8943);
   U1929 : OAI211_X1 port map( C1 => n8972, C2 => n1980, A => n8944, B => n8943
                           , ZN => boothmul_pipelined_i_mux_out_2_7_port);
   U1930 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n8974, B1 => data1_mul_4_port, B2 => n8969, ZN
                           => n8946);
   U1931 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n8953, ZN => n8945);
   U1932 : OAI211_X1 port map( C1 => n8972, C2 => n1979, A => n8946, B => n8945
                           , ZN => boothmul_pipelined_i_mux_out_2_8_port);
   U1933 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n8974, B1 => data1_mul_5_port, B2 => n8966, ZN
                           => n8948);
   U1934 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n8953, ZN => n8947);
   U1935 : OAI211_X1 port map( C1 => n8972, C2 => n1977, A => n8948, B => n8947
                           , ZN => boothmul_pipelined_i_mux_out_2_9_port);
   U1936 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n8974, B1 => data1_mul_6_port, B2 => n8969, ZN
                           => n8950);
   U1937 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n8953, ZN => n8949);
   U1938 : OAI211_X1 port map( C1 => n8972, C2 => n1975, A => n8950, B => n8949
                           , ZN => boothmul_pipelined_i_mux_out_2_10_port);
   U1939 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n8974, B1 => data1_mul_7_port, B2 => n8966, ZN
                           => n8952);
   U1940 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n8953, ZN => n8951);
   U1941 : OAI211_X1 port map( C1 => n8972, C2 => n1973, A => n8952, B => n8951
                           , ZN => boothmul_pipelined_i_mux_out_2_11_port);
   U1942 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n8974, B1 => data1_mul_8_port, B2 => n8969, ZN
                           => n8955);
   U1943 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n8953, ZN => n8954);
   U1944 : OAI211_X1 port map( C1 => n8972, C2 => n1971, A => n8955, B => n8954
                           , ZN => boothmul_pipelined_i_mux_out_2_12_port);
   U1945 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n8974, B1 => data1_mul_9_port, B2 => n8969, ZN
                           => n8957);
   U1946 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n8973, ZN => n8956);
   U1947 : OAI211_X1 port map( C1 => n8972, C2 => n1969, A => n8957, B => n8956
                           , ZN => boothmul_pipelined_i_mux_out_2_13_port);
   U1948 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n8974, B1 => data1_mul_10_port, B2 => n8966, 
                           ZN => n8959);
   U1949 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n8973, ZN => n8958);
   U1950 : OAI211_X1 port map( C1 => n8972, C2 => n1967, A => n8959, B => n8958
                           , ZN => boothmul_pipelined_i_mux_out_2_14_port);
   U1951 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n8974, B1 => data1_mul_11_port, B2 => n8966, 
                           ZN => n8961);
   U1952 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n8973, ZN => n8960);
   U1953 : OAI211_X1 port map( C1 => n8972, C2 => n1965, A => n8961, B => n8960
                           , ZN => boothmul_pipelined_i_mux_out_2_15_port);
   U1954 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n8974, B1 => data1_mul_12_port, B2 => n8969, 
                           ZN => n8963);
   U1955 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n8973, ZN => n8962);
   U1956 : OAI211_X1 port map( C1 => n8972, C2 => n1963, A => n8963, B => n8962
                           , ZN => boothmul_pipelined_i_mux_out_2_16_port);
   U1957 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n8974, B1 => data1_mul_13_port, B2 => n8966, 
                           ZN => n8965);
   U1958 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n8973, ZN => n8964);
   U1959 : OAI211_X1 port map( C1 => n8972, C2 => n1961, A => n8965, B => n8964
                           , ZN => boothmul_pipelined_i_mux_out_2_17_port);
   U1960 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n8974, B1 => data1_mul_14_port, B2 => n8966, 
                           ZN => n8968);
   U1961 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n8973, ZN => n8967);
   U1962 : OAI211_X1 port map( C1 => n8972, C2 => n1959, A => n8968, B => n8967
                           , ZN => boothmul_pipelined_i_mux_out_2_18_port);
   U1963 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n8974, B1 => data1_mul_15_port, B2 => n8969, 
                           ZN => n8971);
   U1964 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n8973, ZN => n8970);
   U1965 : OAI211_X1 port map( C1 => n8972, C2 => n1957, A => n8971, B => n8970
                           , ZN => boothmul_pipelined_i_mux_out_2_19_port);
   U1966 : NAND2_X1 port map( A1 => n3076, A2 => data1_mul_15_port, ZN => n8977
                           );
   U1967 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n8974, B1 => n8973, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n8975);
   U1968 : OAI21_X1 port map( B1 => n8977, B2 => n8976, A => n8975, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1969 : NAND3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n9187);
   U1970 : NOR3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n9185);
   U1971 : INV_X1 port map( A => n9185, ZN => n8981);
   U1972 : INV_X1 port map( A => n8979, ZN => n8978);
   U1973 : NAND2_X1 port map( A1 => n3082, A2 => n8978, ZN => n9188);
   U1974 : INV_X1 port map( A => n9188, ZN => n9007);
   U1975 : NOR2_X1 port map( A1 => n3082, A2 => n8979, ZN => n9011);
   U1976 : CLKBUF_X1 port map( A => n9011, Z => n9184);
   U1977 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_176_port, ZN
                           => n8980);
   U1978 : OAI221_X1 port map( B1 => n3077, B2 => n9187, C1 => n3077, C2 => 
                           n8981, A => n8980, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1979 : INV_X1 port map( A => n9187, ZN => n9010);
   U1980 : CLKBUF_X1 port map( A => n9185, Z => n9006);
   U1981 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_3_60_port, A2
                           => n9010, B1 => n9006, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n8983);
   U1982 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n9011
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n8982);
   U1983 : NAND2_X1 port map( A1 => n8983, A2 => n8982, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1984 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n9185
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n8985);
   U1985 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n9011
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n8984);
   U1986 : NAND2_X1 port map( A1 => n8985, A2 => n8984, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1987 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n9185
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n8987);
   U1988 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n9011
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n8986);
   U1989 : NAND2_X1 port map( A1 => n8987, A2 => n8986, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1990 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n8989);
   U1991 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n8988);
   U1992 : NAND2_X1 port map( A1 => n8989, A2 => n8988, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1993 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n8991);
   U1994 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n9011
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n8990);
   U1995 : NAND2_X1 port map( A1 => n8991, A2 => n8990, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1996 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n8993);
   U1997 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n8992);
   U1998 : NAND2_X1 port map( A1 => n8993, A2 => n8992, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1999 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n8995);
   U2000 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n8994);
   U2001 : NAND2_X1 port map( A1 => n8995, A2 => n8994, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U2002 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n8997);
   U2003 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n8996);
   U2004 : NAND2_X1 port map( A1 => n8997, A2 => n8996, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U2005 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n8999);
   U2006 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n9011
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n8998);
   U2007 : NAND2_X1 port map( A1 => n8999, A2 => n8998, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U2008 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n9001);
   U2009 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n9000);
   U2010 : NAND2_X1 port map( A1 => n9001, A2 => n9000, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U2011 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n9003);
   U2012 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n9002);
   U2013 : NAND2_X1 port map( A1 => n9003, A2 => n9002, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U2014 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n9185
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n9005);
   U2015 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n9184
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n9004);
   U2016 : NAND2_X1 port map( A1 => n9005, A2 => n9004, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U2017 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n9006
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n9009);
   U2018 : AOI22_X1 port map( A1 => n9007, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n9011
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n9008);
   U2019 : NAND2_X1 port map( A1 => n9009, A2 => n9008, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U2020 : AOI22_X1 port map( A1 => n9010, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n9185
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n9013);
   U2021 : NAND2_X1 port map( A1 => n9011, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, ZN => 
                           n9012);
   U2022 : OAI211_X1 port map( C1 => n7164, C2 => n9188, A => n9013, B => n9012
                           , ZN => boothmul_pipelined_i_mux_out_3_21_port);
   U2023 : NAND3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n9172);
   U2024 : NOR3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n9170);
   U2025 : INV_X1 port map( A => n9170, ZN => n9017);
   U2026 : INV_X1 port map( A => n9015, ZN => n9014);
   U2027 : NAND2_X1 port map( A1 => n3078, A2 => n9014, ZN => n9173);
   U2028 : INV_X1 port map( A => n9173, ZN => n9043);
   U2029 : NOR2_X1 port map( A1 => n3078, A2 => n9015, ZN => n9047);
   U2030 : CLKBUF_X1 port map( A => n9047, Z => n9169);
   U2031 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_190_port, ZN
                           => n9016);
   U2032 : OAI221_X1 port map( B1 => n5121, B2 => n9172, C1 => n5121, C2 => 
                           n9017, A => n9016, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U2033 : INV_X1 port map( A => n9172, ZN => n9046);
   U2034 : CLKBUF_X1 port map( A => n9170, Z => n9042);
   U2035 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_64_port, A2
                           => n9046, B1 => n9042, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n9019);
   U2036 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n9047
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n9018);
   U2037 : NAND2_X1 port map( A1 => n9019, A2 => n9018, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U2038 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n9170
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n9021);
   U2039 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n9047
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n9020);
   U2040 : NAND2_X1 port map( A1 => n9021, A2 => n9020, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U2041 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n9170
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n9023);
   U2042 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n9047
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n9022);
   U2043 : NAND2_X1 port map( A1 => n9023, A2 => n9022, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2044 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n9025);
   U2045 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n9024);
   U2046 : NAND2_X1 port map( A1 => n9025, A2 => n9024, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2047 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n9027);
   U2048 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n9047
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n9026);
   U2049 : NAND2_X1 port map( A1 => n9027, A2 => n9026, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2050 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n9029);
   U2051 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n9028);
   U2052 : NAND2_X1 port map( A1 => n9029, A2 => n9028, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2053 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n9031);
   U2054 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n9030);
   U2055 : NAND2_X1 port map( A1 => n9031, A2 => n9030, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2056 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n9033);
   U2057 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n9032);
   U2058 : NAND2_X1 port map( A1 => n9033, A2 => n9032, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2059 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n9035);
   U2060 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n9047
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n9034);
   U2061 : NAND2_X1 port map( A1 => n9035, A2 => n9034, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2062 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n9037);
   U2063 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n9036);
   U2064 : NAND2_X1 port map( A1 => n9037, A2 => n9036, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2065 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n9039);
   U2066 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n9038);
   U2067 : NAND2_X1 port map( A1 => n9039, A2 => n9038, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2068 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n9170
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n9041);
   U2069 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n9169
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n9040);
   U2070 : NAND2_X1 port map( A1 => n9041, A2 => n9040, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2071 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n9042
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n9045);
   U2072 : AOI22_X1 port map( A1 => n9043, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n9047
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n9044);
   U2073 : NAND2_X1 port map( A1 => n9045, A2 => n9044, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2074 : AOI22_X1 port map( A1 => n9046, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n9170
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n9049);
   U2075 : NAND2_X1 port map( A1 => n9047, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, ZN => 
                           n9048);
   U2076 : OAI211_X1 port map( C1 => n5127, C2 => n9173, A => n9049, B => n9048
                           , ZN => boothmul_pipelined_i_mux_out_4_23_port);
   U2077 : NAND3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n9177);
   U2078 : NOR3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n9175);
   U2079 : INV_X1 port map( A => n9175, ZN => n9053);
   U2080 : INV_X1 port map( A => n9051, ZN => n9050);
   U2081 : NAND2_X1 port map( A1 => n3079, A2 => n9050, ZN => n9178);
   U2082 : INV_X1 port map( A => n9178, ZN => n9079);
   U2083 : NOR2_X1 port map( A1 => n3079, A2 => n9051, ZN => n9083);
   U2084 : CLKBUF_X1 port map( A => n9083, Z => n9174);
   U2085 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_204_port, ZN
                           => n9052);
   U2086 : OAI221_X1 port map( B1 => n5122, B2 => n9177, C1 => n5122, C2 => 
                           n9053, A => n9052, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2087 : INV_X1 port map( A => n9177, ZN => n9082);
   U2088 : CLKBUF_X1 port map( A => n9175, Z => n9078);
   U2089 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_5_68_port, A2
                           => n9082, B1 => n9078, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n9055);
   U2090 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n9083
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n9054);
   U2091 : NAND2_X1 port map( A1 => n9055, A2 => n9054, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2092 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n9175
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n9057);
   U2093 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n9083
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n9056);
   U2094 : NAND2_X1 port map( A1 => n9057, A2 => n9056, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2095 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n9175
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n9059);
   U2096 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n9083
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n9058);
   U2097 : NAND2_X1 port map( A1 => n9059, A2 => n9058, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2098 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n9061);
   U2099 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n9060);
   U2100 : NAND2_X1 port map( A1 => n9061, A2 => n9060, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2101 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n9063);
   U2102 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n9083
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n9062);
   U2103 : NAND2_X1 port map( A1 => n9063, A2 => n9062, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2104 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n9065);
   U2105 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n9064);
   U2106 : NAND2_X1 port map( A1 => n9065, A2 => n9064, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2107 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n9067);
   U2108 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n9066);
   U2109 : NAND2_X1 port map( A1 => n9067, A2 => n9066, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2110 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n9069);
   U2111 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n9068);
   U2112 : NAND2_X1 port map( A1 => n9069, A2 => n9068, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2113 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n9071);
   U2114 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n9083
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n9070);
   U2115 : NAND2_X1 port map( A1 => n9071, A2 => n9070, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2116 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n9073);
   U2117 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n9072);
   U2118 : NAND2_X1 port map( A1 => n9073, A2 => n9072, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2119 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n9075);
   U2120 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n9074);
   U2121 : NAND2_X1 port map( A1 => n9075, A2 => n9074, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2122 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n9175
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n9077);
   U2123 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n9174
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n9076);
   U2124 : NAND2_X1 port map( A1 => n9077, A2 => n9076, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2125 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n9078
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n9081);
   U2126 : AOI22_X1 port map( A1 => n9079, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n9083
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n9080);
   U2127 : NAND2_X1 port map( A1 => n9081, A2 => n9080, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2128 : AOI22_X1 port map( A1 => n9082, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n9175
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n9085);
   U2129 : NAND2_X1 port map( A1 => n9083, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, ZN => 
                           n9084);
   U2130 : OAI211_X1 port map( C1 => n5128, C2 => n9178, A => n9085, B => n9084
                           , ZN => boothmul_pipelined_i_mux_out_5_25_port);
   U2131 : NAND3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n9182);
   U2132 : NOR3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n9180);
   U2133 : INV_X1 port map( A => n9180, ZN => n9089);
   U2134 : INV_X1 port map( A => n9087, ZN => n9086);
   U2135 : NAND2_X1 port map( A1 => n3080, A2 => n9086, ZN => n9183);
   U2136 : INV_X1 port map( A => n9183, ZN => n9115);
   U2137 : NOR2_X1 port map( A1 => n3080, A2 => n9087, ZN => n9119);
   U2138 : CLKBUF_X1 port map( A => n9119, Z => n9179);
   U2139 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_218_port, ZN
                           => n9088);
   U2140 : OAI221_X1 port map( B1 => n5123, B2 => n9182, C1 => n5123, C2 => 
                           n9089, A => n9088, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2141 : INV_X1 port map( A => n9182, ZN => n9118);
   U2142 : CLKBUF_X1 port map( A => n9180, Z => n9114);
   U2143 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_6_72_port, A2
                           => n9118, B1 => n9114, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n9091);
   U2144 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n9119
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n9090);
   U2145 : NAND2_X1 port map( A1 => n9091, A2 => n9090, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2146 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n9180
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n9093);
   U2147 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n9119
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n9092);
   U2148 : NAND2_X1 port map( A1 => n9093, A2 => n9092, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2149 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n9180
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n9095);
   U2150 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n9119
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n9094);
   U2151 : NAND2_X1 port map( A1 => n9095, A2 => n9094, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2152 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n9097);
   U2153 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n9096);
   U2154 : NAND2_X1 port map( A1 => n9097, A2 => n9096, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2155 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n9099);
   U2156 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n9119
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n9098);
   U2157 : NAND2_X1 port map( A1 => n9099, A2 => n9098, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2158 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n9101);
   U2159 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n9100);
   U2160 : NAND2_X1 port map( A1 => n9101, A2 => n9100, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2161 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n9103);
   U2162 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n9102);
   U2163 : NAND2_X1 port map( A1 => n9103, A2 => n9102, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2164 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n9105);
   U2165 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n9104);
   U2166 : NAND2_X1 port map( A1 => n9105, A2 => n9104, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2167 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n9107);
   U2168 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n9119
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n9106);
   U2169 : NAND2_X1 port map( A1 => n9107, A2 => n9106, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2170 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n9109);
   U2171 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n9108);
   U2172 : NAND2_X1 port map( A1 => n9109, A2 => n9108, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2173 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n9111);
   U2174 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n9110);
   U2175 : NAND2_X1 port map( A1 => n9111, A2 => n9110, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2176 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n9180
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n9113);
   U2177 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n9179
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n9112);
   U2178 : NAND2_X1 port map( A1 => n9113, A2 => n9112, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2179 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n9114
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n9117);
   U2180 : AOI22_X1 port map( A1 => n9115, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n9119
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n9116);
   U2181 : NAND2_X1 port map( A1 => n9117, A2 => n9116, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2182 : AOI22_X1 port map( A1 => n9118, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n9180
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n9121);
   U2183 : NAND2_X1 port map( A1 => n9119, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, ZN => 
                           n9120);
   U2184 : OAI211_X1 port map( C1 => n5129, C2 => n9183, A => n9121, B => n9120
                           , ZN => boothmul_pipelined_i_mux_out_6_27_port);
   U2185 : NOR2_X1 port map( A1 => n9122, A2 => n9189, ZN => n9139);
   U2186 : INV_X1 port map( A => n9139, ZN => n9126);
   U2187 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A3 => n7165, ZN => n9162);
   U2188 : INV_X1 port map( A => n9162, ZN => n9125);
   U2189 : NOR2_X1 port map( A1 => n9123, A2 => n9189, ZN => n9156);
   U2190 : CLKBUF_X1 port map( A => n9156, Z => n9160);
   U2191 : NOR2_X1 port map( A1 => n7165, A2 => n9123, ZN => n9140);
   U2192 : CLKBUF_X1 port map( A => n9140, Z => n9161);
   U2193 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_76_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_232_port, ZN
                           => n9124);
   U2194 : OAI221_X1 port map( B1 => n5134, B2 => n9126, C1 => n5134, C2 => 
                           n9125, A => n9124, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2195 : CLKBUF_X1 port map( A => n9162, Z => n9155);
   U2196 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_7_76_port, A2
                           => n9139, B1 => n9155, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n9128);
   U2197 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n9127);
   U2198 : NAND2_X1 port map( A1 => n9128, A2 => n9127, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2199 : CLKBUF_X1 port map( A => n9139, Z => n9159);
   U2200 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n9162
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n9130);
   U2201 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n9129);
   U2202 : NAND2_X1 port map( A1 => n9130, A2 => n9129, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2203 : AOI22_X1 port map( A1 => n9139, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n9162
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n9132);
   U2204 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n9131);
   U2205 : NAND2_X1 port map( A1 => n9132, A2 => n9131, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2206 : AOI22_X1 port map( A1 => n9139, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n9134);
   U2207 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n9133);
   U2208 : NAND2_X1 port map( A1 => n9134, A2 => n9133, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2209 : AOI22_X1 port map( A1 => n9139, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n9136);
   U2210 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n9135);
   U2211 : NAND2_X1 port map( A1 => n9136, A2 => n9135, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2212 : AOI22_X1 port map( A1 => n9139, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n9138);
   U2213 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n9137);
   U2214 : NAND2_X1 port map( A1 => n9138, A2 => n9137, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2215 : AOI22_X1 port map( A1 => n9139, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n9142);
   U2216 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n9140
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n9141);
   U2217 : NAND2_X1 port map( A1 => n9142, A2 => n9141, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2218 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n9144);
   U2219 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n9143);
   U2220 : NAND2_X1 port map( A1 => n9144, A2 => n9143, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2221 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n9162
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n9146);
   U2222 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n9145);
   U2223 : NAND2_X1 port map( A1 => n9146, A2 => n9145, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2224 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n9148);
   U2225 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n9147);
   U2226 : NAND2_X1 port map( A1 => n9148, A2 => n9147, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2227 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n9150);
   U2228 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n9149);
   U2229 : NAND2_X1 port map( A1 => n9150, A2 => n9149, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2230 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n9152);
   U2231 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n9151);
   U2232 : NAND2_X1 port map( A1 => n9152, A2 => n9151, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2233 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n9162
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n9154);
   U2234 : AOI22_X1 port map( A1 => n9160, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n9153);
   U2235 : NAND2_X1 port map( A1 => n9154, A2 => n9153, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2236 : AOI22_X1 port map( A1 => n9159, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n9155
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n9158);
   U2237 : AOI22_X1 port map( A1 => n9156, A2 => 
                           boothmul_pipelined_i_muxes_in_7_62_port, B1 => n9161
                           , B2 => boothmul_pipelined_i_muxes_in_7_218_port, ZN
                           => n9157);
   U2238 : NAND2_X1 port map( A1 => n9158, A2 => n9157, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2239 : OAI21_X1 port map( B1 => n9160, B2 => n9159, A => 
                           boothmul_pipelined_i_muxes_in_7_62_port, ZN => n9164
                           );
   U2240 : AOI22_X1 port map( A1 => n9162, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n9161, B2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, ZN => 
                           n9163);
   U2241 : NAND2_X1 port map( A1 => n9164, A2 => n9163, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2242 : AOI22_X1 port map( A1 => n9166, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n9165, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n9167);
   U2243 : OAI21_X1 port map( B1 => n9168, B2 => n1955, A => n9167, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2244 : AOI22_X1 port map( A1 => n9170, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, B1 => 
                           n9169, B2 => 
                           boothmul_pipelined_i_muxes_in_4_175_port, ZN => 
                           n9171);
   U2245 : OAI221_X1 port map( B1 => n5127, B2 => n9173, C1 => n5127, C2 => 
                           n9172, A => n9171, ZN => n1997);
   U2246 : AOI22_X1 port map( A1 => n9175, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, B1 => 
                           n9174, B2 => 
                           boothmul_pipelined_i_muxes_in_5_189_port, ZN => 
                           n9176);
   U2247 : OAI221_X1 port map( B1 => n5128, B2 => n9178, C1 => n5128, C2 => 
                           n9177, A => n9176, ZN => n1996);
   U2248 : AOI22_X1 port map( A1 => n9180, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, B1 => 
                           n9179, B2 => 
                           boothmul_pipelined_i_muxes_in_6_203_port, ZN => 
                           n9181);
   U2249 : OAI221_X1 port map( B1 => n5129, B2 => n9183, C1 => n5129, C2 => 
                           n9182, A => n9181, ZN => n1995);
   U2250 : AOI22_X1 port map( A1 => n9185, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, B1 => 
                           n9184, B2 => 
                           boothmul_pipelined_i_muxes_in_3_161_port, ZN => 
                           n9186);
   U2251 : OAI221_X1 port map( B1 => n7164, B2 => n9188, C1 => n7164, C2 => 
                           n9187, A => n9186, ZN => n1991);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, 
      n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, 
      n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, 
      n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, 
      n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, 
      n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, 
      n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, 
      n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, 
      n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, 
      n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, 
      n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, 
      n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, 
      n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, 
      n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, 
      n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, 
      n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, 
      n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, 
      n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, 
      n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, 
      n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, 
      n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, 
      n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, 
      n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, 
      n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, 
      n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, 
      n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, 
      n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, 
      n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, 
      n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, 
      n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, 
      n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, 
      n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, 
      n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, 
      n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, 
      n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, 
      n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, 
      n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, 
      n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, 
      n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, 
      n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, 
      n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, 
      n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, 
      n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, 
      n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, 
      n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, 
      n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, 
      n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, 
      n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, 
      n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, 
      n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, 
      n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, 
      n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, 
      n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, 
      n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
      n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
      n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, 
      n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, 
      n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, 
      n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, 
      n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, 
      n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, 
      n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, 
      n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, 
      n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, 
      n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, 
      n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, 
      n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, 
      n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, 
      n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, 
      n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, 
      n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, 
      n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, 
      n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, 
      n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, 
      n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, 
      n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, 
      n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, 
      n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, 
      n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, 
      n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, 
      n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, 
      n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, 
      n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, 
      n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, 
      n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, 
      n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, 
      n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, 
      n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, 
      n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, 
      n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, 
      n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, 
      n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, 
      n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, 
      n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, 
      n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, 
      n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, 
      n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, 
      n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, 
      n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, 
      n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, 
      n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, 
      n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, 
      n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, 
      n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, 
      n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, 
      n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, 
      n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, 
      n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, 
      n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, 
      n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, 
      n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, 
      n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, 
      n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, 
      n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, 
      n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, 
      n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, 
      n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, 
      n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, 
      n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, 
      n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, 
      n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, 
      n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, 
      n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, 
      n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, 
      n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, 
      n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, 
      n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, 
      n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, 
      n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, 
      n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, 
      n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, 
      n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, 
      n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, 
      n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, 
      n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, 
      n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, 
      n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, 
      n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, 
      n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, 
      n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, 
      n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, 
      n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, 
      n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, 
      n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, 
      n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, 
      n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, 
      n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, 
      n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, 
      n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, 
      n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, 
      n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, 
      n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, 
      n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, 
      n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, 
      n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, 
      n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, 
      n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, 
      n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, 
      n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, 
      n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, 
      n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, 
      n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, 
      n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, 
      n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, 
      n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, 
      n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, 
      n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, 
      n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, 
      n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, 
      n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, 
      n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, 
      n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, 
      n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, 
      n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, 
      n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, 
      n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, 
      n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, 
      n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, 
      n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, 
      n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, 
      n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, 
      n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, 
      n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, 
      n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, 
      n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, 
      n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, 
      n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, 
      n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, 
      n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, 
      n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, 
      n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, 
      n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, 
      n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, 
      n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, 
      n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, 
      n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, 
      n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, 
      n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, 
      n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, 
      n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, 
      n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, 
      n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, 
      n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, 
      n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, 
      n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, 
      n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, 
      n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, 
      n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, 
      n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, 
      n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, 
      n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, 
      n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, 
      n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, 
      n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, 
      n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, 
      n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, 
      n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, 
      n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, 
      n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, 
      n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, 
      n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, 
      n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, 
      n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, 
      n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, 
      n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, 
      n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, 
      n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, 
      n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, 
      n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, 
      n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, 
      n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, 
      n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, 
      n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, 
      n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, 
      n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, 
      n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, 
      n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, 
      n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, 
      n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, 
      n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, 
      n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, 
      n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, 
      n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, 
      n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, 
      n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, 
      n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, 
      n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, 
      n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, 
      n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, 
      n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, 
      n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, 
      n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, 
      n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, 
      n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, 
      n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, 
      n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, 
      n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, 
      n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, 
      n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, 
      n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, 
      n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, 
      n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, 
      n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, 
      n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, 
      n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, 
      n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, 
      n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, 
      n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, 
      n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, 
      n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, 
      n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, 
      n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, 
      n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, 
      n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, 
      n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, 
      n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, 
      n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, 
      n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, 
      n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, 
      n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, 
      n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, 
      n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, 
      n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, 
      n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, 
      n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, 
      n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, 
      n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, 
      n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, 
      n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, 
      n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, 
      n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, 
      n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, 
      n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, 
      n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, 
      n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, 
      n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, 
      n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, 
      n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, 
      n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, 
      n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, 
      n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, 
      n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, 
      n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, 
      n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, 
      n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, 
      n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, 
      n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, 
      n13998, n13999, n14000, n14001, n14002, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412 : std_logic;

begin
   
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n13744);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n12983);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n13252);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n12984);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n13253);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n13745);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n12985);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n13254);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n13255);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n12986);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n12987);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n13256);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n12988);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n12989);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n13257);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n13746);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n13258);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n13500);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n13501);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n12990);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n13747);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n13502);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n12991);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n13259);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n12992);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n12993);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n13260);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n12994);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n13261);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n13748);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n13503);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n13504);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n12995);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n13749);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n13505);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n13750);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n13506);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n12996);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n13751);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n13507);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n13508);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n13509);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n13510);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n13511);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n13752);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n13512);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n12997);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n12998);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n13753);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n12999);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n13513);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n13514);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n13000);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n13001);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n13754);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n13515);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n13516);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n13755);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n13517);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n13002);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n13518);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n13003);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n13004);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n13756);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n13005);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n13262);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n13757);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n13263);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n13758);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n13264);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n13265);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n13519);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n13266);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n13520);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n13006);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n13007);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n13759);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n13760);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n13521);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n13267);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n13761);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n13268);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n13269);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n13008);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n13762);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n13270);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n13522);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n13271);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n13272);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n13763);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n13009);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n13764);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n13273);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n13274);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n13010);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n13275);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n13276);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n13011);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n13277);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n13012);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n13013);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n13014);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n13015);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n13278);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n13279);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n13016);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n13280);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n13017);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n13018);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n13019);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n13020);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n13021);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n13022);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n13023);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n13281);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n13282);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n13024);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n13283);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n13025);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n13026);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n13284);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n13027);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n13028);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n13285);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n13029);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n13523);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n13286);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n13030);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n13765);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n13524);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n13525);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n13526);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n13287);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n13766);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n13767);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n13288);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n13527);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n13289);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n13528);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n13768);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n13290);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n13291);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n13769);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n13529);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n13031);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n13770);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n13032);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n13292);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n13033);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n13771);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n13772);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n13530);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n13531);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n13034);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n13293);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n13532);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n13533);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n13773);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n13774);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n13775);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n13534);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n13776);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n13535);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n13777);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n13778);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n13779);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n13536);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n13780);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n13781);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n13782);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n13783);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n13784);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n13537);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n13785);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n13786);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n13787);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n13538);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n13788);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n13539);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n13789);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n13540);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n13541);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n13790);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n13791);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n13792);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n13542);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n13793);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n13543);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n13544);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n13545);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n13794);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n13546);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n13547);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n13548);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n13035);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n13795);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n13549);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n13550);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n13551);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n13552);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n13553);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n13796);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n13797);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n13798);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n13799);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n13554);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n13555);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n13556);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n13557);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n13558);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n13800);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n13801);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n13802);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n13559);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n13294);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n13560);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n13561);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n13803);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n13562);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n13804);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n13805);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n13036);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n13295);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n13037);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n13296);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n13297);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n13298);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n13038);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n13039);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n13040);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n13299);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n13041);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n13042);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n13300);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n13301);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n13043);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n13044);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n13302);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n13303);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n13304);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n13305);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n13306);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n13307);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n13563);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n13308);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n13309);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n13045);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n13310);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n13311);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n13312);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n13806);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n13313);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n13314);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n13564);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n13315);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n13316);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n13046);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n13807);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n13047);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n13565);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n13317);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n13808);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n13566);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n13318);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n13319);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n13048);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n13049);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n13320);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n13567);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n13050);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n13321);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n13051);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n13052);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n13568);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n13053);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n13809);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n13054);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n13322);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n13055);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n13323);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n13056);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n13569);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n13324);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n13570);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n13057);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n13810);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n13058);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n13811);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n13812);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n13059);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n13813);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n13571);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n13060);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n13061);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n13325);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n13062);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n13572);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n13814);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n13063);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n13573);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n13064);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n13065);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n13066);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n13574);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n13067);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n13068);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n13815);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n13069);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n13816);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n13326);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n13817);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n13327);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n13328);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n13329);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n13818);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n13070);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n13819);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n13330);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n13575);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n13576);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n13071);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n13331);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n13072);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n13332);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n13577);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n13333);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n13073);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n13334);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n13335);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n13336);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n13074);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n13820);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n13821);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n13822);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n13823);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n13578);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n13824);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n13337);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n13338);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n13825);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n13339);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n13075);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n13340);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n13579);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n13826);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n13580);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n13341);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n13827);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n13076);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n13077);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n13342);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n13343);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n13344);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n13345);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n13346);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n13078);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n13079);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n13080);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n13081);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n13082);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n13347);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n13348);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n13349);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n13350);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n13083);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n13084);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n13085);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n13086);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n13087);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n13088);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n13351);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n13089);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n13352);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n13090);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n13353);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n13091);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n13354);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n13092);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n13093);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n13355);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n13094);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n13828);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n13581);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n13095);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n13829);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n13830);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n13582);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n13356);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n13831);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n13583);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n13832);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n13584);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n13585);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n13096);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n13833);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n13097);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n13357);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n13586);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n13358);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n13359);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n13834);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n13835);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n13836);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n13837);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n13587);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n13588);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n13589);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n13838);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n13590);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n13098);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n13591);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n13592);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n13839);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n13593);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n13594);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n13840);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n13595);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n13596);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n13597);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n13841);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n13842);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n13598);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n13843);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n13844);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n13845);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n13599);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n13846);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n13600);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n13601);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n13847);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n13602);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n13848);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n13603);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n13849);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n13604);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n13605);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n13606);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n13607);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n13608);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n13609);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n13850);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n13851);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n13852);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n13610);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n13853);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n13360);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n13854);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n13611);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n13612);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n13613);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n13855);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n13614);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n13615);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n13856);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n13616);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n13617);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n13618);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n13857);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n13619);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n13620);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n13858);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n13859);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n13860);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n13861);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n13862);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n13863);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n13621);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n13099);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n13864);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n13865);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n13622);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n13866);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n13623);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n13867);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n13624);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n13361);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n13625);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n13100);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n13362);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n13101);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n13363);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n13102);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n13364);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n13365);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n13366);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n13367);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n13368);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n13868);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n13103);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n13626);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n13869);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n13369);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n13370);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n13371);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n13627);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n13372);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n13373);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n13104);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n13105);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n13374);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n13106);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n13870);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n13375);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n13107);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n13108);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n13376);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n13109);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n13377);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n13378);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n12979);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n13110);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n13871);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n13628);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n13872);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n13379);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n13380);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n13629);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n13381);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n13873);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n13630);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n13631);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n13111);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n13382);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n13874);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n13383);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n13875);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n13876);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n13384);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n13877);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n13878);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n13879);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n13112);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n13880);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n13385);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n13386);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n13632);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n13113);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n13114);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n13115);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n13881);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n13882);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n13242);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n13883);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n13116);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n13884);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n13633);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n13885);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n13634);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n13886);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n13887);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n13635);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n13387);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n13888);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n13889);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n13636);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n13637);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n13117);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n13638);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n13118);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n13119);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n13890);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n13891);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n13892);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n13893);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n13894);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n13388);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n13639);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n13389);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n13895);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n13896);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n13897);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n13640);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n13641);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n13243);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n13120);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n13642);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n13390);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n13898);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n13121);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n13643);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n13391);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n13899);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n13122);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n13392);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n13123);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n13124);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n13125);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n13126);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n13900);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n13644);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n13901);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n13645);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n13393);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n13394);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n13395);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n13646);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n13396);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n13127);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n13128);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n13397);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n13129);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n13398);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n13647);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n13902);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n13130);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n12980);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n13399);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n13131);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n13132);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n13133);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n13400);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n13401);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n13402);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n13134);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n13135);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n13403);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n13404);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n13136);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n13405);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n13406);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n13137);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n13407);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n13138);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n13408);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n13139);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n13140);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n13409);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n13141);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n13410);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n13142);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n13143);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n13144);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n13411);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n13412);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n13145);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n13413);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n13146);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n13244);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n13903);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n13414);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n13904);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n13648);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n13415);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n13147);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n13649);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n13650);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n13905);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n13906);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n13651);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n13907);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n13416);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n13652);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n13653);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n13654);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n13908);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n13909);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n13910);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n13417);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n13655);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n13911);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n13656);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n13912);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n13913);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n13657);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n13658);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n13659);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n13660);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n13914);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n13661);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n13245);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n13915);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n13662);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n13916);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n13663);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n13917);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n13918);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n13664);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n13665);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n13919);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n13666);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n13920);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n13667);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n13668);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n13669);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n13921);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n13922);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n13670);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n13923);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n13924);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n13671);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n13672);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n13925);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n13673);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n13674);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n13926);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n13927);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n13928);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n13929);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n13930);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n13418);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n13931);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n13495);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n13932);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n13933);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n13934);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n13675);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n13935);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n13676);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n13677);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n13678);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n13936);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n13937);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n13148);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n13679);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n13680);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n13681);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n13682);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n13419);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n13683);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n13684);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n13685);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n13149);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n13686);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n13938);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n13150);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n13420);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n13687);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n13688);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n13939);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n13940);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n13941);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n13689);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n13942);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n12981);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n13151);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n13152);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n13153);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n13154);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n13155);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n13156);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n13943);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n13421);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n13422);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n13157);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n13158);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n13423);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n13159);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n13424);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n13425);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n13160);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n13426);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n13161);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n13427);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n13428);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n13162);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n13429);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n13944);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n13690);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n13163);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n13691);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n13164);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n13692);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n13430);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n13693);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n13165);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n12982);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n13431);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n13694);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n13166);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n13432);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n13167);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n13168);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n13169);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n13170);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n13695);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n13433);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n13434);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n13435);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n13436);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n13437);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n13171);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n13438);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n13439);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n13172);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n13173);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n13696);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n13440);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n13174);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n13441);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n13175);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n13697);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n13176);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n13177);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n13178);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n13442);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n13179);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n13443);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n13246);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n13698);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n13444);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n13180);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n13181);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n13182);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n13445);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n13183);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n13446);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n13184);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n13447);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n13185);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n13945);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n13186);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n13448);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n13699);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n13187);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n13449);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n13700);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n13946);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n13450);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n13188);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n13189);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n13190);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n13191);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n13451);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n13452);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n13701);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n13453);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n13192);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n13193);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n13454);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n13496);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n13194);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n13455);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n13947);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n13948);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n13702);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n13949);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n13950);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n13951);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n13703);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n13704);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n13456);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n13705);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n13952);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n13953);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n13954);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n13706);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n13707);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n13708);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n13709);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n13710);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n13457);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n13195);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n13711);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n13955);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n13458);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n13459);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n13460);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n13712);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n13956);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n13196);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n13197);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n13247);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n13461);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n13198);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n13462);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n13463);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n13199);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n13957);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n13200);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n13464);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n13465);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n13201);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n13958);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n13202);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n13466);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n13203);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n13467);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n13204);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n13713);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n13205);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n13206);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n13207);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n13468);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n13208);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n13209);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n13714);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n13210);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n13469);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n13470);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n13211);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n13212);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n13471);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n13472);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n13248);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n13473);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n13213);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n13715);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n13474);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n13959);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n13214);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n13475);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n13215);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n13216);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n13217);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n13218);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n13219);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n13716);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n13220);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n13960);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n13221);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n13222);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n13476);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n13477);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n13717);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n13718);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n13961);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n13719);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n13720);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n13962);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n13963);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n13721);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n13478);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n13722);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n13964);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n13479);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n13497);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n13723);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n13965);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n13724);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n13966);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n13725);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n13726);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n13967);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n13727);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n13968);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n13969);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n13970);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n13971);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n13972);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n13973);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n13728);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n13974);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n13975);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n13976);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n13729);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n13977);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n13978);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n13730);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n13979);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n13980);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n13981);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n13731);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n13982);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n13732);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n13983);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n13984);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n13985);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n13249);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n13733);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n13986);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n13223);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n13224);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n13734);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n13987);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n13225);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n13988);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n13480);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n13735);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n13736);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n13989);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n13990);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n13991);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n13481);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n13992);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n13482);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n13483);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n13226);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n13993);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n13737);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n13994);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n13484);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n13485);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n13227);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n13995);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n13738);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n13228);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n13229);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n13230);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n13739);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n13498);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n13740);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n13996);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n13486);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n13487);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n13997);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n13488);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n13489);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n13231);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n13232);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n13741);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n13998);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n13490);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n13742);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n13233);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n13234);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n13491);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n13235);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n13999);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n13236);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n13237);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n13238);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n13492);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n13239);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n14000);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n14001);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n13240);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n13493);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n14002);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n13494);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n13241);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n13743);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1349);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1350);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1351);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1352);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1353);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1354);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1355);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1356);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1357);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1358);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1359);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1360);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1361);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1362);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1363);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1364);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1365);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1366);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1367);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1368);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1369);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1370);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1371);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1372);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1373);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1374);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1375);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1376);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1377);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1378);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1379);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1380);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1381);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1382);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1383);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1384);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1385);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1386);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1387);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1388);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1389);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1390);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1391);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1392);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1393);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1394);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1395);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1396);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1397);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1398);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1399);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1400);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1401);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1402);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1403);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1404);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1405);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1406);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1407);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1408);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1409);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1410);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1411);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1412);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n13250);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n13499);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n13251);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n11226);
   U4 : CLKBUF_X1 port map( A => RESET_BAR, Z => n11227);
   U5 : CLKBUF_X1 port map( A => RESET_BAR, Z => n11228);
   U6 : CLKBUF_X1 port map( A => RESET_BAR, Z => n11229);
   U7 : NAND2_X2 port map( A1 => n11229, A2 => n11285, ZN => n11287);
   U8 : NAND2_X2 port map( A1 => n11229, A2 => n11281, ZN => n11283);
   U9 : NAND2_X2 port map( A1 => n11227, A2 => n11278, ZN => n11280);
   U10 : NAND2_X2 port map( A1 => n11229, A2 => n11275, ZN => n11277);
   U11 : NAND2_X2 port map( A1 => n11226, A2 => n11272, ZN => n11274);
   U12 : NAND2_X2 port map( A1 => n11226, A2 => n11269, ZN => n11271);
   U13 : NAND2_X2 port map( A1 => n11229, A2 => n11262, ZN => n11264);
   U14 : NAND2_X2 port map( A1 => n11226, A2 => n11402, ZN => n11414);
   U15 : NAND2_X2 port map( A1 => n11226, A2 => n11375, ZN => n11377);
   U16 : NAND2_X2 port map( A1 => n11229, A2 => n11371, ZN => n11373);
   U17 : NAND2_X2 port map( A1 => n11226, A2 => n11367, ZN => n11369);
   U18 : NAND2_X2 port map( A1 => n11229, A2 => n11363, ZN => n11365);
   U19 : NAND2_X2 port map( A1 => n11229, A2 => n11359, ZN => n11361);
   U20 : NAND2_X2 port map( A1 => n11226, A2 => n11355, ZN => n11357);
   U21 : NAND2_X2 port map( A1 => n11226, A2 => n11344, ZN => n11346);
   U22 : NAND2_X2 port map( A1 => n11227, A2 => n11339, ZN => n11341);
   U23 : NAND2_X2 port map( A1 => n11226, A2 => n11336, ZN => n11338);
   U24 : NAND2_X2 port map( A1 => n11229, A2 => n11329, ZN => n11331);
   U25 : NAND2_X2 port map( A1 => n11228, A2 => n11316, ZN => n11328);
   U26 : NAND2_X2 port map( A1 => n11227, A2 => n11292, ZN => n11294);
   U27 : NAND2_X2 port map( A1 => n11229, A2 => n11289, ZN => n11291);
   U28 : NAND2_X2 port map( A1 => n11226, A2 => n11259, ZN => n11261);
   U29 : NAND2_X2 port map( A1 => n11226, A2 => n11253, ZN => n11255);
   U30 : NAND2_X2 port map( A1 => n11226, A2 => n11249, ZN => n11251);
   U31 : NAND2_X2 port map( A1 => n11226, A2 => n11245, ZN => n11247);
   U32 : INV_X1 port map( A => ADD_WR(4), ZN => n11348);
   U33 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n11256);
   U34 : NOR2_X1 port map( A1 => n11348, A2 => n11347, ZN => n11378);
   U35 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n11288, ZN => n11258);
   U36 : CLKBUF_X1 port map( A => n12196, Z => n12144);
   U37 : CLKBUF_X1 port map( A => n12978, Z => n12924);
   U38 : CLKBUF_X1 port map( A => n11367, Z => n11368);
   U39 : NAND2_X1 port map( A1 => n11227, A2 => n11350, ZN => n11353);
   U40 : NAND2_X1 port map( A1 => n11228, A2 => n11332, ZN => n11335);
   U41 : CLKBUF_X1 port map( A => n11278, Z => n11279);
   U42 : CLKBUF_X1 port map( A => n11317, Z => n11403);
   U43 : CLKBUF_X1 port map( A => n11301, Z => n11387);
   U44 : NAND2_X1 port map( A1 => n11227, A2 => n11265, ZN => n11268);
   U45 : CLKBUF_X1 port map( A => n11253, Z => n11254);
   U46 : CLKBUF_X1 port map( A => n11242, Z => n11243);
   U47 : NAND2_X1 port map( A1 => n11228, A2 => n11235, ZN => n11238);
   U48 : CLKBUF_X1 port map( A => n11234, Z => n11231);
   U49 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n11349);
   U50 : INV_X1 port map( A => ADD_WR(3), ZN => n11230);
   U51 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n11230, ZN => n11288)
                           ;
   U52 : NAND2_X1 port map( A1 => n11349, A2 => n11258, ZN => n11232);
   U53 : CLKBUF_X1 port map( A => n11232, Z => n11233);
   U54 : NAND2_X1 port map( A1 => n11227, A2 => n11233, ZN => n11234);
   U55 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(31), ZN => n11380);
   U56 : CLKBUF_X1 port map( A => n11380, Z => n11343);
   U57 : OAI22_X1 port map( A1 => n13250, A2 => n11231, B1 => n11343, B2 => 
                           n11233, ZN => n2166);
   U58 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(30), ZN => n11295);
   U59 : OAI22_X1 port map( A1 => n13499, A2 => n11234, B1 => n11233, B2 => 
                           n11295, ZN => n2165);
   U60 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(29), ZN => n11296);
   U61 : OAI22_X1 port map( A1 => n13251, A2 => n11231, B1 => n11233, B2 => 
                           n11296, ZN => n2164);
   U62 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(28), ZN => n11297);
   U63 : OAI22_X1 port map( A1 => n13744, A2 => n11234, B1 => n11233, B2 => 
                           n11297, ZN => n2163);
   U64 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(27), ZN => n11298);
   U65 : OAI22_X1 port map( A1 => n12983, A2 => n11231, B1 => n11233, B2 => 
                           n11298, ZN => n2162);
   U66 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(26), ZN => n11299);
   U67 : OAI22_X1 port map( A1 => n13252, A2 => n11234, B1 => n11233, B2 => 
                           n11299, ZN => n2161);
   U68 : NAND2_X1 port map( A1 => n11229, A2 => DATAIN(25), ZN => n11300);
   U69 : OAI22_X1 port map( A1 => n12984, A2 => n11231, B1 => n11233, B2 => 
                           n11300, ZN => n2160);
   U70 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(24), ZN => n11301);
   U71 : OAI22_X1 port map( A1 => n13253, A2 => n11234, B1 => n11233, B2 => 
                           n11301, ZN => n2159);
   U72 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(23), ZN => n11302);
   U73 : OAI22_X1 port map( A1 => n13745, A2 => n11231, B1 => n11232, B2 => 
                           n11302, ZN => n2158);
   U74 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(22), ZN => n11303);
   U75 : OAI22_X1 port map( A1 => n12985, A2 => n11234, B1 => n11232, B2 => 
                           n11303, ZN => n2157);
   U76 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(21), ZN => n11304);
   U77 : OAI22_X1 port map( A1 => n13254, A2 => n11234, B1 => n11232, B2 => 
                           n11304, ZN => n2156);
   U78 : NAND2_X1 port map( A1 => n11229, A2 => DATAIN(20), ZN => n11305);
   U79 : OAI22_X1 port map( A1 => n13255, A2 => n11234, B1 => n11232, B2 => 
                           n11305, ZN => n2155);
   U80 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(19), ZN => n11306);
   U81 : OAI22_X1 port map( A1 => n12986, A2 => n11231, B1 => n11232, B2 => 
                           n11306, ZN => n2154);
   U82 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(18), ZN => n11307);
   U83 : OAI22_X1 port map( A1 => n12987, A2 => n11231, B1 => n11232, B2 => 
                           n11307, ZN => n2153);
   U84 : NAND2_X1 port map( A1 => n11229, A2 => DATAIN(17), ZN => n11308);
   U85 : OAI22_X1 port map( A1 => n13256, A2 => n11231, B1 => n11232, B2 => 
                           n11308, ZN => n2152);
   U86 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(16), ZN => n11309);
   U87 : OAI22_X1 port map( A1 => n12988, A2 => n11231, B1 => n11232, B2 => 
                           n11309, ZN => n2151);
   U88 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(15), ZN => n11310);
   U89 : OAI22_X1 port map( A1 => n12989, A2 => n11231, B1 => n11233, B2 => 
                           n11310, ZN => n2150);
   U90 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(14), ZN => n11311);
   U91 : OAI22_X1 port map( A1 => n13257, A2 => n11231, B1 => n11232, B2 => 
                           n11311, ZN => n2149);
   U92 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(13), ZN => n11312);
   U93 : OAI22_X1 port map( A1 => n13746, A2 => n11231, B1 => n11233, B2 => 
                           n11312, ZN => n2148);
   U94 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(12), ZN => n11313);
   U95 : OAI22_X1 port map( A1 => n13258, A2 => n11231, B1 => n11232, B2 => 
                           n11313, ZN => n2147);
   U96 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(11), ZN => n11314);
   U97 : OAI22_X1 port map( A1 => n13500, A2 => n11231, B1 => n11232, B2 => 
                           n11314, ZN => n2146);
   U98 : NAND2_X1 port map( A1 => n11229, A2 => DATAIN(10), ZN => n11315);
   U99 : OAI22_X1 port map( A1 => n13501, A2 => n11231, B1 => n11232, B2 => 
                           n11315, ZN => n2145);
   U100 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(9), ZN => n11317);
   U101 : OAI22_X1 port map( A1 => n12990, A2 => n11231, B1 => n11233, B2 => 
                           n11317, ZN => n2144);
   U102 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(8), ZN => n11318);
   U103 : OAI22_X1 port map( A1 => n13747, A2 => n11231, B1 => n11232, B2 => 
                           n11318, ZN => n2143);
   U104 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(7), ZN => n11319);
   U105 : OAI22_X1 port map( A1 => n13502, A2 => n11234, B1 => n11233, B2 => 
                           n11319, ZN => n2142);
   U106 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(6), ZN => n11320);
   U107 : OAI22_X1 port map( A1 => n12991, A2 => n11234, B1 => n11232, B2 => 
                           n11320, ZN => n2141);
   U108 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(5), ZN => n11321);
   U109 : OAI22_X1 port map( A1 => n13259, A2 => n11234, B1 => n11233, B2 => 
                           n11321, ZN => n2140);
   U110 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(4), ZN => n11322);
   U111 : OAI22_X1 port map( A1 => n12992, A2 => n11234, B1 => n11232, B2 => 
                           n11322, ZN => n2139);
   U112 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(3), ZN => n11323);
   U113 : OAI22_X1 port map( A1 => n12993, A2 => n11234, B1 => n11233, B2 => 
                           n11323, ZN => n2138);
   U114 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(2), ZN => n11324);
   U115 : OAI22_X1 port map( A1 => n13260, A2 => n11234, B1 => n11232, B2 => 
                           n11324, ZN => n2137);
   U116 : NAND2_X1 port map( A1 => n11227, A2 => DATAIN(1), ZN => n11325);
   U117 : OAI22_X1 port map( A1 => n12994, A2 => n11234, B1 => n11233, B2 => 
                           n11325, ZN => n2136);
   U118 : NAND2_X1 port map( A1 => n11228, A2 => DATAIN(0), ZN => n11327);
   U119 : OAI22_X1 port map( A1 => n13261, A2 => n11234, B1 => n11233, B2 => 
                           n11327, ZN => n2135);
   U120 : INV_X1 port map( A => ADD_WR(0), ZN => n11248);
   U121 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n11248, ZN 
                           => n11354);
   U122 : NAND2_X1 port map( A1 => n11258, A2 => n11354, ZN => n11235);
   U123 : CLKBUF_X1 port map( A => n11238, Z => n11236);
   U124 : CLKBUF_X1 port map( A => n11235, Z => n11237);
   U125 : OAI22_X1 port map( A1 => n13748, A2 => n11236, B1 => n11380, B2 => 
                           n11237, ZN => n2134);
   U126 : OAI22_X1 port map( A1 => n13503, A2 => n11238, B1 => n11295, B2 => 
                           n11235, ZN => n2133);
   U127 : OAI22_X1 port map( A1 => n13504, A2 => n11236, B1 => n11296, B2 => 
                           n11237, ZN => n2132);
   U128 : OAI22_X1 port map( A1 => n12995, A2 => n11238, B1 => n11297, B2 => 
                           n11235, ZN => n2131);
   U129 : OAI22_X1 port map( A1 => n13749, A2 => n11236, B1 => n11298, B2 => 
                           n11237, ZN => n2130);
   U130 : OAI22_X1 port map( A1 => n13505, A2 => n11238, B1 => n11299, B2 => 
                           n11235, ZN => n2129);
   U131 : OAI22_X1 port map( A1 => n13750, A2 => n11236, B1 => n11300, B2 => 
                           n11237, ZN => n2128);
   U132 : OAI22_X1 port map( A1 => n13506, A2 => n11238, B1 => n11301, B2 => 
                           n11235, ZN => n2127);
   U133 : OAI22_X1 port map( A1 => n12996, A2 => n11236, B1 => n11302, B2 => 
                           n11237, ZN => n2126);
   U134 : OAI22_X1 port map( A1 => n13751, A2 => n11238, B1 => n11303, B2 => 
                           n11235, ZN => n2125);
   U135 : OAI22_X1 port map( A1 => n13507, A2 => n11238, B1 => n11304, B2 => 
                           n11235, ZN => n2124);
   U136 : OAI22_X1 port map( A1 => n13508, A2 => n11238, B1 => n11305, B2 => 
                           n11237, ZN => n2123);
   U137 : OAI22_X1 port map( A1 => n13509, A2 => n11236, B1 => n11306, B2 => 
                           n11235, ZN => n2122);
   U138 : OAI22_X1 port map( A1 => n13510, A2 => n11236, B1 => n11307, B2 => 
                           n11237, ZN => n2121);
   U139 : OAI22_X1 port map( A1 => n13511, A2 => n11236, B1 => n11308, B2 => 
                           n11235, ZN => n2120);
   U140 : OAI22_X1 port map( A1 => n13752, A2 => n11236, B1 => n11309, B2 => 
                           n11237, ZN => n2119);
   U141 : OAI22_X1 port map( A1 => n13512, A2 => n11236, B1 => n11310, B2 => 
                           n11235, ZN => n2118);
   U142 : OAI22_X1 port map( A1 => n12997, A2 => n11236, B1 => n11311, B2 => 
                           n11235, ZN => n2117);
   U143 : OAI22_X1 port map( A1 => n12998, A2 => n11236, B1 => n11312, B2 => 
                           n11235, ZN => n2116);
   U144 : OAI22_X1 port map( A1 => n13753, A2 => n11236, B1 => n11313, B2 => 
                           n11235, ZN => n2115);
   U145 : OAI22_X1 port map( A1 => n12999, A2 => n11236, B1 => n11314, B2 => 
                           n11235, ZN => n2114);
   U146 : OAI22_X1 port map( A1 => n13513, A2 => n11236, B1 => n11315, B2 => 
                           n11235, ZN => n2113);
   U147 : OAI22_X1 port map( A1 => n13514, A2 => n11236, B1 => n11317, B2 => 
                           n11235, ZN => n2112);
   U148 : OAI22_X1 port map( A1 => n13000, A2 => n11236, B1 => n11318, B2 => 
                           n11237, ZN => n2111);
   U149 : OAI22_X1 port map( A1 => n13001, A2 => n11238, B1 => n11319, B2 => 
                           n11237, ZN => n2110);
   U150 : OAI22_X1 port map( A1 => n13754, A2 => n11238, B1 => n11320, B2 => 
                           n11237, ZN => n2109);
   U151 : OAI22_X1 port map( A1 => n13515, A2 => n11238, B1 => n11321, B2 => 
                           n11237, ZN => n2108);
   U152 : OAI22_X1 port map( A1 => n13516, A2 => n11238, B1 => n11322, B2 => 
                           n11237, ZN => n2107);
   U153 : OAI22_X1 port map( A1 => n13755, A2 => n11238, B1 => n11323, B2 => 
                           n11237, ZN => n2106);
   U154 : OAI22_X1 port map( A1 => n13517, A2 => n11238, B1 => n11324, B2 => 
                           n11237, ZN => n2105);
   U155 : OAI22_X1 port map( A1 => n13002, A2 => n11238, B1 => n11325, B2 => 
                           n11237, ZN => n2104);
   U156 : OAI22_X1 port map( A1 => n13518, A2 => n11238, B1 => n11327, B2 => 
                           n11237, ZN => n2103);
   U157 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n11248, ZN => n11252);
   U158 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n11252, ZN => n11358);
   U159 : NAND2_X1 port map( A1 => n11258, A2 => n11358, ZN => n11239);
   U160 : NAND2_X2 port map( A1 => n11226, A2 => n11239, ZN => n11241);
   U161 : CLKBUF_X1 port map( A => n11239, Z => n11240);
   U162 : OAI22_X1 port map( A1 => n13003, A2 => n11241, B1 => n11343, B2 => 
                           n11240, ZN => n2102);
   U163 : OAI22_X1 port map( A1 => n13004, A2 => n11241, B1 => n11295, B2 => 
                           n11239, ZN => n2101);
   U164 : OAI22_X1 port map( A1 => n13756, A2 => n11241, B1 => n11296, B2 => 
                           n11240, ZN => n2100);
   U165 : OAI22_X1 port map( A1 => n13005, A2 => n11241, B1 => n11297, B2 => 
                           n11239, ZN => n2099);
   U166 : OAI22_X1 port map( A1 => n13262, A2 => n11241, B1 => n11298, B2 => 
                           n11240, ZN => n2098);
   U167 : OAI22_X1 port map( A1 => n13757, A2 => n11241, B1 => n11299, B2 => 
                           n11239, ZN => n2097);
   U168 : OAI22_X1 port map( A1 => n13263, A2 => n11241, B1 => n11300, B2 => 
                           n11240, ZN => n2096);
   U169 : OAI22_X1 port map( A1 => n13758, A2 => n11241, B1 => n11301, B2 => 
                           n11239, ZN => n2095);
   U170 : OAI22_X1 port map( A1 => n13264, A2 => n11241, B1 => n11302, B2 => 
                           n11240, ZN => n2094);
   U171 : OAI22_X1 port map( A1 => n13265, A2 => n11241, B1 => n11303, B2 => 
                           n11239, ZN => n2093);
   U172 : OAI22_X1 port map( A1 => n13519, A2 => n11241, B1 => n11304, B2 => 
                           n11239, ZN => n2092);
   U173 : OAI22_X1 port map( A1 => n13266, A2 => n11241, B1 => n11305, B2 => 
                           n11240, ZN => n2091);
   U174 : OAI22_X1 port map( A1 => n13520, A2 => n11241, B1 => n11306, B2 => 
                           n11239, ZN => n2090);
   U175 : OAI22_X1 port map( A1 => n13006, A2 => n11241, B1 => n11307, B2 => 
                           n11240, ZN => n2089);
   U176 : OAI22_X1 port map( A1 => n13007, A2 => n11241, B1 => n11308, B2 => 
                           n11239, ZN => n2088);
   U177 : OAI22_X1 port map( A1 => n13759, A2 => n11241, B1 => n11309, B2 => 
                           n11240, ZN => n2087);
   U178 : OAI22_X1 port map( A1 => n13760, A2 => n11241, B1 => n11310, B2 => 
                           n11239, ZN => n2086);
   U179 : OAI22_X1 port map( A1 => n13521, A2 => n11241, B1 => n11311, B2 => 
                           n11239, ZN => n2085);
   U180 : OAI22_X1 port map( A1 => n13267, A2 => n11241, B1 => n11312, B2 => 
                           n11239, ZN => n2084);
   U181 : OAI22_X1 port map( A1 => n13761, A2 => n11241, B1 => n11313, B2 => 
                           n11239, ZN => n2083);
   U182 : OAI22_X1 port map( A1 => n13268, A2 => n11241, B1 => n11314, B2 => 
                           n11239, ZN => n2082);
   U183 : OAI22_X1 port map( A1 => n13269, A2 => n11241, B1 => n11315, B2 => 
                           n11239, ZN => n2081);
   U184 : OAI22_X1 port map( A1 => n13008, A2 => n11241, B1 => n11317, B2 => 
                           n11239, ZN => n2080);
   U185 : OAI22_X1 port map( A1 => n13762, A2 => n11241, B1 => n11318, B2 => 
                           n11240, ZN => n2079);
   U186 : OAI22_X1 port map( A1 => n13270, A2 => n11241, B1 => n11319, B2 => 
                           n11240, ZN => n2078);
   U187 : OAI22_X1 port map( A1 => n13522, A2 => n11241, B1 => n11320, B2 => 
                           n11240, ZN => n2077);
   U188 : OAI22_X1 port map( A1 => n13271, A2 => n11241, B1 => n11321, B2 => 
                           n11240, ZN => n2076);
   U189 : OAI22_X1 port map( A1 => n13272, A2 => n11241, B1 => n11322, B2 => 
                           n11240, ZN => n2075);
   U190 : OAI22_X1 port map( A1 => n13763, A2 => n11241, B1 => n11323, B2 => 
                           n11240, ZN => n2074);
   U191 : OAI22_X1 port map( A1 => n13009, A2 => n11241, B1 => n11324, B2 => 
                           n11240, ZN => n2073);
   U192 : OAI22_X1 port map( A1 => n13764, A2 => n11241, B1 => n11325, B2 => 
                           n11240, ZN => n2072);
   U193 : OAI22_X1 port map( A1 => n13273, A2 => n11241, B1 => n11327, B2 => 
                           n11240, ZN => n2071);
   U194 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n11256, ZN => n11362);
   U195 : NAND2_X1 port map( A1 => n11258, A2 => n11362, ZN => n11242);
   U196 : NAND2_X2 port map( A1 => n11227, A2 => n11242, ZN => n11244);
   U197 : OAI22_X1 port map( A1 => n13274, A2 => n11244, B1 => n11380, B2 => 
                           n11243, ZN => n2070);
   U198 : OAI22_X1 port map( A1 => n13010, A2 => n11244, B1 => n11295, B2 => 
                           n11242, ZN => n2069);
   U199 : OAI22_X1 port map( A1 => n13275, A2 => n11244, B1 => n11296, B2 => 
                           n11243, ZN => n2068);
   U200 : OAI22_X1 port map( A1 => n13276, A2 => n11244, B1 => n11297, B2 => 
                           n11242, ZN => n2067);
   U201 : OAI22_X1 port map( A1 => n13011, A2 => n11244, B1 => n11298, B2 => 
                           n11243, ZN => n2066);
   U202 : OAI22_X1 port map( A1 => n13277, A2 => n11244, B1 => n11299, B2 => 
                           n11242, ZN => n2065);
   U203 : OAI22_X1 port map( A1 => n13012, A2 => n11244, B1 => n11300, B2 => 
                           n11243, ZN => n2064);
   U204 : OAI22_X1 port map( A1 => n13013, A2 => n11244, B1 => n11301, B2 => 
                           n11242, ZN => n2063);
   U205 : OAI22_X1 port map( A1 => n13014, A2 => n11244, B1 => n11302, B2 => 
                           n11243, ZN => n2062);
   U206 : OAI22_X1 port map( A1 => n13015, A2 => n11244, B1 => n11303, B2 => 
                           n11242, ZN => n2061);
   U207 : OAI22_X1 port map( A1 => n13278, A2 => n11244, B1 => n11304, B2 => 
                           n11242, ZN => n2060);
   U208 : OAI22_X1 port map( A1 => n13279, A2 => n11244, B1 => n11305, B2 => 
                           n11243, ZN => n2059);
   U209 : OAI22_X1 port map( A1 => n13016, A2 => n11244, B1 => n11306, B2 => 
                           n11242, ZN => n2058);
   U210 : OAI22_X1 port map( A1 => n13280, A2 => n11244, B1 => n11307, B2 => 
                           n11243, ZN => n2057);
   U211 : OAI22_X1 port map( A1 => n13017, A2 => n11244, B1 => n11308, B2 => 
                           n11242, ZN => n2056);
   U212 : OAI22_X1 port map( A1 => n13018, A2 => n11244, B1 => n11309, B2 => 
                           n11243, ZN => n2055);
   U213 : OAI22_X1 port map( A1 => n13019, A2 => n11244, B1 => n11310, B2 => 
                           n11242, ZN => n2054);
   U214 : OAI22_X1 port map( A1 => n13020, A2 => n11244, B1 => n11311, B2 => 
                           n11242, ZN => n2053);
   U215 : OAI22_X1 port map( A1 => n13021, A2 => n11244, B1 => n11312, B2 => 
                           n11242, ZN => n2052);
   U216 : OAI22_X1 port map( A1 => n13022, A2 => n11244, B1 => n11313, B2 => 
                           n11242, ZN => n2051);
   U217 : OAI22_X1 port map( A1 => n13023, A2 => n11244, B1 => n11314, B2 => 
                           n11242, ZN => n2050);
   U218 : OAI22_X1 port map( A1 => n13281, A2 => n11244, B1 => n11315, B2 => 
                           n11242, ZN => n2049);
   U219 : OAI22_X1 port map( A1 => n13282, A2 => n11244, B1 => n11317, B2 => 
                           n11242, ZN => n2048);
   U220 : OAI22_X1 port map( A1 => n13024, A2 => n11244, B1 => n11318, B2 => 
                           n11243, ZN => n2047);
   U221 : OAI22_X1 port map( A1 => n13283, A2 => n11244, B1 => n11319, B2 => 
                           n11243, ZN => n2046);
   U222 : OAI22_X1 port map( A1 => n13025, A2 => n11244, B1 => n11320, B2 => 
                           n11243, ZN => n2045);
   U223 : OAI22_X1 port map( A1 => n13026, A2 => n11244, B1 => n11321, B2 => 
                           n11243, ZN => n2044);
   U224 : OAI22_X1 port map( A1 => n13284, A2 => n11244, B1 => n11322, B2 => 
                           n11243, ZN => n2043);
   U225 : OAI22_X1 port map( A1 => n13027, A2 => n11244, B1 => n11323, B2 => 
                           n11243, ZN => n2042);
   U226 : OAI22_X1 port map( A1 => n13028, A2 => n11244, B1 => n11324, B2 => 
                           n11243, ZN => n2041);
   U227 : OAI22_X1 port map( A1 => n13285, A2 => n11244, B1 => n11325, B2 => 
                           n11243, ZN => n2040);
   U228 : OAI22_X1 port map( A1 => n13029, A2 => n11244, B1 => n11327, B2 => 
                           n11243, ZN => n2039);
   U229 : INV_X1 port map( A => ADD_WR(2), ZN => n11257);
   U230 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n11257, ZN 
                           => n11366);
   U231 : NAND2_X1 port map( A1 => n11258, A2 => n11366, ZN => n11245);
   U232 : CLKBUF_X1 port map( A => n11245, Z => n11246);
   U233 : OAI22_X1 port map( A1 => n13523, A2 => n11247, B1 => n11343, B2 => 
                           n11246, ZN => n2038);
   U234 : OAI22_X1 port map( A1 => n13286, A2 => n11247, B1 => n11295, B2 => 
                           n11245, ZN => n2037);
   U235 : OAI22_X1 port map( A1 => n13030, A2 => n11247, B1 => n11296, B2 => 
                           n11246, ZN => n2036);
   U236 : OAI22_X1 port map( A1 => n13765, A2 => n11247, B1 => n11297, B2 => 
                           n11245, ZN => n2035);
   U237 : OAI22_X1 port map( A1 => n13524, A2 => n11247, B1 => n11298, B2 => 
                           n11246, ZN => n2034);
   U238 : OAI22_X1 port map( A1 => n13525, A2 => n11247, B1 => n11299, B2 => 
                           n11245, ZN => n2033);
   U239 : OAI22_X1 port map( A1 => n13526, A2 => n11247, B1 => n11300, B2 => 
                           n11246, ZN => n2032);
   U240 : OAI22_X1 port map( A1 => n13287, A2 => n11247, B1 => n11301, B2 => 
                           n11245, ZN => n2031);
   U241 : OAI22_X1 port map( A1 => n13766, A2 => n11247, B1 => n11302, B2 => 
                           n11246, ZN => n2030);
   U242 : OAI22_X1 port map( A1 => n13767, A2 => n11247, B1 => n11303, B2 => 
                           n11245, ZN => n2029);
   U243 : OAI22_X1 port map( A1 => n13288, A2 => n11247, B1 => n11304, B2 => 
                           n11245, ZN => n2028);
   U244 : OAI22_X1 port map( A1 => n13527, A2 => n11247, B1 => n11305, B2 => 
                           n11246, ZN => n2027);
   U245 : OAI22_X1 port map( A1 => n13289, A2 => n11247, B1 => n11306, B2 => 
                           n11245, ZN => n2026);
   U246 : OAI22_X1 port map( A1 => n13528, A2 => n11247, B1 => n11307, B2 => 
                           n11246, ZN => n2025);
   U247 : OAI22_X1 port map( A1 => n13768, A2 => n11247, B1 => n11308, B2 => 
                           n11245, ZN => n2024);
   U248 : OAI22_X1 port map( A1 => n13290, A2 => n11247, B1 => n11309, B2 => 
                           n11246, ZN => n2023);
   U249 : OAI22_X1 port map( A1 => n13291, A2 => n11247, B1 => n11310, B2 => 
                           n11245, ZN => n2022);
   U250 : OAI22_X1 port map( A1 => n13769, A2 => n11247, B1 => n11311, B2 => 
                           n11245, ZN => n2021);
   U251 : OAI22_X1 port map( A1 => n13529, A2 => n11247, B1 => n11312, B2 => 
                           n11245, ZN => n2020);
   U252 : OAI22_X1 port map( A1 => n13031, A2 => n11247, B1 => n11313, B2 => 
                           n11245, ZN => n2019);
   U253 : OAI22_X1 port map( A1 => n13770, A2 => n11247, B1 => n11314, B2 => 
                           n11245, ZN => n2018);
   U254 : OAI22_X1 port map( A1 => n13032, A2 => n11247, B1 => n11315, B2 => 
                           n11245, ZN => n2017);
   U255 : OAI22_X1 port map( A1 => n13292, A2 => n11247, B1 => n11317, B2 => 
                           n11245, ZN => n2016);
   U256 : OAI22_X1 port map( A1 => n13033, A2 => n11247, B1 => n11318, B2 => 
                           n11246, ZN => n2015);
   U257 : OAI22_X1 port map( A1 => n13771, A2 => n11247, B1 => n11319, B2 => 
                           n11246, ZN => n2014);
   U258 : OAI22_X1 port map( A1 => n13772, A2 => n11247, B1 => n11320, B2 => 
                           n11246, ZN => n2013);
   U259 : OAI22_X1 port map( A1 => n13530, A2 => n11247, B1 => n11321, B2 => 
                           n11246, ZN => n2012);
   U260 : OAI22_X1 port map( A1 => n13531, A2 => n11247, B1 => n11322, B2 => 
                           n11246, ZN => n2011);
   U261 : OAI22_X1 port map( A1 => n13034, A2 => n11247, B1 => n11323, B2 => 
                           n11246, ZN => n2010);
   U262 : OAI22_X1 port map( A1 => n13293, A2 => n11247, B1 => n11324, B2 => 
                           n11246, ZN => n2009);
   U263 : OAI22_X1 port map( A1 => n13532, A2 => n11247, B1 => n11325, B2 => 
                           n11246, ZN => n2008);
   U264 : OAI22_X1 port map( A1 => n13533, A2 => n11247, B1 => n11327, B2 => 
                           n11246, ZN => n2007);
   U265 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n11248, A3 => n11257, ZN => 
                           n11370);
   U266 : NAND2_X1 port map( A1 => n11258, A2 => n11370, ZN => n11249);
   U267 : CLKBUF_X1 port map( A => n11249, Z => n11250);
   U268 : OAI22_X1 port map( A1 => n13773, A2 => n11251, B1 => n11380, B2 => 
                           n11250, ZN => n2006);
   U269 : OAI22_X1 port map( A1 => n13774, A2 => n11251, B1 => n11295, B2 => 
                           n11249, ZN => n2005);
   U270 : OAI22_X1 port map( A1 => n13775, A2 => n11251, B1 => n11296, B2 => 
                           n11250, ZN => n2004);
   U271 : OAI22_X1 port map( A1 => n13534, A2 => n11251, B1 => n11297, B2 => 
                           n11249, ZN => n2003);
   U272 : OAI22_X1 port map( A1 => n13776, A2 => n11251, B1 => n11298, B2 => 
                           n11250, ZN => n2002);
   U273 : OAI22_X1 port map( A1 => n13535, A2 => n11251, B1 => n11299, B2 => 
                           n11249, ZN => n2001);
   U274 : OAI22_X1 port map( A1 => n13777, A2 => n11251, B1 => n11300, B2 => 
                           n11250, ZN => n2000);
   U275 : OAI22_X1 port map( A1 => n13778, A2 => n11251, B1 => n11301, B2 => 
                           n11249, ZN => n1999);
   U276 : OAI22_X1 port map( A1 => n13779, A2 => n11251, B1 => n11302, B2 => 
                           n11250, ZN => n1998);
   U277 : OAI22_X1 port map( A1 => n13536, A2 => n11251, B1 => n11303, B2 => 
                           n11249, ZN => n1997);
   U278 : OAI22_X1 port map( A1 => n13780, A2 => n11251, B1 => n11304, B2 => 
                           n11249, ZN => n1996);
   U279 : OAI22_X1 port map( A1 => n13781, A2 => n11251, B1 => n11305, B2 => 
                           n11250, ZN => n1995);
   U280 : OAI22_X1 port map( A1 => n13782, A2 => n11251, B1 => n11306, B2 => 
                           n11249, ZN => n1994);
   U281 : OAI22_X1 port map( A1 => n13783, A2 => n11251, B1 => n11307, B2 => 
                           n11250, ZN => n1993);
   U282 : OAI22_X1 port map( A1 => n13784, A2 => n11251, B1 => n11308, B2 => 
                           n11249, ZN => n1992);
   U283 : OAI22_X1 port map( A1 => n13537, A2 => n11251, B1 => n11309, B2 => 
                           n11250, ZN => n1991);
   U284 : OAI22_X1 port map( A1 => n13785, A2 => n11251, B1 => n11310, B2 => 
                           n11249, ZN => n1990);
   U285 : OAI22_X1 port map( A1 => n13786, A2 => n11251, B1 => n11311, B2 => 
                           n11249, ZN => n1989);
   U286 : OAI22_X1 port map( A1 => n13787, A2 => n11251, B1 => n11312, B2 => 
                           n11249, ZN => n1988);
   U287 : OAI22_X1 port map( A1 => n13538, A2 => n11251, B1 => n11313, B2 => 
                           n11249, ZN => n1987);
   U288 : OAI22_X1 port map( A1 => n13788, A2 => n11251, B1 => n11314, B2 => 
                           n11249, ZN => n1986);
   U289 : OAI22_X1 port map( A1 => n13539, A2 => n11251, B1 => n11315, B2 => 
                           n11249, ZN => n1985);
   U290 : OAI22_X1 port map( A1 => n13789, A2 => n11251, B1 => n11317, B2 => 
                           n11249, ZN => n1984);
   U291 : OAI22_X1 port map( A1 => n13540, A2 => n11251, B1 => n11318, B2 => 
                           n11250, ZN => n1983);
   U292 : OAI22_X1 port map( A1 => n13541, A2 => n11251, B1 => n11319, B2 => 
                           n11250, ZN => n1982);
   U293 : OAI22_X1 port map( A1 => n13790, A2 => n11251, B1 => n11320, B2 => 
                           n11250, ZN => n1981);
   U294 : OAI22_X1 port map( A1 => n13791, A2 => n11251, B1 => n11321, B2 => 
                           n11250, ZN => n1980);
   U295 : OAI22_X1 port map( A1 => n13792, A2 => n11251, B1 => n11322, B2 => 
                           n11250, ZN => n1979);
   U296 : OAI22_X1 port map( A1 => n13542, A2 => n11251, B1 => n11323, B2 => 
                           n11250, ZN => n1978);
   U297 : OAI22_X1 port map( A1 => n13793, A2 => n11251, B1 => n11324, B2 => 
                           n11250, ZN => n1977);
   U298 : OAI22_X1 port map( A1 => n13543, A2 => n11251, B1 => n11325, B2 => 
                           n11250, ZN => n1976);
   U299 : OAI22_X1 port map( A1 => n13544, A2 => n11251, B1 => n11327, B2 => 
                           n11250, ZN => n1975);
   U300 : NOR2_X1 port map( A1 => n11257, A2 => n11252, ZN => n11374);
   U301 : NAND2_X1 port map( A1 => n11258, A2 => n11374, ZN => n11253);
   U302 : OAI22_X1 port map( A1 => n13545, A2 => n11255, B1 => n11343, B2 => 
                           n11254, ZN => n1974);
   U303 : OAI22_X1 port map( A1 => n13794, A2 => n11255, B1 => n11295, B2 => 
                           n11253, ZN => n1973);
   U304 : OAI22_X1 port map( A1 => n13546, A2 => n11255, B1 => n11296, B2 => 
                           n11254, ZN => n1972);
   U305 : OAI22_X1 port map( A1 => n13547, A2 => n11255, B1 => n11297, B2 => 
                           n11253, ZN => n1971);
   U306 : OAI22_X1 port map( A1 => n13548, A2 => n11255, B1 => n11298, B2 => 
                           n11254, ZN => n1970);
   U307 : OAI22_X1 port map( A1 => n13035, A2 => n11255, B1 => n11299, B2 => 
                           n11253, ZN => n1969);
   U308 : OAI22_X1 port map( A1 => n13795, A2 => n11255, B1 => n11300, B2 => 
                           n11254, ZN => n1968);
   U309 : OAI22_X1 port map( A1 => n13549, A2 => n11255, B1 => n11301, B2 => 
                           n11253, ZN => n1967);
   U310 : OAI22_X1 port map( A1 => n13550, A2 => n11255, B1 => n11302, B2 => 
                           n11254, ZN => n1966);
   U311 : OAI22_X1 port map( A1 => n13551, A2 => n11255, B1 => n11303, B2 => 
                           n11253, ZN => n1965);
   U312 : OAI22_X1 port map( A1 => n13552, A2 => n11255, B1 => n11304, B2 => 
                           n11253, ZN => n1964);
   U313 : OAI22_X1 port map( A1 => n13553, A2 => n11255, B1 => n11305, B2 => 
                           n11254, ZN => n1963);
   U314 : OAI22_X1 port map( A1 => n13796, A2 => n11255, B1 => n11306, B2 => 
                           n11253, ZN => n1962);
   U315 : OAI22_X1 port map( A1 => n13797, A2 => n11255, B1 => n11307, B2 => 
                           n11254, ZN => n1961);
   U316 : OAI22_X1 port map( A1 => n13798, A2 => n11255, B1 => n11308, B2 => 
                           n11253, ZN => n1960);
   U317 : OAI22_X1 port map( A1 => n13799, A2 => n11255, B1 => n11309, B2 => 
                           n11254, ZN => n1959);
   U318 : OAI22_X1 port map( A1 => n13554, A2 => n11255, B1 => n11310, B2 => 
                           n11253, ZN => n1958);
   U319 : OAI22_X1 port map( A1 => n13555, A2 => n11255, B1 => n11311, B2 => 
                           n11253, ZN => n1957);
   U320 : OAI22_X1 port map( A1 => n13556, A2 => n11255, B1 => n11312, B2 => 
                           n11253, ZN => n1956);
   U321 : OAI22_X1 port map( A1 => n13557, A2 => n11255, B1 => n11313, B2 => 
                           n11253, ZN => n1955);
   U322 : OAI22_X1 port map( A1 => n13558, A2 => n11255, B1 => n11314, B2 => 
                           n11253, ZN => n1954);
   U323 : OAI22_X1 port map( A1 => n13800, A2 => n11255, B1 => n11315, B2 => 
                           n11253, ZN => n1953);
   U324 : OAI22_X1 port map( A1 => n13801, A2 => n11255, B1 => n11317, B2 => 
                           n11253, ZN => n1952);
   U325 : OAI22_X1 port map( A1 => n13802, A2 => n11255, B1 => n11318, B2 => 
                           n11254, ZN => n1951);
   U326 : OAI22_X1 port map( A1 => n13559, A2 => n11255, B1 => n11319, B2 => 
                           n11254, ZN => n1950);
   U327 : OAI22_X1 port map( A1 => n13294, A2 => n11255, B1 => n11320, B2 => 
                           n11254, ZN => n1949);
   U328 : OAI22_X1 port map( A1 => n13560, A2 => n11255, B1 => n11321, B2 => 
                           n11254, ZN => n1948);
   U329 : OAI22_X1 port map( A1 => n13561, A2 => n11255, B1 => n11322, B2 => 
                           n11254, ZN => n1947);
   U330 : OAI22_X1 port map( A1 => n13803, A2 => n11255, B1 => n11323, B2 => 
                           n11254, ZN => n1946);
   U331 : OAI22_X1 port map( A1 => n13562, A2 => n11255, B1 => n11324, B2 => 
                           n11254, ZN => n1945);
   U332 : OAI22_X1 port map( A1 => n13804, A2 => n11255, B1 => n11325, B2 => 
                           n11254, ZN => n1944);
   U333 : OAI22_X1 port map( A1 => n13805, A2 => n11255, B1 => n11327, B2 => 
                           n11254, ZN => n1943);
   U334 : NOR2_X1 port map( A1 => n11257, A2 => n11256, ZN => n11379);
   U335 : NAND2_X1 port map( A1 => n11258, A2 => n11379, ZN => n11259);
   U336 : CLKBUF_X1 port map( A => n11259, Z => n11260);
   U337 : OAI22_X1 port map( A1 => n13036, A2 => n11261, B1 => n11380, B2 => 
                           n11260, ZN => n1942);
   U338 : OAI22_X1 port map( A1 => n13295, A2 => n11261, B1 => n11295, B2 => 
                           n11259, ZN => n1941);
   U339 : OAI22_X1 port map( A1 => n13037, A2 => n11261, B1 => n11296, B2 => 
                           n11260, ZN => n1940);
   U340 : OAI22_X1 port map( A1 => n13296, A2 => n11261, B1 => n11297, B2 => 
                           n11259, ZN => n1939);
   U341 : OAI22_X1 port map( A1 => n13297, A2 => n11261, B1 => n11298, B2 => 
                           n11260, ZN => n1938);
   U342 : OAI22_X1 port map( A1 => n13298, A2 => n11261, B1 => n11299, B2 => 
                           n11259, ZN => n1937);
   U343 : OAI22_X1 port map( A1 => n13038, A2 => n11261, B1 => n11300, B2 => 
                           n11260, ZN => n1936);
   U344 : OAI22_X1 port map( A1 => n13039, A2 => n11261, B1 => n11301, B2 => 
                           n11259, ZN => n1935);
   U345 : OAI22_X1 port map( A1 => n13040, A2 => n11261, B1 => n11302, B2 => 
                           n11260, ZN => n1934);
   U346 : OAI22_X1 port map( A1 => n13299, A2 => n11261, B1 => n11303, B2 => 
                           n11259, ZN => n1933);
   U347 : OAI22_X1 port map( A1 => n13041, A2 => n11261, B1 => n11304, B2 => 
                           n11259, ZN => n1932);
   U348 : OAI22_X1 port map( A1 => n13042, A2 => n11261, B1 => n11305, B2 => 
                           n11260, ZN => n1931);
   U349 : OAI22_X1 port map( A1 => n13300, A2 => n11261, B1 => n11306, B2 => 
                           n11259, ZN => n1930);
   U350 : OAI22_X1 port map( A1 => n13301, A2 => n11261, B1 => n11307, B2 => 
                           n11260, ZN => n1929);
   U351 : OAI22_X1 port map( A1 => n13043, A2 => n11261, B1 => n11308, B2 => 
                           n11259, ZN => n1928);
   U352 : OAI22_X1 port map( A1 => n13044, A2 => n11261, B1 => n11309, B2 => 
                           n11260, ZN => n1927);
   U353 : OAI22_X1 port map( A1 => n13302, A2 => n11261, B1 => n11310, B2 => 
                           n11259, ZN => n1926);
   U354 : OAI22_X1 port map( A1 => n13303, A2 => n11261, B1 => n11311, B2 => 
                           n11259, ZN => n1925);
   U355 : OAI22_X1 port map( A1 => n13304, A2 => n11261, B1 => n11312, B2 => 
                           n11259, ZN => n1924);
   U356 : OAI22_X1 port map( A1 => n13305, A2 => n11261, B1 => n11313, B2 => 
                           n11259, ZN => n1923);
   U357 : OAI22_X1 port map( A1 => n13306, A2 => n11261, B1 => n11314, B2 => 
                           n11259, ZN => n1922);
   U358 : OAI22_X1 port map( A1 => n13307, A2 => n11261, B1 => n11315, B2 => 
                           n11259, ZN => n1921);
   U359 : OAI22_X1 port map( A1 => n13563, A2 => n11261, B1 => n11317, B2 => 
                           n11259, ZN => n1920);
   U360 : OAI22_X1 port map( A1 => n13308, A2 => n11261, B1 => n11318, B2 => 
                           n11260, ZN => n1919);
   U361 : OAI22_X1 port map( A1 => n13309, A2 => n11261, B1 => n11319, B2 => 
                           n11260, ZN => n1918);
   U362 : OAI22_X1 port map( A1 => n13045, A2 => n11261, B1 => n11320, B2 => 
                           n11260, ZN => n1917);
   U363 : OAI22_X1 port map( A1 => n13310, A2 => n11261, B1 => n11321, B2 => 
                           n11260, ZN => n1916);
   U364 : OAI22_X1 port map( A1 => n13311, A2 => n11261, B1 => n11322, B2 => 
                           n11260, ZN => n1915);
   U365 : OAI22_X1 port map( A1 => n13312, A2 => n11261, B1 => n11323, B2 => 
                           n11260, ZN => n1914);
   U366 : OAI22_X1 port map( A1 => n13806, A2 => n11261, B1 => n11324, B2 => 
                           n11260, ZN => n1913);
   U367 : OAI22_X1 port map( A1 => n13313, A2 => n11261, B1 => n11325, B2 => 
                           n11260, ZN => n1912);
   U368 : OAI22_X1 port map( A1 => n13314, A2 => n11261, B1 => n11327, B2 => 
                           n11260, ZN => n1911);
   U369 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(3), ZN => 
                           n11347);
   U370 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n11347, ZN => n11284);
   U371 : NAND2_X1 port map( A1 => n11349, A2 => n11284, ZN => n11262);
   U372 : CLKBUF_X1 port map( A => n11262, Z => n11263);
   U373 : OAI22_X1 port map( A1 => n13564, A2 => n11264, B1 => n11343, B2 => 
                           n11263, ZN => n1910);
   U374 : OAI22_X1 port map( A1 => n13315, A2 => n11264, B1 => n11295, B2 => 
                           n11262, ZN => n1909);
   U375 : OAI22_X1 port map( A1 => n13316, A2 => n11264, B1 => n11296, B2 => 
                           n11263, ZN => n1908);
   U376 : OAI22_X1 port map( A1 => n13046, A2 => n11264, B1 => n11297, B2 => 
                           n11262, ZN => n1907);
   U377 : OAI22_X1 port map( A1 => n13807, A2 => n11264, B1 => n11298, B2 => 
                           n11263, ZN => n1906);
   U378 : OAI22_X1 port map( A1 => n13047, A2 => n11264, B1 => n11299, B2 => 
                           n11262, ZN => n1905);
   U379 : OAI22_X1 port map( A1 => n13565, A2 => n11264, B1 => n11300, B2 => 
                           n11263, ZN => n1904);
   U380 : OAI22_X1 port map( A1 => n13317, A2 => n11264, B1 => n11301, B2 => 
                           n11262, ZN => n1903);
   U381 : OAI22_X1 port map( A1 => n13808, A2 => n11264, B1 => n11302, B2 => 
                           n11263, ZN => n1902);
   U382 : OAI22_X1 port map( A1 => n13566, A2 => n11264, B1 => n11303, B2 => 
                           n11262, ZN => n1901);
   U383 : OAI22_X1 port map( A1 => n13318, A2 => n11264, B1 => n11304, B2 => 
                           n11262, ZN => n1900);
   U384 : OAI22_X1 port map( A1 => n13319, A2 => n11264, B1 => n11305, B2 => 
                           n11263, ZN => n1899);
   U385 : OAI22_X1 port map( A1 => n13048, A2 => n11264, B1 => n11306, B2 => 
                           n11262, ZN => n1898);
   U386 : OAI22_X1 port map( A1 => n13049, A2 => n11264, B1 => n11307, B2 => 
                           n11263, ZN => n1897);
   U387 : OAI22_X1 port map( A1 => n13320, A2 => n11264, B1 => n11308, B2 => 
                           n11262, ZN => n1896);
   U388 : OAI22_X1 port map( A1 => n13567, A2 => n11264, B1 => n11309, B2 => 
                           n11263, ZN => n1895);
   U389 : OAI22_X1 port map( A1 => n13050, A2 => n11264, B1 => n11310, B2 => 
                           n11262, ZN => n1894);
   U390 : OAI22_X1 port map( A1 => n13321, A2 => n11264, B1 => n11311, B2 => 
                           n11262, ZN => n1893);
   U391 : OAI22_X1 port map( A1 => n13051, A2 => n11264, B1 => n11312, B2 => 
                           n11262, ZN => n1892);
   U392 : OAI22_X1 port map( A1 => n13052, A2 => n11264, B1 => n11313, B2 => 
                           n11262, ZN => n1891);
   U393 : OAI22_X1 port map( A1 => n13568, A2 => n11264, B1 => n11314, B2 => 
                           n11262, ZN => n1890);
   U394 : OAI22_X1 port map( A1 => n13053, A2 => n11264, B1 => n11315, B2 => 
                           n11262, ZN => n1889);
   U395 : OAI22_X1 port map( A1 => n13809, A2 => n11264, B1 => n11317, B2 => 
                           n11262, ZN => n1888);
   U396 : OAI22_X1 port map( A1 => n13054, A2 => n11264, B1 => n11318, B2 => 
                           n11263, ZN => n1887);
   U397 : OAI22_X1 port map( A1 => n13322, A2 => n11264, B1 => n11319, B2 => 
                           n11263, ZN => n1886);
   U398 : OAI22_X1 port map( A1 => n13055, A2 => n11264, B1 => n11320, B2 => 
                           n11263, ZN => n1885);
   U399 : OAI22_X1 port map( A1 => n13323, A2 => n11264, B1 => n11321, B2 => 
                           n11263, ZN => n1884);
   U400 : OAI22_X1 port map( A1 => n13056, A2 => n11264, B1 => n11322, B2 => 
                           n11263, ZN => n1883);
   U401 : OAI22_X1 port map( A1 => n13569, A2 => n11264, B1 => n11323, B2 => 
                           n11263, ZN => n1882);
   U402 : OAI22_X1 port map( A1 => n13324, A2 => n11264, B1 => n11324, B2 => 
                           n11263, ZN => n1881);
   U403 : OAI22_X1 port map( A1 => n13570, A2 => n11264, B1 => n11325, B2 => 
                           n11263, ZN => n1880);
   U404 : OAI22_X1 port map( A1 => n13057, A2 => n11264, B1 => n11327, B2 => 
                           n11263, ZN => n1879);
   U405 : NAND2_X1 port map( A1 => n11354, A2 => n11284, ZN => n11265);
   U406 : CLKBUF_X1 port map( A => n11268, Z => n11266);
   U407 : CLKBUF_X1 port map( A => n11265, Z => n11267);
   U408 : OAI22_X1 port map( A1 => n13810, A2 => n11266, B1 => n11380, B2 => 
                           n11267, ZN => n1878);
   U409 : OAI22_X1 port map( A1 => n13058, A2 => n11268, B1 => n11295, B2 => 
                           n11265, ZN => n1877);
   U410 : OAI22_X1 port map( A1 => n13811, A2 => n11266, B1 => n11296, B2 => 
                           n11267, ZN => n1876);
   U411 : OAI22_X1 port map( A1 => n13812, A2 => n11268, B1 => n11297, B2 => 
                           n11265, ZN => n1875);
   U412 : OAI22_X1 port map( A1 => n13059, A2 => n11266, B1 => n11298, B2 => 
                           n11267, ZN => n1874);
   U413 : OAI22_X1 port map( A1 => n13813, A2 => n11268, B1 => n11299, B2 => 
                           n11265, ZN => n1873);
   U414 : OAI22_X1 port map( A1 => n13571, A2 => n11266, B1 => n11300, B2 => 
                           n11267, ZN => n1872);
   U415 : OAI22_X1 port map( A1 => n13060, A2 => n11268, B1 => n11301, B2 => 
                           n11265, ZN => n1871);
   U416 : OAI22_X1 port map( A1 => n13061, A2 => n11266, B1 => n11302, B2 => 
                           n11267, ZN => n1870);
   U417 : OAI22_X1 port map( A1 => n13325, A2 => n11268, B1 => n11303, B2 => 
                           n11265, ZN => n1869);
   U418 : OAI22_X1 port map( A1 => n13062, A2 => n11268, B1 => n11304, B2 => 
                           n11265, ZN => n1868);
   U419 : OAI22_X1 port map( A1 => n13572, A2 => n11268, B1 => n11305, B2 => 
                           n11267, ZN => n1867);
   U420 : OAI22_X1 port map( A1 => n13814, A2 => n11266, B1 => n11306, B2 => 
                           n11265, ZN => n1866);
   U421 : OAI22_X1 port map( A1 => n13063, A2 => n11266, B1 => n11307, B2 => 
                           n11267, ZN => n1865);
   U422 : OAI22_X1 port map( A1 => n13573, A2 => n11266, B1 => n11308, B2 => 
                           n11265, ZN => n1864);
   U423 : OAI22_X1 port map( A1 => n13064, A2 => n11266, B1 => n11309, B2 => 
                           n11267, ZN => n1863);
   U424 : OAI22_X1 port map( A1 => n13065, A2 => n11266, B1 => n11310, B2 => 
                           n11265, ZN => n1862);
   U425 : OAI22_X1 port map( A1 => n13066, A2 => n11266, B1 => n11311, B2 => 
                           n11265, ZN => n1861);
   U426 : OAI22_X1 port map( A1 => n13574, A2 => n11266, B1 => n11312, B2 => 
                           n11265, ZN => n1860);
   U427 : OAI22_X1 port map( A1 => n13067, A2 => n11266, B1 => n11313, B2 => 
                           n11265, ZN => n1859);
   U428 : OAI22_X1 port map( A1 => n13068, A2 => n11266, B1 => n11314, B2 => 
                           n11265, ZN => n1858);
   U429 : OAI22_X1 port map( A1 => n13815, A2 => n11266, B1 => n11315, B2 => 
                           n11265, ZN => n1857);
   U430 : OAI22_X1 port map( A1 => n13069, A2 => n11266, B1 => n11317, B2 => 
                           n11265, ZN => n1856);
   U431 : OAI22_X1 port map( A1 => n13816, A2 => n11266, B1 => n11318, B2 => 
                           n11267, ZN => n1855);
   U432 : OAI22_X1 port map( A1 => n13326, A2 => n11268, B1 => n11319, B2 => 
                           n11267, ZN => n1854);
   U433 : OAI22_X1 port map( A1 => n13817, A2 => n11268, B1 => n11320, B2 => 
                           n11267, ZN => n1853);
   U434 : OAI22_X1 port map( A1 => n13327, A2 => n11268, B1 => n11321, B2 => 
                           n11267, ZN => n1852);
   U435 : OAI22_X1 port map( A1 => n13328, A2 => n11268, B1 => n11322, B2 => 
                           n11267, ZN => n1851);
   U436 : OAI22_X1 port map( A1 => n13329, A2 => n11268, B1 => n11323, B2 => 
                           n11267, ZN => n1850);
   U437 : OAI22_X1 port map( A1 => n13818, A2 => n11268, B1 => n11324, B2 => 
                           n11267, ZN => n1849);
   U438 : OAI22_X1 port map( A1 => n13070, A2 => n11268, B1 => n11325, B2 => 
                           n11267, ZN => n1848);
   U439 : OAI22_X1 port map( A1 => n13819, A2 => n11268, B1 => n11327, B2 => 
                           n11267, ZN => n1847);
   U440 : NAND2_X1 port map( A1 => n11358, A2 => n11284, ZN => n11269);
   U441 : CLKBUF_X1 port map( A => n11269, Z => n11270);
   U442 : OAI22_X1 port map( A1 => n13330, A2 => n11271, B1 => n11380, B2 => 
                           n11270, ZN => n1846);
   U443 : OAI22_X1 port map( A1 => n13575, A2 => n11271, B1 => n11295, B2 => 
                           n11269, ZN => n1845);
   U444 : OAI22_X1 port map( A1 => n13576, A2 => n11271, B1 => n11296, B2 => 
                           n11270, ZN => n1844);
   U445 : OAI22_X1 port map( A1 => n13071, A2 => n11271, B1 => n11297, B2 => 
                           n11269, ZN => n1843);
   U446 : OAI22_X1 port map( A1 => n13331, A2 => n11271, B1 => n11298, B2 => 
                           n11270, ZN => n1842);
   U447 : OAI22_X1 port map( A1 => n13072, A2 => n11271, B1 => n11299, B2 => 
                           n11269, ZN => n1841);
   U448 : OAI22_X1 port map( A1 => n13332, A2 => n11271, B1 => n11300, B2 => 
                           n11270, ZN => n1840);
   U449 : OAI22_X1 port map( A1 => n13577, A2 => n11271, B1 => n11301, B2 => 
                           n11269, ZN => n1839);
   U450 : OAI22_X1 port map( A1 => n13333, A2 => n11271, B1 => n11302, B2 => 
                           n11270, ZN => n1838);
   U451 : OAI22_X1 port map( A1 => n13073, A2 => n11271, B1 => n11303, B2 => 
                           n11269, ZN => n1837);
   U452 : OAI22_X1 port map( A1 => n13334, A2 => n11271, B1 => n11304, B2 => 
                           n11269, ZN => n1836);
   U453 : OAI22_X1 port map( A1 => n13335, A2 => n11271, B1 => n11305, B2 => 
                           n11270, ZN => n1835);
   U454 : OAI22_X1 port map( A1 => n13336, A2 => n11271, B1 => n11306, B2 => 
                           n11269, ZN => n1834);
   U455 : OAI22_X1 port map( A1 => n13074, A2 => n11271, B1 => n11307, B2 => 
                           n11270, ZN => n1833);
   U456 : OAI22_X1 port map( A1 => n13820, A2 => n11271, B1 => n11308, B2 => 
                           n11269, ZN => n1832);
   U457 : OAI22_X1 port map( A1 => n13821, A2 => n11271, B1 => n11309, B2 => 
                           n11270, ZN => n1831);
   U458 : OAI22_X1 port map( A1 => n13822, A2 => n11271, B1 => n11310, B2 => 
                           n11269, ZN => n1830);
   U459 : OAI22_X1 port map( A1 => n13823, A2 => n11271, B1 => n11311, B2 => 
                           n11269, ZN => n1829);
   U460 : OAI22_X1 port map( A1 => n13578, A2 => n11271, B1 => n11312, B2 => 
                           n11269, ZN => n1828);
   U461 : OAI22_X1 port map( A1 => n13824, A2 => n11271, B1 => n11313, B2 => 
                           n11269, ZN => n1827);
   U462 : OAI22_X1 port map( A1 => n13337, A2 => n11271, B1 => n11314, B2 => 
                           n11269, ZN => n1826);
   U463 : OAI22_X1 port map( A1 => n13338, A2 => n11271, B1 => n11315, B2 => 
                           n11269, ZN => n1825);
   U464 : OAI22_X1 port map( A1 => n13825, A2 => n11271, B1 => n11317, B2 => 
                           n11269, ZN => n1824);
   U465 : OAI22_X1 port map( A1 => n13339, A2 => n11271, B1 => n11318, B2 => 
                           n11270, ZN => n1823);
   U466 : OAI22_X1 port map( A1 => n13075, A2 => n11271, B1 => n11319, B2 => 
                           n11270, ZN => n1822);
   U467 : OAI22_X1 port map( A1 => n13340, A2 => n11271, B1 => n11320, B2 => 
                           n11270, ZN => n1821);
   U468 : OAI22_X1 port map( A1 => n13579, A2 => n11271, B1 => n11321, B2 => 
                           n11270, ZN => n1820);
   U469 : OAI22_X1 port map( A1 => n13826, A2 => n11271, B1 => n11322, B2 => 
                           n11270, ZN => n1819);
   U470 : OAI22_X1 port map( A1 => n13580, A2 => n11271, B1 => n11323, B2 => 
                           n11270, ZN => n1818);
   U471 : OAI22_X1 port map( A1 => n13341, A2 => n11271, B1 => n11324, B2 => 
                           n11270, ZN => n1817);
   U472 : OAI22_X1 port map( A1 => n13827, A2 => n11271, B1 => n11325, B2 => 
                           n11270, ZN => n1816);
   U473 : OAI22_X1 port map( A1 => n13076, A2 => n11271, B1 => n11327, B2 => 
                           n11270, ZN => n1815);
   U474 : NAND2_X1 port map( A1 => n11362, A2 => n11284, ZN => n11272);
   U475 : CLKBUF_X1 port map( A => n11272, Z => n11273);
   U476 : OAI22_X1 port map( A1 => n13077, A2 => n11274, B1 => n11380, B2 => 
                           n11273, ZN => n1814);
   U477 : CLKBUF_X1 port map( A => n11295, Z => n11381);
   U478 : OAI22_X1 port map( A1 => n13342, A2 => n11274, B1 => n11381, B2 => 
                           n11272, ZN => n1813);
   U479 : CLKBUF_X1 port map( A => n11296, Z => n11382);
   U480 : OAI22_X1 port map( A1 => n13343, A2 => n11274, B1 => n11382, B2 => 
                           n11273, ZN => n1812);
   U481 : CLKBUF_X1 port map( A => n11297, Z => n11383);
   U482 : OAI22_X1 port map( A1 => n13344, A2 => n11274, B1 => n11383, B2 => 
                           n11272, ZN => n1811);
   U483 : CLKBUF_X1 port map( A => n11298, Z => n11384);
   U484 : OAI22_X1 port map( A1 => n13345, A2 => n11274, B1 => n11384, B2 => 
                           n11273, ZN => n1810);
   U485 : CLKBUF_X1 port map( A => n11299, Z => n11385);
   U486 : OAI22_X1 port map( A1 => n13346, A2 => n11274, B1 => n11385, B2 => 
                           n11272, ZN => n1809);
   U487 : CLKBUF_X1 port map( A => n11300, Z => n11386);
   U488 : OAI22_X1 port map( A1 => n13078, A2 => n11274, B1 => n11386, B2 => 
                           n11273, ZN => n1808);
   U489 : OAI22_X1 port map( A1 => n13079, A2 => n11274, B1 => n11387, B2 => 
                           n11272, ZN => n1807);
   U490 : CLKBUF_X1 port map( A => n11302, Z => n11388);
   U491 : OAI22_X1 port map( A1 => n13080, A2 => n11274, B1 => n11388, B2 => 
                           n11273, ZN => n1806);
   U492 : CLKBUF_X1 port map( A => n11303, Z => n11389);
   U493 : OAI22_X1 port map( A1 => n13081, A2 => n11274, B1 => n11389, B2 => 
                           n11272, ZN => n1805);
   U494 : CLKBUF_X1 port map( A => n11304, Z => n11390);
   U495 : OAI22_X1 port map( A1 => n13082, A2 => n11274, B1 => n11390, B2 => 
                           n11272, ZN => n1804);
   U496 : CLKBUF_X1 port map( A => n11305, Z => n11391);
   U497 : OAI22_X1 port map( A1 => n13347, A2 => n11274, B1 => n11391, B2 => 
                           n11273, ZN => n1803);
   U498 : CLKBUF_X1 port map( A => n11306, Z => n11392);
   U499 : OAI22_X1 port map( A1 => n13348, A2 => n11274, B1 => n11392, B2 => 
                           n11272, ZN => n1802);
   U500 : CLKBUF_X1 port map( A => n11307, Z => n11393);
   U501 : OAI22_X1 port map( A1 => n13349, A2 => n11274, B1 => n11393, B2 => 
                           n11273, ZN => n1801);
   U502 : CLKBUF_X1 port map( A => n11308, Z => n11394);
   U503 : OAI22_X1 port map( A1 => n13350, A2 => n11274, B1 => n11394, B2 => 
                           n11272, ZN => n1800);
   U504 : CLKBUF_X1 port map( A => n11309, Z => n11395);
   U505 : OAI22_X1 port map( A1 => n13083, A2 => n11274, B1 => n11395, B2 => 
                           n11273, ZN => n1799);
   U506 : CLKBUF_X1 port map( A => n11310, Z => n11396);
   U507 : OAI22_X1 port map( A1 => n13084, A2 => n11274, B1 => n11396, B2 => 
                           n11272, ZN => n1798);
   U508 : CLKBUF_X1 port map( A => n11311, Z => n11397);
   U509 : OAI22_X1 port map( A1 => n13085, A2 => n11274, B1 => n11397, B2 => 
                           n11272, ZN => n1797);
   U510 : CLKBUF_X1 port map( A => n11312, Z => n11398);
   U511 : OAI22_X1 port map( A1 => n13086, A2 => n11274, B1 => n11398, B2 => 
                           n11272, ZN => n1796);
   U512 : CLKBUF_X1 port map( A => n11313, Z => n11399);
   U513 : OAI22_X1 port map( A1 => n13087, A2 => n11274, B1 => n11399, B2 => 
                           n11272, ZN => n1795);
   U514 : CLKBUF_X1 port map( A => n11314, Z => n11400);
   U515 : OAI22_X1 port map( A1 => n13088, A2 => n11274, B1 => n11400, B2 => 
                           n11272, ZN => n1794);
   U516 : CLKBUF_X1 port map( A => n11315, Z => n11401);
   U517 : OAI22_X1 port map( A1 => n13351, A2 => n11274, B1 => n11401, B2 => 
                           n11272, ZN => n1793);
   U518 : OAI22_X1 port map( A1 => n13089, A2 => n11274, B1 => n11403, B2 => 
                           n11272, ZN => n1792);
   U519 : CLKBUF_X1 port map( A => n11318, Z => n11404);
   U520 : OAI22_X1 port map( A1 => n13352, A2 => n11274, B1 => n11404, B2 => 
                           n11273, ZN => n1791);
   U521 : CLKBUF_X1 port map( A => n11319, Z => n11405);
   U522 : OAI22_X1 port map( A1 => n13090, A2 => n11274, B1 => n11405, B2 => 
                           n11273, ZN => n1790);
   U523 : CLKBUF_X1 port map( A => n11320, Z => n11406);
   U524 : OAI22_X1 port map( A1 => n13353, A2 => n11274, B1 => n11406, B2 => 
                           n11273, ZN => n1789);
   U525 : CLKBUF_X1 port map( A => n11321, Z => n11407);
   U526 : OAI22_X1 port map( A1 => n13091, A2 => n11274, B1 => n11407, B2 => 
                           n11273, ZN => n1788);
   U527 : CLKBUF_X1 port map( A => n11322, Z => n11408);
   U528 : OAI22_X1 port map( A1 => n13354, A2 => n11274, B1 => n11408, B2 => 
                           n11273, ZN => n1787);
   U529 : CLKBUF_X1 port map( A => n11323, Z => n11409);
   U530 : OAI22_X1 port map( A1 => n13092, A2 => n11274, B1 => n11409, B2 => 
                           n11273, ZN => n1786);
   U531 : CLKBUF_X1 port map( A => n11324, Z => n11410);
   U532 : OAI22_X1 port map( A1 => n13093, A2 => n11274, B1 => n11410, B2 => 
                           n11273, ZN => n1785);
   U533 : CLKBUF_X1 port map( A => n11325, Z => n11411);
   U534 : OAI22_X1 port map( A1 => n13355, A2 => n11274, B1 => n11411, B2 => 
                           n11273, ZN => n1784);
   U535 : CLKBUF_X1 port map( A => n11327, Z => n11413);
   U536 : OAI22_X1 port map( A1 => n13094, A2 => n11274, B1 => n11413, B2 => 
                           n11273, ZN => n1783);
   U537 : NAND2_X1 port map( A1 => n11366, A2 => n11284, ZN => n11275);
   U538 : CLKBUF_X1 port map( A => n11275, Z => n11276);
   U539 : OAI22_X1 port map( A1 => n13828, A2 => n11277, B1 => n11343, B2 => 
                           n11276, ZN => n1782);
   U540 : OAI22_X1 port map( A1 => n13581, A2 => n11277, B1 => n11295, B2 => 
                           n11275, ZN => n1781);
   U541 : OAI22_X1 port map( A1 => n13095, A2 => n11277, B1 => n11296, B2 => 
                           n11276, ZN => n1780);
   U542 : OAI22_X1 port map( A1 => n13829, A2 => n11277, B1 => n11297, B2 => 
                           n11275, ZN => n1779);
   U543 : OAI22_X1 port map( A1 => n13830, A2 => n11277, B1 => n11298, B2 => 
                           n11276, ZN => n1778);
   U544 : OAI22_X1 port map( A1 => n13582, A2 => n11277, B1 => n11299, B2 => 
                           n11275, ZN => n1777);
   U545 : OAI22_X1 port map( A1 => n13356, A2 => n11277, B1 => n11300, B2 => 
                           n11276, ZN => n1776);
   U546 : OAI22_X1 port map( A1 => n13831, A2 => n11277, B1 => n11301, B2 => 
                           n11275, ZN => n1775);
   U547 : OAI22_X1 port map( A1 => n13583, A2 => n11277, B1 => n11302, B2 => 
                           n11276, ZN => n1774);
   U548 : OAI22_X1 port map( A1 => n13832, A2 => n11277, B1 => n11303, B2 => 
                           n11275, ZN => n1773);
   U549 : OAI22_X1 port map( A1 => n13584, A2 => n11277, B1 => n11304, B2 => 
                           n11275, ZN => n1772);
   U550 : OAI22_X1 port map( A1 => n13585, A2 => n11277, B1 => n11305, B2 => 
                           n11276, ZN => n1771);
   U551 : OAI22_X1 port map( A1 => n13096, A2 => n11277, B1 => n11306, B2 => 
                           n11275, ZN => n1770);
   U552 : OAI22_X1 port map( A1 => n13833, A2 => n11277, B1 => n11307, B2 => 
                           n11276, ZN => n1769);
   U553 : OAI22_X1 port map( A1 => n13097, A2 => n11277, B1 => n11308, B2 => 
                           n11275, ZN => n1768);
   U554 : OAI22_X1 port map( A1 => n13357, A2 => n11277, B1 => n11309, B2 => 
                           n11276, ZN => n1767);
   U555 : OAI22_X1 port map( A1 => n13586, A2 => n11277, B1 => n11310, B2 => 
                           n11275, ZN => n1766);
   U556 : OAI22_X1 port map( A1 => n13358, A2 => n11277, B1 => n11311, B2 => 
                           n11275, ZN => n1765);
   U557 : OAI22_X1 port map( A1 => n13359, A2 => n11277, B1 => n11312, B2 => 
                           n11275, ZN => n1764);
   U558 : OAI22_X1 port map( A1 => n13834, A2 => n11277, B1 => n11313, B2 => 
                           n11275, ZN => n1763);
   U559 : OAI22_X1 port map( A1 => n13835, A2 => n11277, B1 => n11314, B2 => 
                           n11275, ZN => n1762);
   U560 : OAI22_X1 port map( A1 => n13836, A2 => n11277, B1 => n11315, B2 => 
                           n11275, ZN => n1761);
   U561 : OAI22_X1 port map( A1 => n13837, A2 => n11277, B1 => n11317, B2 => 
                           n11275, ZN => n1760);
   U562 : OAI22_X1 port map( A1 => n13587, A2 => n11277, B1 => n11318, B2 => 
                           n11276, ZN => n1759);
   U563 : OAI22_X1 port map( A1 => n13588, A2 => n11277, B1 => n11319, B2 => 
                           n11276, ZN => n1758);
   U564 : OAI22_X1 port map( A1 => n13589, A2 => n11277, B1 => n11320, B2 => 
                           n11276, ZN => n1757);
   U565 : OAI22_X1 port map( A1 => n13838, A2 => n11277, B1 => n11321, B2 => 
                           n11276, ZN => n1756);
   U566 : OAI22_X1 port map( A1 => n13590, A2 => n11277, B1 => n11322, B2 => 
                           n11276, ZN => n1755);
   U567 : OAI22_X1 port map( A1 => n13098, A2 => n11277, B1 => n11323, B2 => 
                           n11276, ZN => n1754);
   U568 : OAI22_X1 port map( A1 => n13591, A2 => n11277, B1 => n11324, B2 => 
                           n11276, ZN => n1753);
   U569 : OAI22_X1 port map( A1 => n13592, A2 => n11277, B1 => n11325, B2 => 
                           n11276, ZN => n1752);
   U570 : OAI22_X1 port map( A1 => n13839, A2 => n11277, B1 => n11327, B2 => 
                           n11276, ZN => n1751);
   U571 : NAND2_X1 port map( A1 => n11370, A2 => n11284, ZN => n11278);
   U572 : OAI22_X1 port map( A1 => n13593, A2 => n11280, B1 => n11343, B2 => 
                           n11279, ZN => n1750);
   U573 : OAI22_X1 port map( A1 => n13594, A2 => n11280, B1 => n11381, B2 => 
                           n11278, ZN => n1749);
   U574 : OAI22_X1 port map( A1 => n13840, A2 => n11280, B1 => n11382, B2 => 
                           n11279, ZN => n1748);
   U575 : OAI22_X1 port map( A1 => n13595, A2 => n11280, B1 => n11383, B2 => 
                           n11278, ZN => n1747);
   U576 : OAI22_X1 port map( A1 => n13596, A2 => n11280, B1 => n11384, B2 => 
                           n11279, ZN => n1746);
   U577 : OAI22_X1 port map( A1 => n13597, A2 => n11280, B1 => n11385, B2 => 
                           n11278, ZN => n1745);
   U578 : OAI22_X1 port map( A1 => n13841, A2 => n11280, B1 => n11386, B2 => 
                           n11279, ZN => n1744);
   U579 : OAI22_X1 port map( A1 => n13842, A2 => n11280, B1 => n11387, B2 => 
                           n11278, ZN => n1743);
   U580 : OAI22_X1 port map( A1 => n13598, A2 => n11280, B1 => n11388, B2 => 
                           n11279, ZN => n1742);
   U581 : OAI22_X1 port map( A1 => n13843, A2 => n11280, B1 => n11389, B2 => 
                           n11278, ZN => n1741);
   U582 : OAI22_X1 port map( A1 => n13844, A2 => n11280, B1 => n11390, B2 => 
                           n11278, ZN => n1740);
   U583 : OAI22_X1 port map( A1 => n13845, A2 => n11280, B1 => n11391, B2 => 
                           n11279, ZN => n1739);
   U584 : OAI22_X1 port map( A1 => n13599, A2 => n11280, B1 => n11392, B2 => 
                           n11278, ZN => n1738);
   U585 : OAI22_X1 port map( A1 => n13846, A2 => n11280, B1 => n11393, B2 => 
                           n11279, ZN => n1737);
   U586 : OAI22_X1 port map( A1 => n13600, A2 => n11280, B1 => n11394, B2 => 
                           n11278, ZN => n1736);
   U587 : OAI22_X1 port map( A1 => n13601, A2 => n11280, B1 => n11395, B2 => 
                           n11279, ZN => n1735);
   U588 : OAI22_X1 port map( A1 => n13847, A2 => n11280, B1 => n11396, B2 => 
                           n11278, ZN => n1734);
   U589 : OAI22_X1 port map( A1 => n13602, A2 => n11280, B1 => n11397, B2 => 
                           n11278, ZN => n1733);
   U590 : OAI22_X1 port map( A1 => n13848, A2 => n11280, B1 => n11398, B2 => 
                           n11278, ZN => n1732);
   U591 : OAI22_X1 port map( A1 => n13603, A2 => n11280, B1 => n11399, B2 => 
                           n11278, ZN => n1731);
   U592 : OAI22_X1 port map( A1 => n13849, A2 => n11280, B1 => n11400, B2 => 
                           n11278, ZN => n1730);
   U593 : OAI22_X1 port map( A1 => n13604, A2 => n11280, B1 => n11401, B2 => 
                           n11278, ZN => n1729);
   U594 : OAI22_X1 port map( A1 => n13605, A2 => n11280, B1 => n11403, B2 => 
                           n11278, ZN => n1728);
   U595 : OAI22_X1 port map( A1 => n13606, A2 => n11280, B1 => n11404, B2 => 
                           n11279, ZN => n1727);
   U596 : OAI22_X1 port map( A1 => n13607, A2 => n11280, B1 => n11405, B2 => 
                           n11279, ZN => n1726);
   U597 : OAI22_X1 port map( A1 => n13608, A2 => n11280, B1 => n11406, B2 => 
                           n11279, ZN => n1725);
   U598 : OAI22_X1 port map( A1 => n13609, A2 => n11280, B1 => n11407, B2 => 
                           n11279, ZN => n1724);
   U599 : OAI22_X1 port map( A1 => n13850, A2 => n11280, B1 => n11408, B2 => 
                           n11279, ZN => n1723);
   U600 : OAI22_X1 port map( A1 => n13851, A2 => n11280, B1 => n11409, B2 => 
                           n11279, ZN => n1722);
   U601 : OAI22_X1 port map( A1 => n13852, A2 => n11280, B1 => n11410, B2 => 
                           n11279, ZN => n1721);
   U602 : OAI22_X1 port map( A1 => n13610, A2 => n11280, B1 => n11411, B2 => 
                           n11279, ZN => n1720);
   U603 : OAI22_X1 port map( A1 => n13853, A2 => n11280, B1 => n11413, B2 => 
                           n11279, ZN => n1719);
   U604 : NAND2_X1 port map( A1 => n11374, A2 => n11284, ZN => n11281);
   U605 : CLKBUF_X1 port map( A => n11281, Z => n11282);
   U606 : OAI22_X1 port map( A1 => n13360, A2 => n11283, B1 => n11343, B2 => 
                           n11282, ZN => n1718);
   U607 : OAI22_X1 port map( A1 => n13854, A2 => n11283, B1 => n11295, B2 => 
                           n11281, ZN => n1717);
   U608 : OAI22_X1 port map( A1 => n13611, A2 => n11283, B1 => n11296, B2 => 
                           n11282, ZN => n1716);
   U609 : OAI22_X1 port map( A1 => n13612, A2 => n11283, B1 => n11297, B2 => 
                           n11281, ZN => n1715);
   U610 : OAI22_X1 port map( A1 => n13613, A2 => n11283, B1 => n11298, B2 => 
                           n11282, ZN => n1714);
   U611 : OAI22_X1 port map( A1 => n13855, A2 => n11283, B1 => n11299, B2 => 
                           n11281, ZN => n1713);
   U612 : OAI22_X1 port map( A1 => n13614, A2 => n11283, B1 => n11300, B2 => 
                           n11282, ZN => n1712);
   U613 : OAI22_X1 port map( A1 => n13615, A2 => n11283, B1 => n11301, B2 => 
                           n11281, ZN => n1711);
   U614 : OAI22_X1 port map( A1 => n13856, A2 => n11283, B1 => n11302, B2 => 
                           n11282, ZN => n1710);
   U615 : OAI22_X1 port map( A1 => n13616, A2 => n11283, B1 => n11303, B2 => 
                           n11281, ZN => n1709);
   U616 : OAI22_X1 port map( A1 => n13617, A2 => n11283, B1 => n11304, B2 => 
                           n11281, ZN => n1708);
   U617 : OAI22_X1 port map( A1 => n13618, A2 => n11283, B1 => n11305, B2 => 
                           n11282, ZN => n1707);
   U618 : OAI22_X1 port map( A1 => n13857, A2 => n11283, B1 => n11306, B2 => 
                           n11281, ZN => n1706);
   U619 : OAI22_X1 port map( A1 => n13619, A2 => n11283, B1 => n11307, B2 => 
                           n11282, ZN => n1705);
   U620 : OAI22_X1 port map( A1 => n13620, A2 => n11283, B1 => n11308, B2 => 
                           n11281, ZN => n1704);
   U621 : OAI22_X1 port map( A1 => n13858, A2 => n11283, B1 => n11309, B2 => 
                           n11282, ZN => n1703);
   U622 : OAI22_X1 port map( A1 => n13859, A2 => n11283, B1 => n11310, B2 => 
                           n11281, ZN => n1702);
   U623 : OAI22_X1 port map( A1 => n13860, A2 => n11283, B1 => n11311, B2 => 
                           n11281, ZN => n1701);
   U624 : OAI22_X1 port map( A1 => n13861, A2 => n11283, B1 => n11312, B2 => 
                           n11281, ZN => n1700);
   U625 : OAI22_X1 port map( A1 => n13862, A2 => n11283, B1 => n11313, B2 => 
                           n11281, ZN => n1699);
   U626 : OAI22_X1 port map( A1 => n13863, A2 => n11283, B1 => n11314, B2 => 
                           n11281, ZN => n1698);
   U627 : OAI22_X1 port map( A1 => n13621, A2 => n11283, B1 => n11315, B2 => 
                           n11281, ZN => n1697);
   U628 : OAI22_X1 port map( A1 => n13099, A2 => n11283, B1 => n11317, B2 => 
                           n11281, ZN => n1696);
   U629 : OAI22_X1 port map( A1 => n13864, A2 => n11283, B1 => n11318, B2 => 
                           n11282, ZN => n1695);
   U630 : OAI22_X1 port map( A1 => n13865, A2 => n11283, B1 => n11319, B2 => 
                           n11282, ZN => n1694);
   U631 : OAI22_X1 port map( A1 => n13622, A2 => n11283, B1 => n11320, B2 => 
                           n11282, ZN => n1693);
   U632 : OAI22_X1 port map( A1 => n13866, A2 => n11283, B1 => n11321, B2 => 
                           n11282, ZN => n1692);
   U633 : OAI22_X1 port map( A1 => n13623, A2 => n11283, B1 => n11322, B2 => 
                           n11282, ZN => n1691);
   U634 : OAI22_X1 port map( A1 => n13867, A2 => n11283, B1 => n11323, B2 => 
                           n11282, ZN => n1690);
   U635 : OAI22_X1 port map( A1 => n13624, A2 => n11283, B1 => n11324, B2 => 
                           n11282, ZN => n1689);
   U636 : OAI22_X1 port map( A1 => n13361, A2 => n11283, B1 => n11325, B2 => 
                           n11282, ZN => n1688);
   U637 : OAI22_X1 port map( A1 => n13625, A2 => n11283, B1 => n11327, B2 => 
                           n11282, ZN => n1687);
   U638 : NAND2_X1 port map( A1 => n11379, A2 => n11284, ZN => n11285);
   U639 : CLKBUF_X1 port map( A => n11285, Z => n11286);
   U640 : OAI22_X1 port map( A1 => n13100, A2 => n11287, B1 => n11343, B2 => 
                           n11286, ZN => n1686);
   U641 : OAI22_X1 port map( A1 => n13362, A2 => n11287, B1 => n11381, B2 => 
                           n11285, ZN => n1685);
   U642 : OAI22_X1 port map( A1 => n13101, A2 => n11287, B1 => n11382, B2 => 
                           n11286, ZN => n1684);
   U643 : OAI22_X1 port map( A1 => n13363, A2 => n11287, B1 => n11383, B2 => 
                           n11285, ZN => n1683);
   U644 : OAI22_X1 port map( A1 => n13102, A2 => n11287, B1 => n11384, B2 => 
                           n11286, ZN => n1682);
   U645 : OAI22_X1 port map( A1 => n13364, A2 => n11287, B1 => n11385, B2 => 
                           n11285, ZN => n1681);
   U646 : OAI22_X1 port map( A1 => n13365, A2 => n11287, B1 => n11386, B2 => 
                           n11286, ZN => n1680);
   U647 : OAI22_X1 port map( A1 => n13366, A2 => n11287, B1 => n11387, B2 => 
                           n11285, ZN => n1679);
   U648 : OAI22_X1 port map( A1 => n13367, A2 => n11287, B1 => n11388, B2 => 
                           n11286, ZN => n1678);
   U649 : OAI22_X1 port map( A1 => n13368, A2 => n11287, B1 => n11389, B2 => 
                           n11285, ZN => n1677);
   U650 : OAI22_X1 port map( A1 => n13868, A2 => n11287, B1 => n11390, B2 => 
                           n11285, ZN => n1676);
   U651 : OAI22_X1 port map( A1 => n13103, A2 => n11287, B1 => n11391, B2 => 
                           n11286, ZN => n1675);
   U652 : OAI22_X1 port map( A1 => n13626, A2 => n11287, B1 => n11392, B2 => 
                           n11285, ZN => n1674);
   U653 : OAI22_X1 port map( A1 => n13869, A2 => n11287, B1 => n11393, B2 => 
                           n11286, ZN => n1673);
   U654 : OAI22_X1 port map( A1 => n13369, A2 => n11287, B1 => n11394, B2 => 
                           n11285, ZN => n1672);
   U655 : OAI22_X1 port map( A1 => n13370, A2 => n11287, B1 => n11395, B2 => 
                           n11286, ZN => n1671);
   U656 : OAI22_X1 port map( A1 => n13371, A2 => n11287, B1 => n11396, B2 => 
                           n11285, ZN => n1670);
   U657 : OAI22_X1 port map( A1 => n13627, A2 => n11287, B1 => n11397, B2 => 
                           n11285, ZN => n1669);
   U658 : OAI22_X1 port map( A1 => n13372, A2 => n11287, B1 => n11398, B2 => 
                           n11285, ZN => n1668);
   U659 : OAI22_X1 port map( A1 => n13373, A2 => n11287, B1 => n11399, B2 => 
                           n11285, ZN => n1667);
   U660 : OAI22_X1 port map( A1 => n13104, A2 => n11287, B1 => n11400, B2 => 
                           n11285, ZN => n1666);
   U661 : OAI22_X1 port map( A1 => n13105, A2 => n11287, B1 => n11401, B2 => 
                           n11285, ZN => n1665);
   U662 : OAI22_X1 port map( A1 => n13374, A2 => n11287, B1 => n11403, B2 => 
                           n11285, ZN => n1664);
   U663 : OAI22_X1 port map( A1 => n13106, A2 => n11287, B1 => n11404, B2 => 
                           n11286, ZN => n1663);
   U664 : OAI22_X1 port map( A1 => n13870, A2 => n11287, B1 => n11405, B2 => 
                           n11286, ZN => n1662);
   U665 : OAI22_X1 port map( A1 => n13375, A2 => n11287, B1 => n11406, B2 => 
                           n11286, ZN => n1661);
   U666 : OAI22_X1 port map( A1 => n13107, A2 => n11287, B1 => n11407, B2 => 
                           n11286, ZN => n1660);
   U667 : OAI22_X1 port map( A1 => n13108, A2 => n11287, B1 => n11408, B2 => 
                           n11286, ZN => n1659);
   U668 : OAI22_X1 port map( A1 => n13376, A2 => n11287, B1 => n11409, B2 => 
                           n11286, ZN => n1658);
   U669 : OAI22_X1 port map( A1 => n13109, A2 => n11287, B1 => n11410, B2 => 
                           n11286, ZN => n1657);
   U670 : OAI22_X1 port map( A1 => n13377, A2 => n11287, B1 => n11411, B2 => 
                           n11286, ZN => n1656);
   U671 : OAI22_X1 port map( A1 => n13378, A2 => n11287, B1 => n11413, B2 => 
                           n11286, ZN => n1655);
   U672 : NOR2_X1 port map( A1 => n11348, A2 => n11288, ZN => n11342);
   U673 : NAND2_X1 port map( A1 => n11349, A2 => n11342, ZN => n11289);
   U674 : CLKBUF_X1 port map( A => n11289, Z => n11290);
   U675 : OAI22_X1 port map( A1 => n12979, A2 => n11291, B1 => n11343, B2 => 
                           n11290, ZN => n1654);
   U676 : OAI22_X1 port map( A1 => n13110, A2 => n11291, B1 => n11295, B2 => 
                           n11289, ZN => n1653);
   U677 : OAI22_X1 port map( A1 => n13871, A2 => n11291, B1 => n11296, B2 => 
                           n11290, ZN => n1652);
   U678 : OAI22_X1 port map( A1 => n13628, A2 => n11291, B1 => n11297, B2 => 
                           n11289, ZN => n1651);
   U679 : OAI22_X1 port map( A1 => n13872, A2 => n11291, B1 => n11298, B2 => 
                           n11290, ZN => n1650);
   U680 : OAI22_X1 port map( A1 => n13379, A2 => n11291, B1 => n11299, B2 => 
                           n11289, ZN => n1649);
   U681 : OAI22_X1 port map( A1 => n13380, A2 => n11291, B1 => n11300, B2 => 
                           n11290, ZN => n1648);
   U682 : OAI22_X1 port map( A1 => n13629, A2 => n11291, B1 => n11301, B2 => 
                           n11289, ZN => n1647);
   U683 : OAI22_X1 port map( A1 => n13381, A2 => n11291, B1 => n11302, B2 => 
                           n11290, ZN => n1646);
   U684 : OAI22_X1 port map( A1 => n13873, A2 => n11291, B1 => n11303, B2 => 
                           n11289, ZN => n1645);
   U685 : OAI22_X1 port map( A1 => n13630, A2 => n11291, B1 => n11304, B2 => 
                           n11289, ZN => n1644);
   U686 : OAI22_X1 port map( A1 => n13631, A2 => n11291, B1 => n11305, B2 => 
                           n11290, ZN => n1643);
   U687 : OAI22_X1 port map( A1 => n13111, A2 => n11291, B1 => n11306, B2 => 
                           n11289, ZN => n1642);
   U688 : OAI22_X1 port map( A1 => n13382, A2 => n11291, B1 => n11307, B2 => 
                           n11290, ZN => n1641);
   U689 : OAI22_X1 port map( A1 => n13874, A2 => n11291, B1 => n11308, B2 => 
                           n11289, ZN => n1640);
   U690 : OAI22_X1 port map( A1 => n13383, A2 => n11291, B1 => n11309, B2 => 
                           n11290, ZN => n1639);
   U691 : OAI22_X1 port map( A1 => n13875, A2 => n11291, B1 => n11310, B2 => 
                           n11289, ZN => n1638);
   U692 : OAI22_X1 port map( A1 => n13876, A2 => n11291, B1 => n11311, B2 => 
                           n11289, ZN => n1637);
   U693 : OAI22_X1 port map( A1 => n13384, A2 => n11291, B1 => n11312, B2 => 
                           n11289, ZN => n1636);
   U694 : OAI22_X1 port map( A1 => n13877, A2 => n11291, B1 => n11313, B2 => 
                           n11289, ZN => n1635);
   U695 : OAI22_X1 port map( A1 => n13878, A2 => n11291, B1 => n11314, B2 => 
                           n11289, ZN => n1634);
   U696 : OAI22_X1 port map( A1 => n13879, A2 => n11291, B1 => n11315, B2 => 
                           n11289, ZN => n1633);
   U697 : OAI22_X1 port map( A1 => n13112, A2 => n11291, B1 => n11317, B2 => 
                           n11289, ZN => n1632);
   U698 : OAI22_X1 port map( A1 => n13880, A2 => n11291, B1 => n11318, B2 => 
                           n11290, ZN => n1631);
   U699 : OAI22_X1 port map( A1 => n13385, A2 => n11291, B1 => n11319, B2 => 
                           n11290, ZN => n1630);
   U700 : OAI22_X1 port map( A1 => n13386, A2 => n11291, B1 => n11320, B2 => 
                           n11290, ZN => n1629);
   U701 : OAI22_X1 port map( A1 => n13632, A2 => n11291, B1 => n11321, B2 => 
                           n11290, ZN => n1628);
   U702 : OAI22_X1 port map( A1 => n13113, A2 => n11291, B1 => n11322, B2 => 
                           n11290, ZN => n1627);
   U703 : OAI22_X1 port map( A1 => n13114, A2 => n11291, B1 => n11323, B2 => 
                           n11290, ZN => n1626);
   U704 : OAI22_X1 port map( A1 => n13115, A2 => n11291, B1 => n11324, B2 => 
                           n11290, ZN => n1625);
   U705 : OAI22_X1 port map( A1 => n13881, A2 => n11291, B1 => n11325, B2 => 
                           n11290, ZN => n1624);
   U706 : OAI22_X1 port map( A1 => n13882, A2 => n11291, B1 => n11327, B2 => 
                           n11290, ZN => n1623);
   U707 : NAND2_X1 port map( A1 => n11354, A2 => n11342, ZN => n11292);
   U708 : CLKBUF_X1 port map( A => n11292, Z => n11293);
   U709 : OAI22_X1 port map( A1 => n13242, A2 => n11294, B1 => n11343, B2 => 
                           n11293, ZN => n1622);
   U710 : OAI22_X1 port map( A1 => n13883, A2 => n11294, B1 => n11381, B2 => 
                           n11292, ZN => n1621);
   U711 : OAI22_X1 port map( A1 => n13116, A2 => n11294, B1 => n11382, B2 => 
                           n11293, ZN => n1620);
   U712 : OAI22_X1 port map( A1 => n13884, A2 => n11294, B1 => n11383, B2 => 
                           n11292, ZN => n1619);
   U713 : OAI22_X1 port map( A1 => n13633, A2 => n11294, B1 => n11384, B2 => 
                           n11293, ZN => n1618);
   U714 : OAI22_X1 port map( A1 => n13885, A2 => n11294, B1 => n11385, B2 => 
                           n11292, ZN => n1617);
   U715 : OAI22_X1 port map( A1 => n13634, A2 => n11294, B1 => n11386, B2 => 
                           n11293, ZN => n1616);
   U716 : OAI22_X1 port map( A1 => n13886, A2 => n11294, B1 => n11387, B2 => 
                           n11292, ZN => n1615);
   U717 : OAI22_X1 port map( A1 => n13887, A2 => n11294, B1 => n11388, B2 => 
                           n11293, ZN => n1614);
   U718 : OAI22_X1 port map( A1 => n13635, A2 => n11294, B1 => n11389, B2 => 
                           n11292, ZN => n1613);
   U719 : OAI22_X1 port map( A1 => n13387, A2 => n11294, B1 => n11390, B2 => 
                           n11292, ZN => n1612);
   U720 : OAI22_X1 port map( A1 => n13888, A2 => n11294, B1 => n11391, B2 => 
                           n11293, ZN => n1611);
   U721 : OAI22_X1 port map( A1 => n13889, A2 => n11294, B1 => n11392, B2 => 
                           n11292, ZN => n1610);
   U722 : OAI22_X1 port map( A1 => n13636, A2 => n11294, B1 => n11393, B2 => 
                           n11293, ZN => n1609);
   U723 : OAI22_X1 port map( A1 => n13637, A2 => n11294, B1 => n11394, B2 => 
                           n11292, ZN => n1608);
   U724 : OAI22_X1 port map( A1 => n13117, A2 => n11294, B1 => n11395, B2 => 
                           n11293, ZN => n1607);
   U725 : OAI22_X1 port map( A1 => n13638, A2 => n11294, B1 => n11396, B2 => 
                           n11292, ZN => n1606);
   U726 : OAI22_X1 port map( A1 => n13118, A2 => n11294, B1 => n11397, B2 => 
                           n11292, ZN => n1605);
   U727 : OAI22_X1 port map( A1 => n13119, A2 => n11294, B1 => n11398, B2 => 
                           n11292, ZN => n1604);
   U728 : OAI22_X1 port map( A1 => n13890, A2 => n11294, B1 => n11399, B2 => 
                           n11292, ZN => n1603);
   U729 : OAI22_X1 port map( A1 => n13891, A2 => n11294, B1 => n11400, B2 => 
                           n11292, ZN => n1602);
   U730 : OAI22_X1 port map( A1 => n13892, A2 => n11294, B1 => n11401, B2 => 
                           n11292, ZN => n1601);
   U731 : OAI22_X1 port map( A1 => n13893, A2 => n11294, B1 => n11403, B2 => 
                           n11292, ZN => n1600);
   U732 : OAI22_X1 port map( A1 => n13894, A2 => n11294, B1 => n11404, B2 => 
                           n11293, ZN => n1599);
   U733 : OAI22_X1 port map( A1 => n13388, A2 => n11294, B1 => n11405, B2 => 
                           n11293, ZN => n1598);
   U734 : OAI22_X1 port map( A1 => n13639, A2 => n11294, B1 => n11406, B2 => 
                           n11293, ZN => n1597);
   U735 : OAI22_X1 port map( A1 => n13389, A2 => n11294, B1 => n11407, B2 => 
                           n11293, ZN => n1596);
   U736 : OAI22_X1 port map( A1 => n13895, A2 => n11294, B1 => n11408, B2 => 
                           n11293, ZN => n1595);
   U737 : OAI22_X1 port map( A1 => n13896, A2 => n11294, B1 => n11409, B2 => 
                           n11293, ZN => n1594);
   U738 : OAI22_X1 port map( A1 => n13897, A2 => n11294, B1 => n11410, B2 => 
                           n11293, ZN => n1593);
   U739 : OAI22_X1 port map( A1 => n13640, A2 => n11294, B1 => n11411, B2 => 
                           n11293, ZN => n1592);
   U740 : OAI22_X1 port map( A1 => n13641, A2 => n11294, B1 => n11413, B2 => 
                           n11293, ZN => n1591);
   U741 : NAND2_X1 port map( A1 => n11358, A2 => n11342, ZN => n11316);
   U742 : CLKBUF_X1 port map( A => n11316, Z => n11326);
   U743 : OAI22_X1 port map( A1 => n13243, A2 => n11328, B1 => n11343, B2 => 
                           n11326, ZN => n1590);
   U744 : OAI22_X1 port map( A1 => n13120, A2 => n11328, B1 => n11295, B2 => 
                           n11316, ZN => n1589);
   U745 : OAI22_X1 port map( A1 => n13642, A2 => n11328, B1 => n11296, B2 => 
                           n11326, ZN => n1588);
   U746 : OAI22_X1 port map( A1 => n13390, A2 => n11328, B1 => n11297, B2 => 
                           n11316, ZN => n1587);
   U747 : OAI22_X1 port map( A1 => n13898, A2 => n11328, B1 => n11298, B2 => 
                           n11326, ZN => n1586);
   U748 : OAI22_X1 port map( A1 => n13121, A2 => n11328, B1 => n11299, B2 => 
                           n11316, ZN => n1585);
   U749 : OAI22_X1 port map( A1 => n13643, A2 => n11328, B1 => n11300, B2 => 
                           n11326, ZN => n1584);
   U750 : OAI22_X1 port map( A1 => n13391, A2 => n11328, B1 => n11301, B2 => 
                           n11316, ZN => n1583);
   U751 : OAI22_X1 port map( A1 => n13899, A2 => n11328, B1 => n11302, B2 => 
                           n11326, ZN => n1582);
   U752 : OAI22_X1 port map( A1 => n13122, A2 => n11328, B1 => n11303, B2 => 
                           n11316, ZN => n1581);
   U753 : OAI22_X1 port map( A1 => n13392, A2 => n11328, B1 => n11304, B2 => 
                           n11316, ZN => n1580);
   U754 : OAI22_X1 port map( A1 => n13123, A2 => n11328, B1 => n11305, B2 => 
                           n11326, ZN => n1579);
   U755 : OAI22_X1 port map( A1 => n13124, A2 => n11328, B1 => n11306, B2 => 
                           n11316, ZN => n1578);
   U756 : OAI22_X1 port map( A1 => n13125, A2 => n11328, B1 => n11307, B2 => 
                           n11326, ZN => n1577);
   U757 : OAI22_X1 port map( A1 => n13126, A2 => n11328, B1 => n11308, B2 => 
                           n11316, ZN => n1576);
   U758 : OAI22_X1 port map( A1 => n13900, A2 => n11328, B1 => n11309, B2 => 
                           n11326, ZN => n1575);
   U759 : OAI22_X1 port map( A1 => n13644, A2 => n11328, B1 => n11310, B2 => 
                           n11316, ZN => n1574);
   U760 : OAI22_X1 port map( A1 => n13901, A2 => n11328, B1 => n11311, B2 => 
                           n11316, ZN => n1573);
   U761 : OAI22_X1 port map( A1 => n13645, A2 => n11328, B1 => n11312, B2 => 
                           n11316, ZN => n1572);
   U762 : OAI22_X1 port map( A1 => n13393, A2 => n11328, B1 => n11313, B2 => 
                           n11316, ZN => n1571);
   U763 : OAI22_X1 port map( A1 => n13394, A2 => n11328, B1 => n11314, B2 => 
                           n11316, ZN => n1570);
   U764 : OAI22_X1 port map( A1 => n13395, A2 => n11328, B1 => n11315, B2 => 
                           n11316, ZN => n1569);
   U765 : OAI22_X1 port map( A1 => n13646, A2 => n11328, B1 => n11317, B2 => 
                           n11316, ZN => n1568);
   U766 : OAI22_X1 port map( A1 => n13396, A2 => n11328, B1 => n11318, B2 => 
                           n11326, ZN => n1567);
   U767 : OAI22_X1 port map( A1 => n13127, A2 => n11328, B1 => n11319, B2 => 
                           n11326, ZN => n1566);
   U768 : OAI22_X1 port map( A1 => n13128, A2 => n11328, B1 => n11320, B2 => 
                           n11326, ZN => n1565);
   U769 : OAI22_X1 port map( A1 => n13397, A2 => n11328, B1 => n11321, B2 => 
                           n11326, ZN => n1564);
   U770 : OAI22_X1 port map( A1 => n13129, A2 => n11328, B1 => n11322, B2 => 
                           n11326, ZN => n1563);
   U771 : OAI22_X1 port map( A1 => n13398, A2 => n11328, B1 => n11323, B2 => 
                           n11326, ZN => n1562);
   U772 : OAI22_X1 port map( A1 => n13647, A2 => n11328, B1 => n11324, B2 => 
                           n11326, ZN => n1561);
   U773 : OAI22_X1 port map( A1 => n13902, A2 => n11328, B1 => n11325, B2 => 
                           n11326, ZN => n1560);
   U774 : OAI22_X1 port map( A1 => n13130, A2 => n11328, B1 => n11327, B2 => 
                           n11326, ZN => n1559);
   U775 : NAND2_X1 port map( A1 => n11362, A2 => n11342, ZN => n11329);
   U776 : CLKBUF_X1 port map( A => n11329, Z => n11330);
   U777 : OAI22_X1 port map( A1 => n12980, A2 => n11331, B1 => n11343, B2 => 
                           n11330, ZN => n1558);
   U778 : OAI22_X1 port map( A1 => n13399, A2 => n11331, B1 => n11381, B2 => 
                           n11329, ZN => n1557);
   U779 : OAI22_X1 port map( A1 => n13131, A2 => n11331, B1 => n11382, B2 => 
                           n11330, ZN => n1556);
   U780 : OAI22_X1 port map( A1 => n13132, A2 => n11331, B1 => n11383, B2 => 
                           n11329, ZN => n1555);
   U781 : OAI22_X1 port map( A1 => n13133, A2 => n11331, B1 => n11384, B2 => 
                           n11330, ZN => n1554);
   U782 : OAI22_X1 port map( A1 => n13400, A2 => n11331, B1 => n11385, B2 => 
                           n11329, ZN => n1553);
   U783 : OAI22_X1 port map( A1 => n13401, A2 => n11331, B1 => n11386, B2 => 
                           n11330, ZN => n1552);
   U784 : OAI22_X1 port map( A1 => n13402, A2 => n11331, B1 => n11387, B2 => 
                           n11329, ZN => n1551);
   U785 : OAI22_X1 port map( A1 => n13134, A2 => n11331, B1 => n11388, B2 => 
                           n11330, ZN => n1550);
   U786 : OAI22_X1 port map( A1 => n13135, A2 => n11331, B1 => n11389, B2 => 
                           n11329, ZN => n1549);
   U787 : OAI22_X1 port map( A1 => n13403, A2 => n11331, B1 => n11390, B2 => 
                           n11329, ZN => n1548);
   U788 : OAI22_X1 port map( A1 => n13404, A2 => n11331, B1 => n11391, B2 => 
                           n11330, ZN => n1547);
   U789 : OAI22_X1 port map( A1 => n13136, A2 => n11331, B1 => n11392, B2 => 
                           n11329, ZN => n1546);
   U790 : OAI22_X1 port map( A1 => n13405, A2 => n11331, B1 => n11393, B2 => 
                           n11330, ZN => n1545);
   U791 : OAI22_X1 port map( A1 => n13406, A2 => n11331, B1 => n11394, B2 => 
                           n11329, ZN => n1544);
   U792 : OAI22_X1 port map( A1 => n13137, A2 => n11331, B1 => n11395, B2 => 
                           n11330, ZN => n1543);
   U793 : OAI22_X1 port map( A1 => n13407, A2 => n11331, B1 => n11396, B2 => 
                           n11329, ZN => n1542);
   U794 : OAI22_X1 port map( A1 => n13138, A2 => n11331, B1 => n11397, B2 => 
                           n11329, ZN => n1541);
   U795 : OAI22_X1 port map( A1 => n13408, A2 => n11331, B1 => n11398, B2 => 
                           n11329, ZN => n1540);
   U796 : OAI22_X1 port map( A1 => n13139, A2 => n11331, B1 => n11399, B2 => 
                           n11329, ZN => n1539);
   U797 : OAI22_X1 port map( A1 => n13140, A2 => n11331, B1 => n11400, B2 => 
                           n11329, ZN => n1538);
   U798 : OAI22_X1 port map( A1 => n13409, A2 => n11331, B1 => n11401, B2 => 
                           n11329, ZN => n1537);
   U799 : OAI22_X1 port map( A1 => n13141, A2 => n11331, B1 => n11403, B2 => 
                           n11329, ZN => n1536);
   U800 : OAI22_X1 port map( A1 => n13410, A2 => n11331, B1 => n11404, B2 => 
                           n11330, ZN => n1535);
   U801 : OAI22_X1 port map( A1 => n13142, A2 => n11331, B1 => n11405, B2 => 
                           n11330, ZN => n1534);
   U802 : OAI22_X1 port map( A1 => n13143, A2 => n11331, B1 => n11406, B2 => 
                           n11330, ZN => n1533);
   U803 : OAI22_X1 port map( A1 => n13144, A2 => n11331, B1 => n11407, B2 => 
                           n11330, ZN => n1532);
   U804 : OAI22_X1 port map( A1 => n13411, A2 => n11331, B1 => n11408, B2 => 
                           n11330, ZN => n1531);
   U805 : OAI22_X1 port map( A1 => n13412, A2 => n11331, B1 => n11409, B2 => 
                           n11330, ZN => n1530);
   U806 : OAI22_X1 port map( A1 => n13145, A2 => n11331, B1 => n11410, B2 => 
                           n11330, ZN => n1529);
   U807 : OAI22_X1 port map( A1 => n13413, A2 => n11331, B1 => n11411, B2 => 
                           n11330, ZN => n1528);
   U808 : OAI22_X1 port map( A1 => n13146, A2 => n11331, B1 => n11413, B2 => 
                           n11330, ZN => n1527);
   U809 : NAND2_X1 port map( A1 => n11366, A2 => n11342, ZN => n11332);
   U810 : CLKBUF_X1 port map( A => n11335, Z => n11333);
   U811 : CLKBUF_X1 port map( A => n11332, Z => n11334);
   U812 : OAI22_X1 port map( A1 => n13244, A2 => n11333, B1 => n11343, B2 => 
                           n11334, ZN => n1526);
   U813 : OAI22_X1 port map( A1 => n13903, A2 => n11335, B1 => n11381, B2 => 
                           n11332, ZN => n1525);
   U814 : OAI22_X1 port map( A1 => n13414, A2 => n11333, B1 => n11382, B2 => 
                           n11334, ZN => n1524);
   U815 : OAI22_X1 port map( A1 => n13904, A2 => n11335, B1 => n11383, B2 => 
                           n11332, ZN => n1523);
   U816 : OAI22_X1 port map( A1 => n13648, A2 => n11333, B1 => n11384, B2 => 
                           n11334, ZN => n1522);
   U817 : OAI22_X1 port map( A1 => n13415, A2 => n11335, B1 => n11385, B2 => 
                           n11332, ZN => n1521);
   U818 : OAI22_X1 port map( A1 => n13147, A2 => n11333, B1 => n11386, B2 => 
                           n11334, ZN => n1520);
   U819 : OAI22_X1 port map( A1 => n13649, A2 => n11335, B1 => n11387, B2 => 
                           n11332, ZN => n1519);
   U820 : OAI22_X1 port map( A1 => n13650, A2 => n11333, B1 => n11388, B2 => 
                           n11334, ZN => n1518);
   U821 : OAI22_X1 port map( A1 => n13905, A2 => n11335, B1 => n11389, B2 => 
                           n11332, ZN => n1517);
   U822 : OAI22_X1 port map( A1 => n13906, A2 => n11335, B1 => n11390, B2 => 
                           n11332, ZN => n1516);
   U823 : OAI22_X1 port map( A1 => n13651, A2 => n11335, B1 => n11391, B2 => 
                           n11334, ZN => n1515);
   U824 : OAI22_X1 port map( A1 => n13907, A2 => n11333, B1 => n11392, B2 => 
                           n11332, ZN => n1514);
   U825 : OAI22_X1 port map( A1 => n13416, A2 => n11333, B1 => n11393, B2 => 
                           n11334, ZN => n1513);
   U826 : OAI22_X1 port map( A1 => n13652, A2 => n11333, B1 => n11394, B2 => 
                           n11332, ZN => n1512);
   U827 : OAI22_X1 port map( A1 => n13653, A2 => n11333, B1 => n11395, B2 => 
                           n11334, ZN => n1511);
   U828 : OAI22_X1 port map( A1 => n13654, A2 => n11333, B1 => n11396, B2 => 
                           n11332, ZN => n1510);
   U829 : OAI22_X1 port map( A1 => n13908, A2 => n11333, B1 => n11397, B2 => 
                           n11332, ZN => n1509);
   U830 : OAI22_X1 port map( A1 => n13909, A2 => n11333, B1 => n11398, B2 => 
                           n11332, ZN => n1508);
   U831 : OAI22_X1 port map( A1 => n13910, A2 => n11333, B1 => n11399, B2 => 
                           n11332, ZN => n1507);
   U832 : OAI22_X1 port map( A1 => n13417, A2 => n11333, B1 => n11400, B2 => 
                           n11332, ZN => n1506);
   U833 : OAI22_X1 port map( A1 => n13655, A2 => n11333, B1 => n11401, B2 => 
                           n11332, ZN => n1505);
   U834 : OAI22_X1 port map( A1 => n13911, A2 => n11333, B1 => n11403, B2 => 
                           n11332, ZN => n1504);
   U835 : OAI22_X1 port map( A1 => n13656, A2 => n11333, B1 => n11404, B2 => 
                           n11334, ZN => n1503);
   U836 : OAI22_X1 port map( A1 => n13912, A2 => n11335, B1 => n11405, B2 => 
                           n11334, ZN => n1502);
   U837 : OAI22_X1 port map( A1 => n13913, A2 => n11335, B1 => n11406, B2 => 
                           n11334, ZN => n1501);
   U838 : OAI22_X1 port map( A1 => n13657, A2 => n11335, B1 => n11407, B2 => 
                           n11334, ZN => n1500);
   U839 : OAI22_X1 port map( A1 => n13658, A2 => n11335, B1 => n11408, B2 => 
                           n11334, ZN => n1499);
   U840 : OAI22_X1 port map( A1 => n13659, A2 => n11335, B1 => n11409, B2 => 
                           n11334, ZN => n1498);
   U841 : OAI22_X1 port map( A1 => n13660, A2 => n11335, B1 => n11410, B2 => 
                           n11334, ZN => n1497);
   U842 : OAI22_X1 port map( A1 => n13914, A2 => n11335, B1 => n11411, B2 => 
                           n11334, ZN => n1496);
   U843 : OAI22_X1 port map( A1 => n13661, A2 => n11335, B1 => n11413, B2 => 
                           n11334, ZN => n1495);
   U844 : NAND2_X1 port map( A1 => n11370, A2 => n11342, ZN => n11336);
   U845 : CLKBUF_X1 port map( A => n11336, Z => n11337);
   U846 : OAI22_X1 port map( A1 => n13245, A2 => n11338, B1 => n11343, B2 => 
                           n11337, ZN => n1494);
   U847 : OAI22_X1 port map( A1 => n13915, A2 => n11338, B1 => n11381, B2 => 
                           n11336, ZN => n1493);
   U848 : OAI22_X1 port map( A1 => n13662, A2 => n11338, B1 => n11382, B2 => 
                           n11337, ZN => n1492);
   U849 : OAI22_X1 port map( A1 => n13916, A2 => n11338, B1 => n11383, B2 => 
                           n11336, ZN => n1491);
   U850 : OAI22_X1 port map( A1 => n13663, A2 => n11338, B1 => n11384, B2 => 
                           n11337, ZN => n1490);
   U851 : OAI22_X1 port map( A1 => n13917, A2 => n11338, B1 => n11385, B2 => 
                           n11336, ZN => n1489);
   U852 : OAI22_X1 port map( A1 => n13918, A2 => n11338, B1 => n11386, B2 => 
                           n11337, ZN => n1488);
   U853 : OAI22_X1 port map( A1 => n13664, A2 => n11338, B1 => n11387, B2 => 
                           n11336, ZN => n1487);
   U854 : OAI22_X1 port map( A1 => n13665, A2 => n11338, B1 => n11388, B2 => 
                           n11337, ZN => n1486);
   U855 : OAI22_X1 port map( A1 => n13919, A2 => n11338, B1 => n11389, B2 => 
                           n11336, ZN => n1485);
   U856 : OAI22_X1 port map( A1 => n13666, A2 => n11338, B1 => n11390, B2 => 
                           n11336, ZN => n1484);
   U857 : OAI22_X1 port map( A1 => n13920, A2 => n11338, B1 => n11391, B2 => 
                           n11337, ZN => n1483);
   U858 : OAI22_X1 port map( A1 => n13667, A2 => n11338, B1 => n11392, B2 => 
                           n11336, ZN => n1482);
   U859 : OAI22_X1 port map( A1 => n13668, A2 => n11338, B1 => n11393, B2 => 
                           n11337, ZN => n1481);
   U860 : OAI22_X1 port map( A1 => n13669, A2 => n11338, B1 => n11394, B2 => 
                           n11336, ZN => n1480);
   U861 : OAI22_X1 port map( A1 => n13921, A2 => n11338, B1 => n11395, B2 => 
                           n11337, ZN => n1479);
   U862 : OAI22_X1 port map( A1 => n13922, A2 => n11338, B1 => n11396, B2 => 
                           n11336, ZN => n1478);
   U863 : OAI22_X1 port map( A1 => n13670, A2 => n11338, B1 => n11397, B2 => 
                           n11336, ZN => n1477);
   U864 : OAI22_X1 port map( A1 => n13923, A2 => n11338, B1 => n11398, B2 => 
                           n11336, ZN => n1476);
   U865 : OAI22_X1 port map( A1 => n13924, A2 => n11338, B1 => n11399, B2 => 
                           n11336, ZN => n1475);
   U866 : OAI22_X1 port map( A1 => n13671, A2 => n11338, B1 => n11400, B2 => 
                           n11336, ZN => n1474);
   U867 : OAI22_X1 port map( A1 => n13672, A2 => n11338, B1 => n11401, B2 => 
                           n11336, ZN => n1473);
   U868 : OAI22_X1 port map( A1 => n13925, A2 => n11338, B1 => n11403, B2 => 
                           n11336, ZN => n1472);
   U869 : OAI22_X1 port map( A1 => n13673, A2 => n11338, B1 => n11404, B2 => 
                           n11337, ZN => n1471);
   U870 : OAI22_X1 port map( A1 => n13674, A2 => n11338, B1 => n11405, B2 => 
                           n11337, ZN => n1470);
   U871 : OAI22_X1 port map( A1 => n13926, A2 => n11338, B1 => n11406, B2 => 
                           n11337, ZN => n1469);
   U872 : OAI22_X1 port map( A1 => n13927, A2 => n11338, B1 => n11407, B2 => 
                           n11337, ZN => n1468);
   U873 : OAI22_X1 port map( A1 => n13928, A2 => n11338, B1 => n11408, B2 => 
                           n11337, ZN => n1467);
   U874 : OAI22_X1 port map( A1 => n13929, A2 => n11338, B1 => n11409, B2 => 
                           n11337, ZN => n1466);
   U875 : OAI22_X1 port map( A1 => n13930, A2 => n11338, B1 => n11410, B2 => 
                           n11337, ZN => n1465);
   U876 : OAI22_X1 port map( A1 => n13418, A2 => n11338, B1 => n11411, B2 => 
                           n11337, ZN => n1464);
   U877 : OAI22_X1 port map( A1 => n13931, A2 => n11338, B1 => n11413, B2 => 
                           n11337, ZN => n1463);
   U878 : NAND2_X1 port map( A1 => n11374, A2 => n11342, ZN => n11339);
   U879 : CLKBUF_X1 port map( A => n11339, Z => n11340);
   U880 : OAI22_X1 port map( A1 => n13495, A2 => n11341, B1 => n11343, B2 => 
                           n11340, ZN => n1462);
   U881 : OAI22_X1 port map( A1 => n13932, A2 => n11341, B1 => n11381, B2 => 
                           n11339, ZN => n1461);
   U882 : OAI22_X1 port map( A1 => n13933, A2 => n11341, B1 => n11382, B2 => 
                           n11340, ZN => n1460);
   U883 : OAI22_X1 port map( A1 => n13934, A2 => n11341, B1 => n11383, B2 => 
                           n11339, ZN => n1459);
   U884 : OAI22_X1 port map( A1 => n13675, A2 => n11341, B1 => n11384, B2 => 
                           n11340, ZN => n1458);
   U885 : OAI22_X1 port map( A1 => n13935, A2 => n11341, B1 => n11385, B2 => 
                           n11339, ZN => n1457);
   U886 : OAI22_X1 port map( A1 => n13676, A2 => n11341, B1 => n11386, B2 => 
                           n11340, ZN => n1456);
   U887 : OAI22_X1 port map( A1 => n13677, A2 => n11341, B1 => n11387, B2 => 
                           n11339, ZN => n1455);
   U888 : OAI22_X1 port map( A1 => n13678, A2 => n11341, B1 => n11388, B2 => 
                           n11340, ZN => n1454);
   U889 : OAI22_X1 port map( A1 => n13936, A2 => n11341, B1 => n11389, B2 => 
                           n11339, ZN => n1453);
   U890 : OAI22_X1 port map( A1 => n13937, A2 => n11341, B1 => n11390, B2 => 
                           n11339, ZN => n1452);
   U891 : OAI22_X1 port map( A1 => n13148, A2 => n11341, B1 => n11391, B2 => 
                           n11340, ZN => n1451);
   U892 : OAI22_X1 port map( A1 => n13679, A2 => n11341, B1 => n11392, B2 => 
                           n11339, ZN => n1450);
   U893 : OAI22_X1 port map( A1 => n13680, A2 => n11341, B1 => n11393, B2 => 
                           n11340, ZN => n1449);
   U894 : OAI22_X1 port map( A1 => n13681, A2 => n11341, B1 => n11394, B2 => 
                           n11339, ZN => n1448);
   U895 : OAI22_X1 port map( A1 => n13682, A2 => n11341, B1 => n11395, B2 => 
                           n11340, ZN => n1447);
   U896 : OAI22_X1 port map( A1 => n13419, A2 => n11341, B1 => n11396, B2 => 
                           n11339, ZN => n1446);
   U897 : OAI22_X1 port map( A1 => n13683, A2 => n11341, B1 => n11397, B2 => 
                           n11339, ZN => n1445);
   U898 : OAI22_X1 port map( A1 => n13684, A2 => n11341, B1 => n11398, B2 => 
                           n11339, ZN => n1444);
   U899 : OAI22_X1 port map( A1 => n13685, A2 => n11341, B1 => n11399, B2 => 
                           n11339, ZN => n1443);
   U900 : OAI22_X1 port map( A1 => n13149, A2 => n11341, B1 => n11400, B2 => 
                           n11339, ZN => n1442);
   U901 : OAI22_X1 port map( A1 => n13686, A2 => n11341, B1 => n11401, B2 => 
                           n11339, ZN => n1441);
   U902 : OAI22_X1 port map( A1 => n13938, A2 => n11341, B1 => n11403, B2 => 
                           n11339, ZN => n1440);
   U903 : OAI22_X1 port map( A1 => n13150, A2 => n11341, B1 => n11404, B2 => 
                           n11340, ZN => n1439);
   U904 : OAI22_X1 port map( A1 => n13420, A2 => n11341, B1 => n11405, B2 => 
                           n11340, ZN => n1438);
   U905 : OAI22_X1 port map( A1 => n13687, A2 => n11341, B1 => n11406, B2 => 
                           n11340, ZN => n1437);
   U906 : OAI22_X1 port map( A1 => n13688, A2 => n11341, B1 => n11407, B2 => 
                           n11340, ZN => n1436);
   U907 : OAI22_X1 port map( A1 => n13939, A2 => n11341, B1 => n11408, B2 => 
                           n11340, ZN => n1435);
   U908 : OAI22_X1 port map( A1 => n13940, A2 => n11341, B1 => n11409, B2 => 
                           n11340, ZN => n1434);
   U909 : OAI22_X1 port map( A1 => n13941, A2 => n11341, B1 => n11410, B2 => 
                           n11340, ZN => n1433);
   U910 : OAI22_X1 port map( A1 => n13689, A2 => n11341, B1 => n11411, B2 => 
                           n11340, ZN => n1432);
   U911 : OAI22_X1 port map( A1 => n13942, A2 => n11341, B1 => n11413, B2 => 
                           n11340, ZN => n1431);
   U912 : NAND2_X1 port map( A1 => n11379, A2 => n11342, ZN => n11344);
   U913 : CLKBUF_X1 port map( A => n11344, Z => n11345);
   U914 : OAI22_X1 port map( A1 => n12981, A2 => n11346, B1 => n11343, B2 => 
                           n11345, ZN => n1430);
   U915 : OAI22_X1 port map( A1 => n13151, A2 => n11346, B1 => n11381, B2 => 
                           n11344, ZN => n1429);
   U916 : OAI22_X1 port map( A1 => n13152, A2 => n11346, B1 => n11382, B2 => 
                           n11345, ZN => n1428);
   U917 : OAI22_X1 port map( A1 => n13153, A2 => n11346, B1 => n11383, B2 => 
                           n11344, ZN => n1427);
   U918 : OAI22_X1 port map( A1 => n13154, A2 => n11346, B1 => n11384, B2 => 
                           n11345, ZN => n1426);
   U919 : OAI22_X1 port map( A1 => n13155, A2 => n11346, B1 => n11385, B2 => 
                           n11344, ZN => n1425);
   U920 : OAI22_X1 port map( A1 => n13156, A2 => n11346, B1 => n11386, B2 => 
                           n11345, ZN => n1424);
   U921 : OAI22_X1 port map( A1 => n13943, A2 => n11346, B1 => n11387, B2 => 
                           n11344, ZN => n1423);
   U922 : OAI22_X1 port map( A1 => n13421, A2 => n11346, B1 => n11388, B2 => 
                           n11345, ZN => n1422);
   U923 : OAI22_X1 port map( A1 => n13422, A2 => n11346, B1 => n11389, B2 => 
                           n11344, ZN => n1421);
   U924 : OAI22_X1 port map( A1 => n13157, A2 => n11346, B1 => n11390, B2 => 
                           n11344, ZN => n1420);
   U925 : OAI22_X1 port map( A1 => n13158, A2 => n11346, B1 => n11391, B2 => 
                           n11345, ZN => n1419);
   U926 : OAI22_X1 port map( A1 => n13423, A2 => n11346, B1 => n11392, B2 => 
                           n11344, ZN => n1418);
   U927 : OAI22_X1 port map( A1 => n13159, A2 => n11346, B1 => n11393, B2 => 
                           n11345, ZN => n1417);
   U928 : OAI22_X1 port map( A1 => n13424, A2 => n11346, B1 => n11394, B2 => 
                           n11344, ZN => n1416);
   U929 : OAI22_X1 port map( A1 => n13425, A2 => n11346, B1 => n11395, B2 => 
                           n11345, ZN => n1415);
   U930 : OAI22_X1 port map( A1 => n13160, A2 => n11346, B1 => n11396, B2 => 
                           n11344, ZN => n1414);
   U931 : OAI22_X1 port map( A1 => n13426, A2 => n11346, B1 => n11397, B2 => 
                           n11344, ZN => n1413);
   U932 : OAI22_X1 port map( A1 => n13161, A2 => n11346, B1 => n11398, B2 => 
                           n11344, ZN => n1412);
   U933 : OAI22_X1 port map( A1 => n13427, A2 => n11346, B1 => n11399, B2 => 
                           n11344, ZN => n1411);
   U934 : OAI22_X1 port map( A1 => n13428, A2 => n11346, B1 => n11400, B2 => 
                           n11344, ZN => n1410);
   U935 : OAI22_X1 port map( A1 => n13162, A2 => n11346, B1 => n11401, B2 => 
                           n11344, ZN => n1409);
   U936 : OAI22_X1 port map( A1 => n13429, A2 => n11346, B1 => n11403, B2 => 
                           n11344, ZN => n1408);
   U937 : OAI22_X1 port map( A1 => n13944, A2 => n11346, B1 => n11404, B2 => 
                           n11345, ZN => n1407);
   U938 : OAI22_X1 port map( A1 => n13690, A2 => n11346, B1 => n11405, B2 => 
                           n11345, ZN => n1406);
   U939 : OAI22_X1 port map( A1 => n13163, A2 => n11346, B1 => n11406, B2 => 
                           n11345, ZN => n1405);
   U940 : OAI22_X1 port map( A1 => n13691, A2 => n11346, B1 => n11407, B2 => 
                           n11345, ZN => n1404);
   U941 : OAI22_X1 port map( A1 => n13164, A2 => n11346, B1 => n11408, B2 => 
                           n11345, ZN => n1403);
   U942 : OAI22_X1 port map( A1 => n13692, A2 => n11346, B1 => n11409, B2 => 
                           n11345, ZN => n1402);
   U943 : OAI22_X1 port map( A1 => n13430, A2 => n11346, B1 => n11410, B2 => 
                           n11345, ZN => n1401);
   U944 : OAI22_X1 port map( A1 => n13693, A2 => n11346, B1 => n11411, B2 => 
                           n11345, ZN => n1400);
   U945 : OAI22_X1 port map( A1 => n13165, A2 => n11346, B1 => n11413, B2 => 
                           n11345, ZN => n1399);
   U946 : NAND2_X1 port map( A1 => n11349, A2 => n11378, ZN => n11350);
   U947 : CLKBUF_X1 port map( A => n11353, Z => n11351);
   U948 : CLKBUF_X1 port map( A => n11350, Z => n11352);
   U949 : OAI22_X1 port map( A1 => n12982, A2 => n11351, B1 => n11380, B2 => 
                           n11352, ZN => n1398);
   U950 : OAI22_X1 port map( A1 => n13431, A2 => n11353, B1 => n11381, B2 => 
                           n11350, ZN => n1397);
   U951 : OAI22_X1 port map( A1 => n13694, A2 => n11351, B1 => n11382, B2 => 
                           n11352, ZN => n1396);
   U952 : OAI22_X1 port map( A1 => n13166, A2 => n11353, B1 => n11383, B2 => 
                           n11350, ZN => n1395);
   U953 : OAI22_X1 port map( A1 => n13432, A2 => n11351, B1 => n11384, B2 => 
                           n11352, ZN => n1394);
   U954 : OAI22_X1 port map( A1 => n13167, A2 => n11353, B1 => n11385, B2 => 
                           n11350, ZN => n1393);
   U955 : OAI22_X1 port map( A1 => n13168, A2 => n11351, B1 => n11386, B2 => 
                           n11352, ZN => n1392);
   U956 : OAI22_X1 port map( A1 => n13169, A2 => n11353, B1 => n11387, B2 => 
                           n11350, ZN => n1391);
   U957 : OAI22_X1 port map( A1 => n13170, A2 => n11351, B1 => n11388, B2 => 
                           n11352, ZN => n1390);
   U958 : OAI22_X1 port map( A1 => n13695, A2 => n11353, B1 => n11389, B2 => 
                           n11350, ZN => n1389);
   U959 : OAI22_X1 port map( A1 => n13433, A2 => n11353, B1 => n11390, B2 => 
                           n11350, ZN => n1388);
   U960 : OAI22_X1 port map( A1 => n13434, A2 => n11353, B1 => n11391, B2 => 
                           n11352, ZN => n1387);
   U961 : OAI22_X1 port map( A1 => n13435, A2 => n11351, B1 => n11392, B2 => 
                           n11350, ZN => n1386);
   U962 : OAI22_X1 port map( A1 => n13436, A2 => n11351, B1 => n11393, B2 => 
                           n11352, ZN => n1385);
   U963 : OAI22_X1 port map( A1 => n13437, A2 => n11351, B1 => n11394, B2 => 
                           n11350, ZN => n1384);
   U964 : OAI22_X1 port map( A1 => n13171, A2 => n11351, B1 => n11395, B2 => 
                           n11352, ZN => n1383);
   U965 : OAI22_X1 port map( A1 => n13438, A2 => n11351, B1 => n11396, B2 => 
                           n11350, ZN => n1382);
   U966 : OAI22_X1 port map( A1 => n13439, A2 => n11351, B1 => n11397, B2 => 
                           n11350, ZN => n1381);
   U967 : OAI22_X1 port map( A1 => n13172, A2 => n11351, B1 => n11398, B2 => 
                           n11350, ZN => n1380);
   U968 : OAI22_X1 port map( A1 => n13173, A2 => n11351, B1 => n11399, B2 => 
                           n11350, ZN => n1379);
   U969 : OAI22_X1 port map( A1 => n13696, A2 => n11351, B1 => n11400, B2 => 
                           n11350, ZN => n1378);
   U970 : OAI22_X1 port map( A1 => n13440, A2 => n11351, B1 => n11401, B2 => 
                           n11350, ZN => n1377);
   U971 : OAI22_X1 port map( A1 => n13174, A2 => n11351, B1 => n11403, B2 => 
                           n11350, ZN => n1376);
   U972 : OAI22_X1 port map( A1 => n13441, A2 => n11351, B1 => n11404, B2 => 
                           n11352, ZN => n1375);
   U973 : OAI22_X1 port map( A1 => n13175, A2 => n11353, B1 => n11405, B2 => 
                           n11352, ZN => n1374);
   U974 : OAI22_X1 port map( A1 => n13697, A2 => n11353, B1 => n11406, B2 => 
                           n11352, ZN => n1373);
   U975 : OAI22_X1 port map( A1 => n13176, A2 => n11353, B1 => n11407, B2 => 
                           n11352, ZN => n1372);
   U976 : OAI22_X1 port map( A1 => n13177, A2 => n11353, B1 => n11408, B2 => 
                           n11352, ZN => n1371);
   U977 : OAI22_X1 port map( A1 => n13178, A2 => n11353, B1 => n11409, B2 => 
                           n11352, ZN => n1370);
   U978 : OAI22_X1 port map( A1 => n13442, A2 => n11353, B1 => n11410, B2 => 
                           n11352, ZN => n1369);
   U979 : OAI22_X1 port map( A1 => n13179, A2 => n11353, B1 => n11411, B2 => 
                           n11352, ZN => n1368);
   U980 : OAI22_X1 port map( A1 => n13443, A2 => n11353, B1 => n11413, B2 => 
                           n11352, ZN => n1367);
   U981 : NAND2_X1 port map( A1 => n11354, A2 => n11378, ZN => n11355);
   U982 : CLKBUF_X1 port map( A => n11355, Z => n11356);
   U983 : OAI22_X1 port map( A1 => n13246, A2 => n11357, B1 => n11380, B2 => 
                           n11356, ZN => n1366);
   U984 : OAI22_X1 port map( A1 => n13698, A2 => n11357, B1 => n11381, B2 => 
                           n11355, ZN => n1365);
   U985 : OAI22_X1 port map( A1 => n13444, A2 => n11357, B1 => n11382, B2 => 
                           n11356, ZN => n1364);
   U986 : OAI22_X1 port map( A1 => n13180, A2 => n11357, B1 => n11383, B2 => 
                           n11355, ZN => n1363);
   U987 : OAI22_X1 port map( A1 => n13181, A2 => n11357, B1 => n11384, B2 => 
                           n11356, ZN => n1362);
   U988 : OAI22_X1 port map( A1 => n13182, A2 => n11357, B1 => n11385, B2 => 
                           n11355, ZN => n1361);
   U989 : OAI22_X1 port map( A1 => n13445, A2 => n11357, B1 => n11386, B2 => 
                           n11356, ZN => n1360);
   U990 : OAI22_X1 port map( A1 => n13183, A2 => n11357, B1 => n11387, B2 => 
                           n11355, ZN => n1359);
   U991 : OAI22_X1 port map( A1 => n13446, A2 => n11357, B1 => n11388, B2 => 
                           n11356, ZN => n1358);
   U992 : OAI22_X1 port map( A1 => n13184, A2 => n11357, B1 => n11389, B2 => 
                           n11355, ZN => n1357);
   U993 : OAI22_X1 port map( A1 => n13447, A2 => n11357, B1 => n11390, B2 => 
                           n11355, ZN => n1356);
   U994 : OAI22_X1 port map( A1 => n13185, A2 => n11357, B1 => n11391, B2 => 
                           n11356, ZN => n1355);
   U995 : OAI22_X1 port map( A1 => n13945, A2 => n11357, B1 => n11392, B2 => 
                           n11355, ZN => n1354);
   U996 : OAI22_X1 port map( A1 => n13186, A2 => n11357, B1 => n11393, B2 => 
                           n11356, ZN => n1353);
   U997 : OAI22_X1 port map( A1 => n13448, A2 => n11357, B1 => n11394, B2 => 
                           n11355, ZN => n1352);
   U998 : OAI22_X1 port map( A1 => n13699, A2 => n11357, B1 => n11395, B2 => 
                           n11356, ZN => n1351);
   U999 : OAI22_X1 port map( A1 => n13187, A2 => n11357, B1 => n11396, B2 => 
                           n11355, ZN => n1350);
   U1000 : OAI22_X1 port map( A1 => n13449, A2 => n11357, B1 => n11397, B2 => 
                           n11355, ZN => n1349);
   U1001 : OAI22_X1 port map( A1 => n13700, A2 => n11357, B1 => n11398, B2 => 
                           n11355, ZN => n1348);
   U1002 : OAI22_X1 port map( A1 => n13946, A2 => n11357, B1 => n11399, B2 => 
                           n11355, ZN => n1347);
   U1003 : OAI22_X1 port map( A1 => n13450, A2 => n11357, B1 => n11400, B2 => 
                           n11355, ZN => n1346);
   U1004 : OAI22_X1 port map( A1 => n13188, A2 => n11357, B1 => n11401, B2 => 
                           n11355, ZN => n1345);
   U1005 : OAI22_X1 port map( A1 => n13189, A2 => n11357, B1 => n11403, B2 => 
                           n11355, ZN => n1344);
   U1006 : OAI22_X1 port map( A1 => n13190, A2 => n11357, B1 => n11404, B2 => 
                           n11356, ZN => n1343);
   U1007 : OAI22_X1 port map( A1 => n13191, A2 => n11357, B1 => n11405, B2 => 
                           n11356, ZN => n1342);
   U1008 : OAI22_X1 port map( A1 => n13451, A2 => n11357, B1 => n11406, B2 => 
                           n11356, ZN => n1341);
   U1009 : OAI22_X1 port map( A1 => n13452, A2 => n11357, B1 => n11407, B2 => 
                           n11356, ZN => n1340);
   U1010 : OAI22_X1 port map( A1 => n13701, A2 => n11357, B1 => n11408, B2 => 
                           n11356, ZN => n1339);
   U1011 : OAI22_X1 port map( A1 => n13453, A2 => n11357, B1 => n11409, B2 => 
                           n11356, ZN => n1338);
   U1012 : OAI22_X1 port map( A1 => n13192, A2 => n11357, B1 => n11410, B2 => 
                           n11356, ZN => n1337);
   U1013 : OAI22_X1 port map( A1 => n13193, A2 => n11357, B1 => n11411, B2 => 
                           n11356, ZN => n1336);
   U1014 : OAI22_X1 port map( A1 => n13454, A2 => n11357, B1 => n11413, B2 => 
                           n11356, ZN => n1335);
   U1015 : NAND2_X1 port map( A1 => n11358, A2 => n11378, ZN => n11359);
   U1016 : CLKBUF_X1 port map( A => n11359, Z => n11360);
   U1017 : OAI22_X1 port map( A1 => n13496, A2 => n11361, B1 => n11380, B2 => 
                           n11360, ZN => n1334);
   U1018 : OAI22_X1 port map( A1 => n13194, A2 => n11361, B1 => n11381, B2 => 
                           n11359, ZN => n1333);
   U1019 : OAI22_X1 port map( A1 => n13455, A2 => n11361, B1 => n11382, B2 => 
                           n11360, ZN => n1332);
   U1020 : OAI22_X1 port map( A1 => n13947, A2 => n11361, B1 => n11383, B2 => 
                           n11359, ZN => n1331);
   U1021 : OAI22_X1 port map( A1 => n13948, A2 => n11361, B1 => n11384, B2 => 
                           n11360, ZN => n1330);
   U1022 : OAI22_X1 port map( A1 => n13702, A2 => n11361, B1 => n11385, B2 => 
                           n11359, ZN => n1329);
   U1023 : OAI22_X1 port map( A1 => n13949, A2 => n11361, B1 => n11386, B2 => 
                           n11360, ZN => n1328);
   U1024 : OAI22_X1 port map( A1 => n13950, A2 => n11361, B1 => n11387, B2 => 
                           n11359, ZN => n1327);
   U1025 : OAI22_X1 port map( A1 => n13951, A2 => n11361, B1 => n11388, B2 => 
                           n11360, ZN => n1326);
   U1026 : OAI22_X1 port map( A1 => n13703, A2 => n11361, B1 => n11389, B2 => 
                           n11359, ZN => n1325);
   U1027 : OAI22_X1 port map( A1 => n13704, A2 => n11361, B1 => n11390, B2 => 
                           n11359, ZN => n1324);
   U1028 : OAI22_X1 port map( A1 => n13456, A2 => n11361, B1 => n11391, B2 => 
                           n11360, ZN => n1323);
   U1029 : OAI22_X1 port map( A1 => n13705, A2 => n11361, B1 => n11392, B2 => 
                           n11359, ZN => n1322);
   U1030 : OAI22_X1 port map( A1 => n13952, A2 => n11361, B1 => n11393, B2 => 
                           n11360, ZN => n1321);
   U1031 : OAI22_X1 port map( A1 => n13953, A2 => n11361, B1 => n11394, B2 => 
                           n11359, ZN => n1320);
   U1032 : OAI22_X1 port map( A1 => n13954, A2 => n11361, B1 => n11395, B2 => 
                           n11360, ZN => n1319);
   U1033 : OAI22_X1 port map( A1 => n13706, A2 => n11361, B1 => n11396, B2 => 
                           n11359, ZN => n1318);
   U1034 : OAI22_X1 port map( A1 => n13707, A2 => n11361, B1 => n11397, B2 => 
                           n11359, ZN => n1317);
   U1035 : OAI22_X1 port map( A1 => n13708, A2 => n11361, B1 => n11398, B2 => 
                           n11359, ZN => n1316);
   U1036 : OAI22_X1 port map( A1 => n13709, A2 => n11361, B1 => n11399, B2 => 
                           n11359, ZN => n1315);
   U1037 : OAI22_X1 port map( A1 => n13710, A2 => n11361, B1 => n11400, B2 => 
                           n11359, ZN => n1314);
   U1038 : OAI22_X1 port map( A1 => n13457, A2 => n11361, B1 => n11401, B2 => 
                           n11359, ZN => n1313);
   U1039 : OAI22_X1 port map( A1 => n13195, A2 => n11361, B1 => n11403, B2 => 
                           n11359, ZN => n1312);
   U1040 : OAI22_X1 port map( A1 => n13711, A2 => n11361, B1 => n11404, B2 => 
                           n11360, ZN => n1311);
   U1041 : OAI22_X1 port map( A1 => n13955, A2 => n11361, B1 => n11405, B2 => 
                           n11360, ZN => n1310);
   U1042 : OAI22_X1 port map( A1 => n13458, A2 => n11361, B1 => n11406, B2 => 
                           n11360, ZN => n1309);
   U1043 : OAI22_X1 port map( A1 => n13459, A2 => n11361, B1 => n11407, B2 => 
                           n11360, ZN => n1308);
   U1044 : OAI22_X1 port map( A1 => n13460, A2 => n11361, B1 => n11408, B2 => 
                           n11360, ZN => n1307);
   U1045 : OAI22_X1 port map( A1 => n13712, A2 => n11361, B1 => n11409, B2 => 
                           n11360, ZN => n1306);
   U1046 : OAI22_X1 port map( A1 => n13956, A2 => n11361, B1 => n11410, B2 => 
                           n11360, ZN => n1305);
   U1047 : OAI22_X1 port map( A1 => n13196, A2 => n11361, B1 => n11411, B2 => 
                           n11360, ZN => n1304);
   U1048 : OAI22_X1 port map( A1 => n13197, A2 => n11361, B1 => n11413, B2 => 
                           n11360, ZN => n1303);
   U1049 : NAND2_X1 port map( A1 => n11362, A2 => n11378, ZN => n11363);
   U1050 : CLKBUF_X1 port map( A => n11363, Z => n11364);
   U1051 : OAI22_X1 port map( A1 => n13247, A2 => n11365, B1 => n11380, B2 => 
                           n11364, ZN => n1302);
   U1052 : OAI22_X1 port map( A1 => n13461, A2 => n11365, B1 => n11381, B2 => 
                           n11363, ZN => n1301);
   U1053 : OAI22_X1 port map( A1 => n13198, A2 => n11365, B1 => n11382, B2 => 
                           n11364, ZN => n1300);
   U1054 : OAI22_X1 port map( A1 => n13462, A2 => n11365, B1 => n11383, B2 => 
                           n11363, ZN => n1299);
   U1055 : OAI22_X1 port map( A1 => n13463, A2 => n11365, B1 => n11384, B2 => 
                           n11364, ZN => n1298);
   U1056 : OAI22_X1 port map( A1 => n13199, A2 => n11365, B1 => n11385, B2 => 
                           n11363, ZN => n1297);
   U1057 : OAI22_X1 port map( A1 => n13957, A2 => n11365, B1 => n11386, B2 => 
                           n11364, ZN => n1296);
   U1058 : OAI22_X1 port map( A1 => n13200, A2 => n11365, B1 => n11387, B2 => 
                           n11363, ZN => n1295);
   U1059 : OAI22_X1 port map( A1 => n13464, A2 => n11365, B1 => n11388, B2 => 
                           n11364, ZN => n1294);
   U1060 : OAI22_X1 port map( A1 => n13465, A2 => n11365, B1 => n11389, B2 => 
                           n11363, ZN => n1293);
   U1061 : OAI22_X1 port map( A1 => n13201, A2 => n11365, B1 => n11390, B2 => 
                           n11363, ZN => n1292);
   U1062 : OAI22_X1 port map( A1 => n13958, A2 => n11365, B1 => n11391, B2 => 
                           n11364, ZN => n1291);
   U1063 : OAI22_X1 port map( A1 => n13202, A2 => n11365, B1 => n11392, B2 => 
                           n11363, ZN => n1290);
   U1064 : OAI22_X1 port map( A1 => n13466, A2 => n11365, B1 => n11393, B2 => 
                           n11364, ZN => n1289);
   U1065 : OAI22_X1 port map( A1 => n13203, A2 => n11365, B1 => n11394, B2 => 
                           n11363, ZN => n1288);
   U1066 : OAI22_X1 port map( A1 => n13467, A2 => n11365, B1 => n11395, B2 => 
                           n11364, ZN => n1287);
   U1067 : OAI22_X1 port map( A1 => n13204, A2 => n11365, B1 => n11396, B2 => 
                           n11363, ZN => n1286);
   U1068 : OAI22_X1 port map( A1 => n13713, A2 => n11365, B1 => n11397, B2 => 
                           n11363, ZN => n1285);
   U1069 : OAI22_X1 port map( A1 => n13205, A2 => n11365, B1 => n11398, B2 => 
                           n11363, ZN => n1284);
   U1070 : OAI22_X1 port map( A1 => n13206, A2 => n11365, B1 => n11399, B2 => 
                           n11363, ZN => n1283);
   U1071 : OAI22_X1 port map( A1 => n13207, A2 => n11365, B1 => n11400, B2 => 
                           n11363, ZN => n1282);
   U1072 : OAI22_X1 port map( A1 => n13468, A2 => n11365, B1 => n11401, B2 => 
                           n11363, ZN => n1281);
   U1073 : OAI22_X1 port map( A1 => n13208, A2 => n11365, B1 => n11403, B2 => 
                           n11363, ZN => n1280);
   U1074 : OAI22_X1 port map( A1 => n13209, A2 => n11365, B1 => n11404, B2 => 
                           n11364, ZN => n1279);
   U1075 : OAI22_X1 port map( A1 => n13714, A2 => n11365, B1 => n11405, B2 => 
                           n11364, ZN => n1278);
   U1076 : OAI22_X1 port map( A1 => n13210, A2 => n11365, B1 => n11406, B2 => 
                           n11364, ZN => n1277);
   U1077 : OAI22_X1 port map( A1 => n13469, A2 => n11365, B1 => n11407, B2 => 
                           n11364, ZN => n1276);
   U1078 : OAI22_X1 port map( A1 => n13470, A2 => n11365, B1 => n11408, B2 => 
                           n11364, ZN => n1275);
   U1079 : OAI22_X1 port map( A1 => n13211, A2 => n11365, B1 => n11409, B2 => 
                           n11364, ZN => n1274);
   U1080 : OAI22_X1 port map( A1 => n13212, A2 => n11365, B1 => n11410, B2 => 
                           n11364, ZN => n1273);
   U1081 : OAI22_X1 port map( A1 => n13471, A2 => n11365, B1 => n11411, B2 => 
                           n11364, ZN => n1272);
   U1082 : OAI22_X1 port map( A1 => n13472, A2 => n11365, B1 => n11413, B2 => 
                           n11364, ZN => n1271);
   U1083 : NAND2_X1 port map( A1 => n11366, A2 => n11378, ZN => n11367);
   U1084 : OAI22_X1 port map( A1 => n13248, A2 => n11369, B1 => n11380, B2 => 
                           n11368, ZN => n1270);
   U1085 : OAI22_X1 port map( A1 => n13473, A2 => n11369, B1 => n11381, B2 => 
                           n11367, ZN => n1269);
   U1086 : OAI22_X1 port map( A1 => n13213, A2 => n11369, B1 => n11382, B2 => 
                           n11368, ZN => n1268);
   U1087 : OAI22_X1 port map( A1 => n13715, A2 => n11369, B1 => n11383, B2 => 
                           n11367, ZN => n1267);
   U1088 : OAI22_X1 port map( A1 => n13474, A2 => n11369, B1 => n11384, B2 => 
                           n11368, ZN => n1266);
   U1089 : OAI22_X1 port map( A1 => n13959, A2 => n11369, B1 => n11385, B2 => 
                           n11367, ZN => n1265);
   U1090 : OAI22_X1 port map( A1 => n13214, A2 => n11369, B1 => n11386, B2 => 
                           n11368, ZN => n1264);
   U1091 : OAI22_X1 port map( A1 => n13475, A2 => n11369, B1 => n11387, B2 => 
                           n11367, ZN => n1263);
   U1092 : OAI22_X1 port map( A1 => n13215, A2 => n11369, B1 => n11388, B2 => 
                           n11368, ZN => n1262);
   U1093 : OAI22_X1 port map( A1 => n13216, A2 => n11369, B1 => n11389, B2 => 
                           n11367, ZN => n1261);
   U1094 : OAI22_X1 port map( A1 => n13217, A2 => n11369, B1 => n11390, B2 => 
                           n11367, ZN => n1260);
   U1095 : OAI22_X1 port map( A1 => n13218, A2 => n11369, B1 => n11391, B2 => 
                           n11368, ZN => n1259);
   U1096 : OAI22_X1 port map( A1 => n13219, A2 => n11369, B1 => n11392, B2 => 
                           n11367, ZN => n1258);
   U1097 : OAI22_X1 port map( A1 => n13716, A2 => n11369, B1 => n11393, B2 => 
                           n11368, ZN => n1257);
   U1098 : OAI22_X1 port map( A1 => n13220, A2 => n11369, B1 => n11394, B2 => 
                           n11367, ZN => n1256);
   U1099 : OAI22_X1 port map( A1 => n13960, A2 => n11369, B1 => n11395, B2 => 
                           n11368, ZN => n1255);
   U1100 : OAI22_X1 port map( A1 => n13221, A2 => n11369, B1 => n11396, B2 => 
                           n11367, ZN => n1254);
   U1101 : OAI22_X1 port map( A1 => n13222, A2 => n11369, B1 => n11397, B2 => 
                           n11367, ZN => n1253);
   U1102 : OAI22_X1 port map( A1 => n13476, A2 => n11369, B1 => n11398, B2 => 
                           n11367, ZN => n1252);
   U1103 : OAI22_X1 port map( A1 => n13477, A2 => n11369, B1 => n11399, B2 => 
                           n11367, ZN => n1251);
   U1104 : OAI22_X1 port map( A1 => n13717, A2 => n11369, B1 => n11400, B2 => 
                           n11367, ZN => n1250);
   U1105 : OAI22_X1 port map( A1 => n13718, A2 => n11369, B1 => n11401, B2 => 
                           n11367, ZN => n1249);
   U1106 : OAI22_X1 port map( A1 => n13961, A2 => n11369, B1 => n11403, B2 => 
                           n11367, ZN => n1248);
   U1107 : OAI22_X1 port map( A1 => n13719, A2 => n11369, B1 => n11404, B2 => 
                           n11368, ZN => n1247);
   U1108 : OAI22_X1 port map( A1 => n13720, A2 => n11369, B1 => n11405, B2 => 
                           n11368, ZN => n1246);
   U1109 : OAI22_X1 port map( A1 => n13962, A2 => n11369, B1 => n11406, B2 => 
                           n11368, ZN => n1245);
   U1110 : OAI22_X1 port map( A1 => n13963, A2 => n11369, B1 => n11407, B2 => 
                           n11368, ZN => n1244);
   U1111 : OAI22_X1 port map( A1 => n13721, A2 => n11369, B1 => n11408, B2 => 
                           n11368, ZN => n1243);
   U1112 : OAI22_X1 port map( A1 => n13478, A2 => n11369, B1 => n11409, B2 => 
                           n11368, ZN => n1242);
   U1113 : OAI22_X1 port map( A1 => n13722, A2 => n11369, B1 => n11410, B2 => 
                           n11368, ZN => n1241);
   U1114 : OAI22_X1 port map( A1 => n13964, A2 => n11369, B1 => n11411, B2 => 
                           n11368, ZN => n1240);
   U1115 : OAI22_X1 port map( A1 => n13479, A2 => n11369, B1 => n11413, B2 => 
                           n11368, ZN => n1239);
   U1116 : NAND2_X1 port map( A1 => n11370, A2 => n11378, ZN => n11371);
   U1117 : CLKBUF_X1 port map( A => n11371, Z => n11372);
   U1118 : OAI22_X1 port map( A1 => n13497, A2 => n11373, B1 => n11380, B2 => 
                           n11372, ZN => n1238);
   U1119 : OAI22_X1 port map( A1 => n13723, A2 => n11373, B1 => n11381, B2 => 
                           n11371, ZN => n1237);
   U1120 : OAI22_X1 port map( A1 => n13965, A2 => n11373, B1 => n11382, B2 => 
                           n11372, ZN => n1236);
   U1121 : OAI22_X1 port map( A1 => n13724, A2 => n11373, B1 => n11383, B2 => 
                           n11371, ZN => n1235);
   U1122 : OAI22_X1 port map( A1 => n13966, A2 => n11373, B1 => n11384, B2 => 
                           n11372, ZN => n1234);
   U1123 : OAI22_X1 port map( A1 => n13725, A2 => n11373, B1 => n11385, B2 => 
                           n11371, ZN => n1233);
   U1124 : OAI22_X1 port map( A1 => n13726, A2 => n11373, B1 => n11386, B2 => 
                           n11372, ZN => n1232);
   U1125 : OAI22_X1 port map( A1 => n13967, A2 => n11373, B1 => n11387, B2 => 
                           n11371, ZN => n1231);
   U1126 : OAI22_X1 port map( A1 => n13727, A2 => n11373, B1 => n11388, B2 => 
                           n11372, ZN => n1230);
   U1127 : OAI22_X1 port map( A1 => n13968, A2 => n11373, B1 => n11389, B2 => 
                           n11371, ZN => n1229);
   U1128 : OAI22_X1 port map( A1 => n13969, A2 => n11373, B1 => n11390, B2 => 
                           n11371, ZN => n1228);
   U1129 : OAI22_X1 port map( A1 => n13970, A2 => n11373, B1 => n11391, B2 => 
                           n11372, ZN => n1227);
   U1130 : OAI22_X1 port map( A1 => n13971, A2 => n11373, B1 => n11392, B2 => 
                           n11371, ZN => n1226);
   U1131 : OAI22_X1 port map( A1 => n13972, A2 => n11373, B1 => n11393, B2 => 
                           n11372, ZN => n1225);
   U1132 : OAI22_X1 port map( A1 => n13973, A2 => n11373, B1 => n11394, B2 => 
                           n11371, ZN => n1224);
   U1133 : OAI22_X1 port map( A1 => n13728, A2 => n11373, B1 => n11395, B2 => 
                           n11372, ZN => n1223);
   U1134 : OAI22_X1 port map( A1 => n13974, A2 => n11373, B1 => n11396, B2 => 
                           n11371, ZN => n1222);
   U1135 : OAI22_X1 port map( A1 => n13975, A2 => n11373, B1 => n11397, B2 => 
                           n11371, ZN => n1221);
   U1136 : OAI22_X1 port map( A1 => n13976, A2 => n11373, B1 => n11398, B2 => 
                           n11371, ZN => n1220);
   U1137 : OAI22_X1 port map( A1 => n13729, A2 => n11373, B1 => n11399, B2 => 
                           n11371, ZN => n1219);
   U1138 : OAI22_X1 port map( A1 => n13977, A2 => n11373, B1 => n11400, B2 => 
                           n11371, ZN => n1218);
   U1139 : OAI22_X1 port map( A1 => n13978, A2 => n11373, B1 => n11401, B2 => 
                           n11371, ZN => n1217);
   U1140 : OAI22_X1 port map( A1 => n13730, A2 => n11373, B1 => n11403, B2 => 
                           n11371, ZN => n1216);
   U1141 : OAI22_X1 port map( A1 => n13979, A2 => n11373, B1 => n11404, B2 => 
                           n11372, ZN => n1215);
   U1142 : OAI22_X1 port map( A1 => n13980, A2 => n11373, B1 => n11405, B2 => 
                           n11372, ZN => n1214);
   U1143 : OAI22_X1 port map( A1 => n13981, A2 => n11373, B1 => n11406, B2 => 
                           n11372, ZN => n1213);
   U1144 : OAI22_X1 port map( A1 => n13731, A2 => n11373, B1 => n11407, B2 => 
                           n11372, ZN => n1212);
   U1145 : OAI22_X1 port map( A1 => n13982, A2 => n11373, B1 => n11408, B2 => 
                           n11372, ZN => n1211);
   U1146 : OAI22_X1 port map( A1 => n13732, A2 => n11373, B1 => n11409, B2 => 
                           n11372, ZN => n1210);
   U1147 : OAI22_X1 port map( A1 => n13983, A2 => n11373, B1 => n11410, B2 => 
                           n11372, ZN => n1209);
   U1148 : OAI22_X1 port map( A1 => n13984, A2 => n11373, B1 => n11411, B2 => 
                           n11372, ZN => n1208);
   U1149 : OAI22_X1 port map( A1 => n13985, A2 => n11373, B1 => n11413, B2 => 
                           n11372, ZN => n1207);
   U1150 : NAND2_X1 port map( A1 => n11374, A2 => n11378, ZN => n11375);
   U1151 : CLKBUF_X1 port map( A => n11375, Z => n11376);
   U1152 : OAI22_X1 port map( A1 => n13249, A2 => n11377, B1 => n11380, B2 => 
                           n11376, ZN => n1206);
   U1153 : OAI22_X1 port map( A1 => n13733, A2 => n11377, B1 => n11381, B2 => 
                           n11375, ZN => n1205);
   U1154 : OAI22_X1 port map( A1 => n13986, A2 => n11377, B1 => n11382, B2 => 
                           n11376, ZN => n1204);
   U1155 : OAI22_X1 port map( A1 => n13223, A2 => n11377, B1 => n11383, B2 => 
                           n11375, ZN => n1203);
   U1156 : OAI22_X1 port map( A1 => n13224, A2 => n11377, B1 => n11384, B2 => 
                           n11376, ZN => n1202);
   U1157 : OAI22_X1 port map( A1 => n13734, A2 => n11377, B1 => n11385, B2 => 
                           n11375, ZN => n1201);
   U1158 : OAI22_X1 port map( A1 => n13987, A2 => n11377, B1 => n11386, B2 => 
                           n11376, ZN => n1200);
   U1159 : OAI22_X1 port map( A1 => n13225, A2 => n11377, B1 => n11387, B2 => 
                           n11375, ZN => n1199);
   U1160 : OAI22_X1 port map( A1 => n13988, A2 => n11377, B1 => n11388, B2 => 
                           n11376, ZN => n1198);
   U1161 : OAI22_X1 port map( A1 => n13480, A2 => n11377, B1 => n11389, B2 => 
                           n11375, ZN => n1197);
   U1162 : OAI22_X1 port map( A1 => n13735, A2 => n11377, B1 => n11390, B2 => 
                           n11375, ZN => n1196);
   U1163 : OAI22_X1 port map( A1 => n13736, A2 => n11377, B1 => n11391, B2 => 
                           n11376, ZN => n1195);
   U1164 : OAI22_X1 port map( A1 => n13989, A2 => n11377, B1 => n11392, B2 => 
                           n11375, ZN => n1194);
   U1165 : OAI22_X1 port map( A1 => n13990, A2 => n11377, B1 => n11393, B2 => 
                           n11376, ZN => n1193);
   U1166 : OAI22_X1 port map( A1 => n13991, A2 => n11377, B1 => n11394, B2 => 
                           n11375, ZN => n1192);
   U1167 : OAI22_X1 port map( A1 => n13481, A2 => n11377, B1 => n11395, B2 => 
                           n11376, ZN => n1191);
   U1168 : OAI22_X1 port map( A1 => n13992, A2 => n11377, B1 => n11396, B2 => 
                           n11375, ZN => n1190);
   U1169 : OAI22_X1 port map( A1 => n13482, A2 => n11377, B1 => n11397, B2 => 
                           n11375, ZN => n1189);
   U1170 : OAI22_X1 port map( A1 => n13483, A2 => n11377, B1 => n11398, B2 => 
                           n11375, ZN => n1188);
   U1171 : OAI22_X1 port map( A1 => n13226, A2 => n11377, B1 => n11399, B2 => 
                           n11375, ZN => n1187);
   U1172 : OAI22_X1 port map( A1 => n13993, A2 => n11377, B1 => n11400, B2 => 
                           n11375, ZN => n1186);
   U1173 : OAI22_X1 port map( A1 => n13737, A2 => n11377, B1 => n11401, B2 => 
                           n11375, ZN => n1185);
   U1174 : OAI22_X1 port map( A1 => n13994, A2 => n11377, B1 => n11403, B2 => 
                           n11375, ZN => n1184);
   U1175 : OAI22_X1 port map( A1 => n13484, A2 => n11377, B1 => n11404, B2 => 
                           n11376, ZN => n1183);
   U1176 : OAI22_X1 port map( A1 => n13485, A2 => n11377, B1 => n11405, B2 => 
                           n11376, ZN => n1182);
   U1177 : OAI22_X1 port map( A1 => n13227, A2 => n11377, B1 => n11406, B2 => 
                           n11376, ZN => n1181);
   U1178 : OAI22_X1 port map( A1 => n13995, A2 => n11377, B1 => n11407, B2 => 
                           n11376, ZN => n1180);
   U1179 : OAI22_X1 port map( A1 => n13738, A2 => n11377, B1 => n11408, B2 => 
                           n11376, ZN => n1179);
   U1180 : OAI22_X1 port map( A1 => n13228, A2 => n11377, B1 => n11409, B2 => 
                           n11376, ZN => n1178);
   U1181 : OAI22_X1 port map( A1 => n13229, A2 => n11377, B1 => n11410, B2 => 
                           n11376, ZN => n1177);
   U1182 : OAI22_X1 port map( A1 => n13230, A2 => n11377, B1 => n11411, B2 => 
                           n11376, ZN => n1176);
   U1183 : OAI22_X1 port map( A1 => n13739, A2 => n11377, B1 => n11413, B2 => 
                           n11376, ZN => n1175);
   U1184 : NAND2_X1 port map( A1 => n11379, A2 => n11378, ZN => n11402);
   U1185 : CLKBUF_X1 port map( A => n11402, Z => n11412);
   U1186 : OAI22_X1 port map( A1 => n13498, A2 => n11414, B1 => n11380, B2 => 
                           n11412, ZN => n1174);
   U1187 : OAI22_X1 port map( A1 => n13740, A2 => n11414, B1 => n11381, B2 => 
                           n11402, ZN => n1173);
   U1188 : OAI22_X1 port map( A1 => n13996, A2 => n11414, B1 => n11382, B2 => 
                           n11412, ZN => n1172);
   U1189 : OAI22_X1 port map( A1 => n13486, A2 => n11414, B1 => n11383, B2 => 
                           n11402, ZN => n1171);
   U1190 : OAI22_X1 port map( A1 => n13487, A2 => n11414, B1 => n11384, B2 => 
                           n11412, ZN => n1170);
   U1191 : OAI22_X1 port map( A1 => n13997, A2 => n11414, B1 => n11385, B2 => 
                           n11402, ZN => n1169);
   U1192 : OAI22_X1 port map( A1 => n13488, A2 => n11414, B1 => n11386, B2 => 
                           n11412, ZN => n1168);
   U1193 : OAI22_X1 port map( A1 => n13489, A2 => n11414, B1 => n11387, B2 => 
                           n11402, ZN => n1167);
   U1194 : OAI22_X1 port map( A1 => n13231, A2 => n11414, B1 => n11388, B2 => 
                           n11412, ZN => n1166);
   U1195 : OAI22_X1 port map( A1 => n13232, A2 => n11414, B1 => n11389, B2 => 
                           n11402, ZN => n1165);
   U1196 : OAI22_X1 port map( A1 => n13741, A2 => n11414, B1 => n11390, B2 => 
                           n11402, ZN => n1164);
   U1197 : OAI22_X1 port map( A1 => n13998, A2 => n11414, B1 => n11391, B2 => 
                           n11412, ZN => n1163);
   U1198 : OAI22_X1 port map( A1 => n13490, A2 => n11414, B1 => n11392, B2 => 
                           n11402, ZN => n1162);
   U1199 : OAI22_X1 port map( A1 => n13742, A2 => n11414, B1 => n11393, B2 => 
                           n11412, ZN => n1161);
   U1200 : OAI22_X1 port map( A1 => n13233, A2 => n11414, B1 => n11394, B2 => 
                           n11402, ZN => n1160);
   U1201 : OAI22_X1 port map( A1 => n13234, A2 => n11414, B1 => n11395, B2 => 
                           n11412, ZN => n1159);
   U1202 : OAI22_X1 port map( A1 => n13491, A2 => n11414, B1 => n11396, B2 => 
                           n11402, ZN => n1158);
   U1203 : OAI22_X1 port map( A1 => n13235, A2 => n11414, B1 => n11397, B2 => 
                           n11402, ZN => n1157);
   U1204 : OAI22_X1 port map( A1 => n13999, A2 => n11414, B1 => n11398, B2 => 
                           n11402, ZN => n1156);
   U1205 : OAI22_X1 port map( A1 => n13236, A2 => n11414, B1 => n11399, B2 => 
                           n11402, ZN => n1155);
   U1206 : OAI22_X1 port map( A1 => n13237, A2 => n11414, B1 => n11400, B2 => 
                           n11402, ZN => n1154);
   U1207 : OAI22_X1 port map( A1 => n13238, A2 => n11414, B1 => n11401, B2 => 
                           n11402, ZN => n1153);
   U1208 : OAI22_X1 port map( A1 => n13492, A2 => n11414, B1 => n11403, B2 => 
                           n11402, ZN => n1152);
   U1209 : OAI22_X1 port map( A1 => n13239, A2 => n11414, B1 => n11404, B2 => 
                           n11412, ZN => n1151);
   U1210 : OAI22_X1 port map( A1 => n14000, A2 => n11414, B1 => n11405, B2 => 
                           n11412, ZN => n1150);
   U1211 : OAI22_X1 port map( A1 => n14001, A2 => n11414, B1 => n11406, B2 => 
                           n11412, ZN => n1149);
   U1212 : OAI22_X1 port map( A1 => n13240, A2 => n11414, B1 => n11407, B2 => 
                           n11412, ZN => n1148);
   U1213 : OAI22_X1 port map( A1 => n13493, A2 => n11414, B1 => n11408, B2 => 
                           n11412, ZN => n1147);
   U1214 : OAI22_X1 port map( A1 => n14002, A2 => n11414, B1 => n11409, B2 => 
                           n11412, ZN => n1146);
   U1215 : OAI22_X1 port map( A1 => n13494, A2 => n11414, B1 => n11410, B2 => 
                           n11412, ZN => n1145);
   U1216 : OAI22_X1 port map( A1 => n13241, A2 => n11414, B1 => n11411, B2 => 
                           n11412, ZN => n1144);
   U1217 : OAI22_X1 port map( A1 => n13743, A2 => n11414, B1 => n11413, B2 => 
                           n11412, ZN => n1143);
   U1218 : NAND3_X1 port map( A1 => n11229, A2 => ENABLE, A3 => RD2, ZN => 
                           n12196);
   U1219 : INV_X1 port map( A => ADD_RD2(3), ZN => n11443);
   U1220 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n11443, ZN => n11423);
   U1221 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), ZN => n11416);
   U1222 : NAND2_X1 port map( A1 => ADD_RD2(1), A2 => n11416, ZN => n11438);
   U1223 : NOR2_X1 port map( A1 => n11423, A2 => n11438, ZN => n11826);
   U1224 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n11436);
   U1225 : NOR2_X1 port map( A1 => n11423, A2 => n11436, ZN => n12013);
   U1226 : CLKBUF_X1 port map( A => n12013, Z => n12149);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_18_31_port, A2 => n11826, B1 => 
                           REGISTERS_23_31_port, B2 => n12149, ZN => n11420);
   U1228 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n11424)
                           ;
   U1229 : NOR2_X1 port map( A1 => n11424, A2 => n11436, ZN => n12150);
   U1230 : INV_X1 port map( A => ADD_RD2(1), ZN => n11422);
   U1231 : INV_X1 port map( A => ADD_RD2(0), ZN => n11421);
   U1232 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => n11422, A3 => n11421, ZN 
                           => n11431);
   U1233 : NOR2_X1 port map( A1 => n11424, A2 => n11431, ZN => n12163);
   U1234 : CLKBUF_X1 port map( A => n12163, Z => n12119);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_31_31_port, A2 => n12150, B1 => 
                           REGISTERS_28_31_port, B2 => n12119, ZN => n11419);
   U1236 : INV_X1 port map( A => ADD_RD2(2), ZN => n11415);
   U1237 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => n11415,
                           ZN => n11434);
   U1238 : NOR2_X1 port map( A1 => n11424, A2 => n11434, ZN => n11965);
   U1239 : NOR2_X1 port map( A1 => n11423, A2 => n11434, ZN => n12145);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n11965, B1 => 
                           REGISTERS_19_31_port, B2 => n12145, ZN => n11418);
   U1241 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n11422, A3 => n11415, ZN 
                           => n11437);
   U1242 : NOR2_X1 port map( A1 => n11424, A2 => n11437, ZN => n11853);
   U1243 : NAND2_X1 port map( A1 => n11416, A2 => n11422, ZN => n11432);
   U1244 : NOR2_X1 port map( A1 => n11424, A2 => n11432, ZN => n11989);
   U1245 : CLKBUF_X1 port map( A => n11989, Z => n12157);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n11853, B1 => 
                           REGISTERS_24_31_port, B2 => n12157, ZN => n11417);
   U1247 : NAND4_X1 port map( A1 => n11420, A2 => n11419, A3 => n11418, A4 => 
                           n11417, ZN => n11430);
   U1248 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => n11421,
                           ZN => n11435);
   U1249 : NOR2_X1 port map( A1 => n11423, A2 => n11435, ZN => n11970);
   U1250 : NOR2_X1 port map( A1 => n11423, A2 => n11431, ZN => n11900);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n11970, B1 => 
                           REGISTERS_20_31_port, B2 => n11900, ZN => n11428);
   U1252 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => n11422,
                           ZN => n11433);
   U1253 : NOR2_X1 port map( A1 => n11424, A2 => n11433, ZN => n12164);
   U1254 : NOR2_X1 port map( A1 => n11433, A2 => n11423, ZN => n12120);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n12164, B1 => 
                           REGISTERS_21_31_port, B2 => n12120, ZN => n11427);
   U1256 : NOR2_X1 port map( A1 => n11424, A2 => n11438, ZN => n12112);
   U1257 : NOR2_X1 port map( A1 => n11423, A2 => n11432, ZN => n12086);
   U1258 : CLKBUF_X1 port map( A => n12086, Z => n12158);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n12112, B1 => 
                           REGISTERS_16_31_port, B2 => n12158, ZN => n11426);
   U1260 : NOR2_X1 port map( A1 => n11423, A2 => n11437, ZN => n12018);
   U1261 : NOR2_X1 port map( A1 => n11424, A2 => n11435, ZN => n12113);
   U1262 : CLKBUF_X1 port map( A => n12113, Z => n12146);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n12018, B1 => 
                           REGISTERS_30_31_port, B2 => n12146, ZN => n11425);
   U1264 : NAND4_X1 port map( A1 => n11428, A2 => n11427, A3 => n11426, A4 => 
                           n11425, ZN => n11429);
   U1265 : NOR2_X1 port map( A1 => n11430, A2 => n11429, ZN => n11451);
   U1266 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n12144, 
                           ZN => n12193);
   U1267 : CLKBUF_X1 port map( A => n12193, Z => n12010);
   U1268 : INV_X1 port map( A => n11431, ZN => n12077);
   U1269 : CLKBUF_X1 port map( A => n12077, Z => n12183);
   U1270 : INV_X1 port map( A => n11432, ZN => n12127);
   U1271 : CLKBUF_X1 port map( A => n12127, Z => n12134);
   U1272 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_31_port, B1 => 
                           n12134, B2 => REGISTERS_0_31_port, ZN => n11442);
   U1273 : INV_X1 port map( A => n11433, ZN => n12098);
   U1274 : CLKBUF_X1 port map( A => n12098, Z => n11886);
   U1275 : INV_X1 port map( A => n11434, ZN => n12099);
   U1276 : CLKBUF_X1 port map( A => n12099, Z => n11887);
   U1277 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_31_port, B1 => 
                           n11887, B2 => REGISTERS_3_31_port, ZN => n11441);
   U1278 : INV_X1 port map( A => n11435, ZN => n12185);
   U1279 : CLKBUF_X1 port map( A => n12185, Z => n12171);
   U1280 : INV_X1 port map( A => n11436, ZN => n12049);
   U1281 : CLKBUF_X1 port map( A => n12049, Z => n12172);
   U1282 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_31_port, B1 => 
                           n12172, B2 => REGISTERS_7_31_port, ZN => n11440);
   U1283 : INV_X1 port map( A => n11437, ZN => n12054);
   U1284 : CLKBUF_X1 port map( A => n12054, Z => n12181);
   U1285 : INV_X1 port map( A => n11438, ZN => n12182);
   U1286 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_31_port, B1 => 
                           n12182, B2 => REGISTERS_2_31_port, ZN => n11439);
   U1287 : NAND4_X1 port map( A1 => n11442, A2 => n11441, A3 => n11440, A4 => 
                           n11439, ZN => n11449);
   U1288 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n11443, A3 => n12144, ZN 
                           => n12191);
   U1289 : CLKBUF_X1 port map( A => n12191, Z => n12034);
   U1290 : CLKBUF_X1 port map( A => n12182, Z => n12173);
   U1291 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_31_port, B1 => 
                           n12173, B2 => REGISTERS_10_31_port, ZN => n11447);
   U1292 : CLKBUF_X1 port map( A => n12185, Z => n12133);
   U1293 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_31_port, B1 => 
                           n12133, B2 => REGISTERS_14_31_port, ZN => n11446);
   U1294 : CLKBUF_X1 port map( A => n12077, Z => n12097);
   U1295 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_12_31_port, B1 => 
                           n11887, B2 => REGISTERS_11_31_port, ZN => n11445);
   U1296 : CLKBUF_X1 port map( A => n12049, Z => n12178);
   U1297 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_31_port, B1 => 
                           n12178, B2 => REGISTERS_15_31_port, ZN => n11444);
   U1298 : NAND4_X1 port map( A1 => n11447, A2 => n11446, A3 => n11445, A4 => 
                           n11444, ZN => n11448);
   U1299 : AOI22_X1 port map( A1 => n12010, A2 => n11449, B1 => n12034, B2 => 
                           n11448, ZN => n11450);
   U1300 : OAI21_X1 port map( B1 => n12144, B2 => n11451, A => n11450, ZN => 
                           N448);
   U1301 : AOI22_X1 port map( A1 => n11900, A2 => REGISTERS_20_30_port, B1 => 
                           n12086, B2 => REGISTERS_16_30_port, ZN => n11455);
   U1302 : CLKBUF_X1 port map( A => n12150, Z => n12114);
   U1303 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_30_port, B1 => 
                           n12149, B2 => REGISTERS_23_30_port, ZN => n11454);
   U1304 : CLKBUF_X1 port map( A => n12164, Z => n11946);
   U1305 : CLKBUF_X1 port map( A => n11826, Z => n12161);
   U1306 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_30_port, B1 => 
                           n12161, B2 => REGISTERS_18_30_port, ZN => n11453);
   U1307 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_30_port, B1 => 
                           n12112, B2 => REGISTERS_26_30_port, ZN => n11452);
   U1308 : NAND4_X1 port map( A1 => n11455, A2 => n11454, A3 => n11453, A4 => 
                           n11452, ZN => n11461);
   U1309 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_30_port, B1 => 
                           n12119, B2 => REGISTERS_28_30_port, ZN => n11459);
   U1310 : CLKBUF_X1 port map( A => n12018, Z => n12162);
   U1311 : CLKBUF_X1 port map( A => n12145, Z => n11941);
   U1312 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_30_port, B1 => 
                           n11941, B2 => REGISTERS_19_30_port, ZN => n11458);
   U1313 : CLKBUF_X1 port map( A => n11970, Z => n12148);
   U1314 : CLKBUF_X1 port map( A => n11965, Z => n12147);
   U1315 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_30_port, B1 => 
                           n12147, B2 => REGISTERS_27_30_port, ZN => n11457);
   U1316 : CLKBUF_X1 port map( A => n11853, Z => n12159);
   U1317 : AOI22_X1 port map( A1 => n12159, A2 => REGISTERS_25_30_port, B1 => 
                           n12157, B2 => REGISTERS_24_30_port, ZN => n11456);
   U1318 : NAND4_X1 port map( A1 => n11459, A2 => n11458, A3 => n11457, A4 => 
                           n11456, ZN => n11460);
   U1319 : NOR2_X1 port map( A1 => n11461, A2 => n11460, ZN => n11473);
   U1320 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_30_port, B1 => 
                           n12178, B2 => REGISTERS_7_30_port, ZN => n11465);
   U1321 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_30_port, B1 => 
                           n12097, B2 => REGISTERS_4_30_port, ZN => n11464);
   U1322 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_30_port, B1 => 
                           n12173, B2 => REGISTERS_2_30_port, ZN => n11463);
   U1323 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_0_30_port, B1 => 
                           n11887, B2 => REGISTERS_3_30_port, ZN => n11462);
   U1324 : NAND4_X1 port map( A1 => n11465, A2 => n11464, A3 => n11463, A4 => 
                           n11462, ZN => n11471);
   U1325 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_30_port, B1 => 
                           n12178, B2 => REGISTERS_15_30_port, ZN => n11469);
   U1326 : CLKBUF_X1 port map( A => n12182, Z => n12132);
   U1327 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_30_port, B1 => 
                           n11887, B2 => REGISTERS_11_30_port, ZN => n11468);
   U1328 : CLKBUF_X1 port map( A => n12127, Z => n12180);
   U1329 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_30_port, B1 => 
                           n12180, B2 => REGISTERS_8_30_port, ZN => n11467);
   U1330 : CLKBUF_X1 port map( A => n12054, Z => n12135);
   U1331 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_30_port, B1 => 
                           n12135, B2 => REGISTERS_9_30_port, ZN => n11466);
   U1332 : NAND4_X1 port map( A1 => n11469, A2 => n11468, A3 => n11467, A4 => 
                           n11466, ZN => n11470);
   U1333 : AOI22_X1 port map( A1 => n12010, A2 => n11471, B1 => n12034, B2 => 
                           n11470, ZN => n11472);
   U1334 : OAI21_X1 port map( B1 => n12144, B2 => n11473, A => n11472, ZN => 
                           N447);
   U1335 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_29_port, B1 => 
                           n11941, B2 => REGISTERS_19_29_port, ZN => n11477);
   U1336 : AOI22_X1 port map( A1 => n12157, A2 => REGISTERS_24_29_port, B1 => 
                           n11965, B2 => REGISTERS_27_29_port, ZN => n11476);
   U1337 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_29_port, B1 => 
                           n12018, B2 => REGISTERS_17_29_port, ZN => n11475);
   U1338 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_29_port, B1 => 
                           n12013, B2 => REGISTERS_23_29_port, ZN => n11474);
   U1339 : NAND4_X1 port map( A1 => n11477, A2 => n11476, A3 => n11475, A4 => 
                           n11474, ZN => n11483);
   U1340 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_29_port, B1 => 
                           n11900, B2 => REGISTERS_20_29_port, ZN => n11481);
   U1341 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_29_port, B1 => 
                           n12112, B2 => REGISTERS_26_29_port, ZN => n11480);
   U1342 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_29_port, B1 => 
                           n12163, B2 => REGISTERS_28_29_port, ZN => n11479);
   U1343 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_29_port, B1 => 
                           n12159, B2 => REGISTERS_25_29_port, ZN => n11478);
   U1344 : NAND4_X1 port map( A1 => n11481, A2 => n11480, A3 => n11479, A4 => 
                           n11478, ZN => n11482);
   U1345 : NOR2_X1 port map( A1 => n11483, A2 => n11482, ZN => n11495);
   U1346 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_29_port, B1 => 
                           n12180, B2 => REGISTERS_0_29_port, ZN => n11487);
   U1347 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_29_port, B1 => 
                           n12097, B2 => REGISTERS_4_29_port, ZN => n11486);
   U1348 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_29_port, B1 => 
                           n11887, B2 => REGISTERS_3_29_port, ZN => n11485);
   U1349 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_29_port, B1 => 
                           n12178, B2 => REGISTERS_7_29_port, ZN => n11484);
   U1350 : NAND4_X1 port map( A1 => n11487, A2 => n11486, A3 => n11485, A4 => 
                           n11484, ZN => n11493);
   U1351 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_9_29_port, B1 => 
                           n11887, B2 => REGISTERS_11_29_port, ZN => n11491);
   U1352 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_29_port, B1 => 
                           n12180, B2 => REGISTERS_8_29_port, ZN => n11490);
   U1353 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_14_29_port, B1 => 
                           n12097, B2 => REGISTERS_12_29_port, ZN => n11489);
   U1354 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_29_port, B1 => 
                           n12178, B2 => REGISTERS_15_29_port, ZN => n11488);
   U1355 : NAND4_X1 port map( A1 => n11491, A2 => n11490, A3 => n11489, A4 => 
                           n11488, ZN => n11492);
   U1356 : AOI22_X1 port map( A1 => n12010, A2 => n11493, B1 => n12034, B2 => 
                           n11492, ZN => n11494);
   U1357 : OAI21_X1 port map( B1 => n12144, B2 => n11495, A => n11494, ZN => 
                           N446);
   U1358 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_28_port, B1 => 
                           n12114, B2 => REGISTERS_31_28_port, ZN => n11499);
   U1359 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_28_port, B1 => 
                           n12113, B2 => REGISTERS_30_28_port, ZN => n11498);
   U1360 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_28_port, B1 => 
                           n11989, B2 => REGISTERS_24_28_port, ZN => n11497);
   U1361 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_28_port, B1 => 
                           n11941, B2 => REGISTERS_19_28_port, ZN => n11496);
   U1362 : NAND4_X1 port map( A1 => n11499, A2 => n11498, A3 => n11497, A4 => 
                           n11496, ZN => n11505);
   U1363 : AOI22_X1 port map( A1 => n11970, A2 => REGISTERS_22_28_port, B1 => 
                           n11965, B2 => REGISTERS_27_28_port, ZN => n11503);
   U1364 : CLKBUF_X1 port map( A => n11900, Z => n12152);
   U1365 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_28_port, B1 => 
                           n11826, B2 => REGISTERS_18_28_port, ZN => n11502);
   U1366 : AOI22_X1 port map( A1 => n12018, A2 => REGISTERS_17_28_port, B1 => 
                           n11853, B2 => REGISTERS_25_28_port, ZN => n11501);
   U1367 : CLKBUF_X1 port map( A => n12112, Z => n12151);
   U1368 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_28_port, B1 => 
                           n12013, B2 => REGISTERS_23_28_port, ZN => n11500);
   U1369 : NAND4_X1 port map( A1 => n11503, A2 => n11502, A3 => n11501, A4 => 
                           n11500, ZN => n11504);
   U1370 : NOR2_X1 port map( A1 => n11505, A2 => n11504, ZN => n11517);
   U1371 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_4_28_port, B1 => 
                           n12135, B2 => REGISTERS_1_28_port, ZN => n11509);
   U1372 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_0_28_port, B1 => 
                           n11887, B2 => REGISTERS_3_28_port, ZN => n11508);
   U1373 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_28_port, B1 => 
                           n12049, B2 => REGISTERS_7_28_port, ZN => n11507);
   U1374 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_28_port, B1 => 
                           n12173, B2 => REGISTERS_2_28_port, ZN => n11506);
   U1375 : NAND4_X1 port map( A1 => n11509, A2 => n11508, A3 => n11507, A4 => 
                           n11506, ZN => n11515);
   U1376 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_9_28_port, B1 => 
                           n11887, B2 => REGISTERS_11_28_port, ZN => n11513);
   U1377 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_28_port, B1 => 
                           n12178, B2 => REGISTERS_15_28_port, ZN => n11512);
   U1378 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_28_port, B1 => 
                           n12173, B2 => REGISTERS_10_28_port, ZN => n11511);
   U1379 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_28_port, B1 => 
                           n12180, B2 => REGISTERS_8_28_port, ZN => n11510);
   U1380 : NAND4_X1 port map( A1 => n11513, A2 => n11512, A3 => n11511, A4 => 
                           n11510, ZN => n11514);
   U1381 : AOI22_X1 port map( A1 => n12010, A2 => n11515, B1 => n12034, B2 => 
                           n11514, ZN => n11516);
   U1382 : OAI21_X1 port map( B1 => n12144, B2 => n11517, A => n11516, ZN => 
                           N445);
   U1383 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_27_port, B1 => 
                           n11853, B2 => REGISTERS_25_27_port, ZN => n11521);
   U1384 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_27_port, B1 => 
                           n12150, B2 => REGISTERS_31_27_port, ZN => n11520);
   U1385 : AOI22_X1 port map( A1 => n11900, A2 => REGISTERS_20_27_port, B1 => 
                           n12113, B2 => REGISTERS_30_27_port, ZN => n11519);
   U1386 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_27_port, B1 => 
                           n11941, B2 => REGISTERS_19_27_port, ZN => n11518);
   U1387 : NAND4_X1 port map( A1 => n11521, A2 => n11520, A3 => n11519, A4 => 
                           n11518, ZN => n11527);
   U1388 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_27_port, B1 => 
                           n11965, B2 => REGISTERS_27_27_port, ZN => n11525);
   U1389 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_27_port, B1 => 
                           n11989, B2 => REGISTERS_24_27_port, ZN => n11524);
   U1390 : AOI22_X1 port map( A1 => n11970, A2 => REGISTERS_22_27_port, B1 => 
                           n12013, B2 => REGISTERS_23_27_port, ZN => n11523);
   U1391 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_27_port, B1 => 
                           n12163, B2 => REGISTERS_28_27_port, ZN => n11522);
   U1392 : NAND4_X1 port map( A1 => n11525, A2 => n11524, A3 => n11523, A4 => 
                           n11522, ZN => n11526);
   U1393 : NOR2_X1 port map( A1 => n11527, A2 => n11526, ZN => n11539);
   U1394 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_27_port, B1 => 
                           n12173, B2 => REGISTERS_2_27_port, ZN => n11531);
   U1395 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_27_port, B1 => 
                           n12049, B2 => REGISTERS_7_27_port, ZN => n11530);
   U1396 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_4_27_port, B1 => 
                           n11887, B2 => REGISTERS_3_27_port, ZN => n11529);
   U1397 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_27_port, B1 => 
                           n12180, B2 => REGISTERS_0_27_port, ZN => n11528);
   U1398 : NAND4_X1 port map( A1 => n11531, A2 => n11530, A3 => n11529, A4 => 
                           n11528, ZN => n11537);
   U1399 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_12_27_port, B1 => 
                           n12182, B2 => REGISTERS_10_27_port, ZN => n11535);
   U1400 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_27_port, B1 => 
                           n11887, B2 => REGISTERS_11_27_port, ZN => n11534);
   U1401 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_27_port, B1 => 
                           n12178, B2 => REGISTERS_15_27_port, ZN => n11533);
   U1402 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_27_port, B1 => 
                           n12054, B2 => REGISTERS_9_27_port, ZN => n11532);
   U1403 : NAND4_X1 port map( A1 => n11535, A2 => n11534, A3 => n11533, A4 => 
                           n11532, ZN => n11536);
   U1404 : AOI22_X1 port map( A1 => n12010, A2 => n11537, B1 => n12034, B2 => 
                           n11536, ZN => n11538);
   U1405 : OAI21_X1 port map( B1 => n12144, B2 => n11539, A => n11538, ZN => 
                           N444);
   U1406 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_26_port, B1 => 
                           n11965, B2 => REGISTERS_27_26_port, ZN => n11543);
   U1407 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_26_port, B1 => 
                           n11900, B2 => REGISTERS_20_26_port, ZN => n11542);
   U1408 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_26_port, B1 => 
                           n11826, B2 => REGISTERS_18_26_port, ZN => n11541);
   U1409 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_26_port, B1 => 
                           n11853, B2 => REGISTERS_25_26_port, ZN => n11540);
   U1410 : NAND4_X1 port map( A1 => n11543, A2 => n11542, A3 => n11541, A4 => 
                           n11540, ZN => n11549);
   U1411 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_26_port, B1 => 
                           n11941, B2 => REGISTERS_19_26_port, ZN => n11547);
   U1412 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_26_port, B1 => 
                           n12158, B2 => REGISTERS_16_26_port, ZN => n11546);
   U1413 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_26_port, B1 => 
                           n12013, B2 => REGISTERS_23_26_port, ZN => n11545);
   U1414 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_26_port, B1 => 
                           n11989, B2 => REGISTERS_24_26_port, ZN => n11544);
   U1415 : NAND4_X1 port map( A1 => n11547, A2 => n11546, A3 => n11545, A4 => 
                           n11544, ZN => n11548);
   U1416 : NOR2_X1 port map( A1 => n11549, A2 => n11548, ZN => n11561);
   U1417 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_26_port, B1 => 
                           n12049, B2 => REGISTERS_7_26_port, ZN => n11553);
   U1418 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_26_port, B1 => 
                           n12127, B2 => REGISTERS_0_26_port, ZN => n11552);
   U1419 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_26_port, B1 => 
                           n11887, B2 => REGISTERS_3_26_port, ZN => n11551);
   U1420 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_26_port, B1 => 
                           n12133, B2 => REGISTERS_6_26_port, ZN => n11550);
   U1421 : NAND4_X1 port map( A1 => n11553, A2 => n11552, A3 => n11551, A4 => 
                           n11550, ZN => n11559);
   U1422 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_26_port, B1 => 
                           n11887, B2 => REGISTERS_11_26_port, ZN => n11557);
   U1423 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_26_port, B1 => 
                           n12180, B2 => REGISTERS_8_26_port, ZN => n11556);
   U1424 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_26_port, B1 => 
                           n12178, B2 => REGISTERS_15_26_port, ZN => n11555);
   U1425 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_26_port, B1 => 
                           n12173, B2 => REGISTERS_10_26_port, ZN => n11554);
   U1426 : NAND4_X1 port map( A1 => n11557, A2 => n11556, A3 => n11555, A4 => 
                           n11554, ZN => n11558);
   U1427 : AOI22_X1 port map( A1 => n12010, A2 => n11559, B1 => n12034, B2 => 
                           n11558, ZN => n11560);
   U1428 : OAI21_X1 port map( B1 => n12144, B2 => n11561, A => n11560, ZN => 
                           N443);
   U1429 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_25_port, B1 => 
                           n12086, B2 => REGISTERS_16_25_port, ZN => n11565);
   U1430 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_25_port, B1 => 
                           n12150, B2 => REGISTERS_31_25_port, ZN => n11564);
   U1431 : AOI22_X1 port map( A1 => n11970, A2 => REGISTERS_22_25_port, B1 => 
                           n11900, B2 => REGISTERS_20_25_port, ZN => n11563);
   U1432 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_25_port, B1 => 
                           n12163, B2 => REGISTERS_28_25_port, ZN => n11562);
   U1433 : NAND4_X1 port map( A1 => n11565, A2 => n11564, A3 => n11563, A4 => 
                           n11562, ZN => n11571);
   U1434 : AOI22_X1 port map( A1 => n11965, A2 => REGISTERS_27_25_port, B1 => 
                           n11941, B2 => REGISTERS_19_25_port, ZN => n11569);
   U1435 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_25_port, B1 => 
                           n12013, B2 => REGISTERS_23_25_port, ZN => n11568);
   U1436 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_25_port, B1 => 
                           n11853, B2 => REGISTERS_25_25_port, ZN => n11567);
   U1437 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_25_port, B1 => 
                           n11989, B2 => REGISTERS_24_25_port, ZN => n11566);
   U1438 : NAND4_X1 port map( A1 => n11569, A2 => n11568, A3 => n11567, A4 => 
                           n11566, ZN => n11570);
   U1439 : NOR2_X1 port map( A1 => n11571, A2 => n11570, ZN => n11583);
   U1440 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_25_port, B1 => 
                           n12182, B2 => REGISTERS_2_25_port, ZN => n11575);
   U1441 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_25_port, B1 => 
                           n12049, B2 => REGISTERS_7_25_port, ZN => n11574);
   U1442 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_4_25_port, B1 => 
                           n11887, B2 => REGISTERS_3_25_port, ZN => n11573);
   U1443 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_6_25_port, B1 => 
                           n12127, B2 => REGISTERS_0_25_port, ZN => n11572);
   U1444 : NAND4_X1 port map( A1 => n11575, A2 => n11574, A3 => n11573, A4 => 
                           n11572, ZN => n11581);
   U1445 : CLKBUF_X1 port map( A => n12098, Z => n12179);
   U1446 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_25_port, B1 => 
                           n12077, B2 => REGISTERS_12_25_port, ZN => n11579);
   U1447 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_25_port, B1 => 
                           n12173, B2 => REGISTERS_10_25_port, ZN => n11578);
   U1448 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_25_port, B1 => 
                           n12178, B2 => REGISTERS_15_25_port, ZN => n11577);
   U1449 : CLKBUF_X1 port map( A => n12099, Z => n12184);
   U1450 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_9_25_port, B1 => 
                           n12184, B2 => REGISTERS_11_25_port, ZN => n11576);
   U1451 : NAND4_X1 port map( A1 => n11579, A2 => n11578, A3 => n11577, A4 => 
                           n11576, ZN => n11580);
   U1452 : AOI22_X1 port map( A1 => n12010, A2 => n11581, B1 => n12034, B2 => 
                           n11580, ZN => n11582);
   U1453 : OAI21_X1 port map( B1 => n12144, B2 => n11583, A => n11582, ZN => 
                           N442);
   U1454 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_24_port, B1 => 
                           n11826, B2 => REGISTERS_18_24_port, ZN => n11587);
   U1455 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_24_port, B1 => 
                           n11853, B2 => REGISTERS_25_24_port, ZN => n11586);
   U1456 : CLKBUF_X1 port map( A => n12120, Z => n12160);
   U1457 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_24_port, B1 => 
                           n11989, B2 => REGISTERS_24_24_port, ZN => n11585);
   U1458 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_24_port, B1 => 
                           n12113, B2 => REGISTERS_30_24_port, ZN => n11584);
   U1459 : NAND4_X1 port map( A1 => n11587, A2 => n11586, A3 => n11585, A4 => 
                           n11584, ZN => n11593);
   U1460 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_24_port, B1 => 
                           n11941, B2 => REGISTERS_19_24_port, ZN => n11591);
   U1461 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_24_port, B1 => 
                           n12163, B2 => REGISTERS_28_24_port, ZN => n11590);
   U1462 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_24_port, B1 => 
                           n12150, B2 => REGISTERS_31_24_port, ZN => n11589);
   U1463 : AOI22_X1 port map( A1 => n12149, A2 => REGISTERS_23_24_port, B1 => 
                           n11965, B2 => REGISTERS_27_24_port, ZN => n11588);
   U1464 : NAND4_X1 port map( A1 => n11591, A2 => n11590, A3 => n11589, A4 => 
                           n11588, ZN => n11592);
   U1465 : NOR2_X1 port map( A1 => n11593, A2 => n11592, ZN => n11605);
   U1466 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_24_port, B1 => 
                           n12077, B2 => REGISTERS_4_24_port, ZN => n11597);
   U1467 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_24_port, B1 => 
                           n12180, B2 => REGISTERS_0_24_port, ZN => n11596);
   U1468 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_24_port, B1 => 
                           n12049, B2 => REGISTERS_7_24_port, ZN => n11595);
   U1469 : AOI22_X1 port map( A1 => n12182, A2 => REGISTERS_2_24_port, B1 => 
                           n12099, B2 => REGISTERS_3_24_port, ZN => n11594);
   U1470 : NAND4_X1 port map( A1 => n11597, A2 => n11596, A3 => n11595, A4 => 
                           n11594, ZN => n11603);
   U1471 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_24_port, B1 => 
                           n12127, B2 => REGISTERS_8_24_port, ZN => n11601);
   U1472 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_24_port, B1 => 
                           n12135, B2 => REGISTERS_9_24_port, ZN => n11600);
   U1473 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_24_port, B1 => 
                           n12178, B2 => REGISTERS_15_24_port, ZN => n11599);
   U1474 : AOI22_X1 port map( A1 => n12173, A2 => REGISTERS_10_24_port, B1 => 
                           n11887, B2 => REGISTERS_11_24_port, ZN => n11598);
   U1475 : NAND4_X1 port map( A1 => n11601, A2 => n11600, A3 => n11599, A4 => 
                           n11598, ZN => n11602);
   U1476 : AOI22_X1 port map( A1 => n12010, A2 => n11603, B1 => n12034, B2 => 
                           n11602, ZN => n11604);
   U1477 : OAI21_X1 port map( B1 => n12144, B2 => n11605, A => n11604, ZN => 
                           N441);
   U1478 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_23_port, B1 => 
                           n12150, B2 => REGISTERS_31_23_port, ZN => n11609);
   U1479 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_23_port, B1 => 
                           n12013, B2 => REGISTERS_23_23_port, ZN => n11608);
   U1480 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_23_port, B1 => 
                           n12119, B2 => REGISTERS_28_23_port, ZN => n11607);
   U1481 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_23_port, B1 => 
                           n11989, B2 => REGISTERS_24_23_port, ZN => n11606);
   U1482 : NAND4_X1 port map( A1 => n11609, A2 => n11608, A3 => n11607, A4 => 
                           n11606, ZN => n11615);
   U1483 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_23_port, B1 => 
                           n11853, B2 => REGISTERS_25_23_port, ZN => n11613);
   U1484 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_23_port, B1 => 
                           n12158, B2 => REGISTERS_16_23_port, ZN => n11612);
   U1485 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_23_port, B1 => 
                           n11941, B2 => REGISTERS_19_23_port, ZN => n11611);
   U1486 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_23_port, B1 => 
                           n11965, B2 => REGISTERS_27_23_port, ZN => n11610);
   U1487 : NAND4_X1 port map( A1 => n11613, A2 => n11612, A3 => n11611, A4 => 
                           n11610, ZN => n11614);
   U1488 : NOR2_X1 port map( A1 => n11615, A2 => n11614, ZN => n11627);
   U1489 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_0_23_port, B1 => 
                           n12184, B2 => REGISTERS_3_23_port, ZN => n11619);
   U1490 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_4_23_port, B1 => 
                           n12049, B2 => REGISTERS_7_23_port, ZN => n11618);
   U1491 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_23_port, B1 => 
                           n12182, B2 => REGISTERS_2_23_port, ZN => n11617);
   U1492 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_23_port, B1 => 
                           n12054, B2 => REGISTERS_1_23_port, ZN => n11616);
   U1493 : NAND4_X1 port map( A1 => n11619, A2 => n11618, A3 => n11617, A4 => 
                           n11616, ZN => n11625);
   U1494 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_23_port, B1 => 
                           n12049, B2 => REGISTERS_15_23_port, ZN => n11623);
   U1495 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_14_23_port, B1 => 
                           n12173, B2 => REGISTERS_10_23_port, ZN => n11622);
   U1496 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_23_port, B1 => 
                           n12099, B2 => REGISTERS_11_23_port, ZN => n11621);
   U1497 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_23_port, B1 => 
                           n12181, B2 => REGISTERS_9_23_port, ZN => n11620);
   U1498 : NAND4_X1 port map( A1 => n11623, A2 => n11622, A3 => n11621, A4 => 
                           n11620, ZN => n11624);
   U1499 : AOI22_X1 port map( A1 => n12010, A2 => n11625, B1 => n12034, B2 => 
                           n11624, ZN => n11626);
   U1500 : OAI21_X1 port map( B1 => n12196, B2 => n11627, A => n11626, ZN => 
                           N440);
   U1501 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_22_port, B1 => 
                           n12013, B2 => REGISTERS_23_22_port, ZN => n11631);
   U1502 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_22_port, B1 => 
                           n12150, B2 => REGISTERS_31_22_port, ZN => n11630);
   U1503 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_22_port, B1 => 
                           n12163, B2 => REGISTERS_28_22_port, ZN => n11629);
   U1504 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_22_port, B1 => 
                           n11826, B2 => REGISTERS_18_22_port, ZN => n11628);
   U1505 : NAND4_X1 port map( A1 => n11631, A2 => n11630, A3 => n11629, A4 => 
                           n11628, ZN => n11637);
   U1506 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_22_port, B1 => 
                           n12146, B2 => REGISTERS_30_22_port, ZN => n11635);
   U1507 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_22_port, B1 => 
                           n11941, B2 => REGISTERS_19_22_port, ZN => n11634);
   U1508 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_22_port, B1 => 
                           n11853, B2 => REGISTERS_25_22_port, ZN => n11633);
   U1509 : AOI22_X1 port map( A1 => n11989, A2 => REGISTERS_24_22_port, B1 => 
                           n11965, B2 => REGISTERS_27_22_port, ZN => n11632);
   U1510 : NAND4_X1 port map( A1 => n11635, A2 => n11634, A3 => n11633, A4 => 
                           n11632, ZN => n11636);
   U1511 : NOR2_X1 port map( A1 => n11637, A2 => n11636, ZN => n11649);
   U1512 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_4_22_port, B1 => 
                           n12182, B2 => REGISTERS_2_22_port, ZN => n11641);
   U1513 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_22_port, B1 => 
                           n12178, B2 => REGISTERS_7_22_port, ZN => n11640);
   U1514 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_22_port, B1 => 
                           n12180, B2 => REGISTERS_0_22_port, ZN => n11639);
   U1515 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_6_22_port, B1 => 
                           n11887, B2 => REGISTERS_3_22_port, ZN => n11638);
   U1516 : NAND4_X1 port map( A1 => n11641, A2 => n11640, A3 => n11639, A4 => 
                           n11638, ZN => n11647);
   U1517 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_22_port, B1 => 
                           n12049, B2 => REGISTERS_15_22_port, ZN => n11645);
   U1518 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_22_port, B1 => 
                           n12135, B2 => REGISTERS_9_22_port, ZN => n11644);
   U1519 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_22_port, B1 => 
                           n12184, B2 => REGISTERS_11_22_port, ZN => n11643);
   U1520 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_14_22_port, B1 => 
                           n12173, B2 => REGISTERS_10_22_port, ZN => n11642);
   U1521 : NAND4_X1 port map( A1 => n11645, A2 => n11644, A3 => n11643, A4 => 
                           n11642, ZN => n11646);
   U1522 : AOI22_X1 port map( A1 => n12010, A2 => n11647, B1 => n12034, B2 => 
                           n11646, ZN => n11648);
   U1523 : OAI21_X1 port map( B1 => n12196, B2 => n11649, A => n11648, ZN => 
                           N439);
   U1524 : AOI22_X1 port map( A1 => n12113, A2 => REGISTERS_30_21_port, B1 => 
                           n12013, B2 => REGISTERS_23_21_port, ZN => n11653);
   U1525 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_21_port, B1 => 
                           n11853, B2 => REGISTERS_25_21_port, ZN => n11652);
   U1526 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_21_port, B1 => 
                           n11965, B2 => REGISTERS_27_21_port, ZN => n11651);
   U1527 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_21_port, B1 => 
                           n12145, B2 => REGISTERS_19_21_port, ZN => n11650);
   U1528 : NAND4_X1 port map( A1 => n11653, A2 => n11652, A3 => n11651, A4 => 
                           n11650, ZN => n11659);
   U1529 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_21_port, B1 => 
                           n11826, B2 => REGISTERS_18_21_port, ZN => n11657);
   U1530 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_21_port, B1 => 
                           n11989, B2 => REGISTERS_24_21_port, ZN => n11656);
   U1531 : AOI22_X1 port map( A1 => n12086, A2 => REGISTERS_16_21_port, B1 => 
                           n12163, B2 => REGISTERS_28_21_port, ZN => n11655);
   U1532 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_21_port, B1 => 
                           n12018, B2 => REGISTERS_17_21_port, ZN => n11654);
   U1533 : NAND4_X1 port map( A1 => n11657, A2 => n11656, A3 => n11655, A4 => 
                           n11654, ZN => n11658);
   U1534 : NOR2_X1 port map( A1 => n11659, A2 => n11658, ZN => n11671);
   U1535 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_21_port, B1 => 
                           n12097, B2 => REGISTERS_4_21_port, ZN => n11663);
   U1536 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_21_port, B1 => 
                           n12099, B2 => REGISTERS_3_21_port, ZN => n11662);
   U1537 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_21_port, B1 => 
                           n12127, B2 => REGISTERS_0_21_port, ZN => n11661);
   U1538 : AOI22_X1 port map( A1 => n12173, A2 => REGISTERS_2_21_port, B1 => 
                           n12178, B2 => REGISTERS_7_21_port, ZN => n11660);
   U1539 : NAND4_X1 port map( A1 => n11663, A2 => n11662, A3 => n11661, A4 => 
                           n11660, ZN => n11669);
   U1540 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_21_port, B1 => 
                           n12180, B2 => REGISTERS_8_21_port, ZN => n11667);
   U1541 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_21_port, B1 => 
                           n12182, B2 => REGISTERS_10_21_port, ZN => n11666);
   U1542 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_15_21_port, B1 => 
                           n11887, B2 => REGISTERS_11_21_port, ZN => n11665);
   U1543 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_21_port, B1 => 
                           n12181, B2 => REGISTERS_9_21_port, ZN => n11664);
   U1544 : NAND4_X1 port map( A1 => n11667, A2 => n11666, A3 => n11665, A4 => 
                           n11664, ZN => n11668);
   U1545 : AOI22_X1 port map( A1 => n12010, A2 => n11669, B1 => n12034, B2 => 
                           n11668, ZN => n11670);
   U1546 : OAI21_X1 port map( B1 => n12196, B2 => n11671, A => n11670, ZN => 
                           N438);
   U1547 : AOI22_X1 port map( A1 => n12113, A2 => REGISTERS_30_20_port, B1 => 
                           n12159, B2 => REGISTERS_25_20_port, ZN => n11675);
   U1548 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_20_port, B1 => 
                           n11970, B2 => REGISTERS_22_20_port, ZN => n11674);
   U1549 : AOI22_X1 port map( A1 => n12086, A2 => REGISTERS_16_20_port, B1 => 
                           n12163, B2 => REGISTERS_28_20_port, ZN => n11673);
   U1550 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_20_port, B1 => 
                           n12149, B2 => REGISTERS_23_20_port, ZN => n11672);
   U1551 : NAND4_X1 port map( A1 => n11675, A2 => n11674, A3 => n11673, A4 => 
                           n11672, ZN => n11681);
   U1552 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_20_port, B1 => 
                           n11826, B2 => REGISTERS_18_20_port, ZN => n11679);
   U1553 : AOI22_X1 port map( A1 => n12147, A2 => REGISTERS_27_20_port, B1 => 
                           n12145, B2 => REGISTERS_19_20_port, ZN => n11678);
   U1554 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_20_port, B1 => 
                           n12112, B2 => REGISTERS_26_20_port, ZN => n11677);
   U1555 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_20_port, B1 => 
                           n11989, B2 => REGISTERS_24_20_port, ZN => n11676);
   U1556 : NAND4_X1 port map( A1 => n11679, A2 => n11678, A3 => n11677, A4 => 
                           n11676, ZN => n11680);
   U1557 : NOR2_X1 port map( A1 => n11681, A2 => n11680, ZN => n11693);
   U1558 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_20_port, B1 => 
                           n12127, B2 => REGISTERS_0_20_port, ZN => n11685);
   U1559 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_20_port, B1 => 
                           n12184, B2 => REGISTERS_3_20_port, ZN => n11684);
   U1560 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_6_20_port, B1 => 
                           n12173, B2 => REGISTERS_2_20_port, ZN => n11683);
   U1561 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_4_20_port, B1 => 
                           n12049, B2 => REGISTERS_7_20_port, ZN => n11682);
   U1562 : NAND4_X1 port map( A1 => n11685, A2 => n11684, A3 => n11683, A4 => 
                           n11682, ZN => n11691);
   U1563 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_20_port, B1 => 
                           n12180, B2 => REGISTERS_8_20_port, ZN => n11689);
   U1564 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_9_20_port, B1 => 
                           n12182, B2 => REGISTERS_10_20_port, ZN => n11688);
   U1565 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_20_port, B1 => 
                           n12099, B2 => REGISTERS_11_20_port, ZN => n11687);
   U1566 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_20_port, B1 => 
                           n12178, B2 => REGISTERS_15_20_port, ZN => n11686);
   U1567 : NAND4_X1 port map( A1 => n11689, A2 => n11688, A3 => n11687, A4 => 
                           n11686, ZN => n11690);
   U1568 : AOI22_X1 port map( A1 => n12010, A2 => n11691, B1 => n12191, B2 => 
                           n11690, ZN => n11692);
   U1569 : OAI21_X1 port map( B1 => n12196, B2 => n11693, A => n11692, ZN => 
                           N437);
   U1570 : AOI22_X1 port map( A1 => n12159, A2 => REGISTERS_25_19_port, B1 => 
                           n12147, B2 => REGISTERS_27_19_port, ZN => n11697);
   U1571 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_19_port, B1 => 
                           n12119, B2 => REGISTERS_28_19_port, ZN => n11696);
   U1572 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_19_port, B1 => 
                           n12158, B2 => REGISTERS_16_19_port, ZN => n11695);
   U1573 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_19_port, B1 => 
                           n11826, B2 => REGISTERS_18_19_port, ZN => n11694);
   U1574 : NAND4_X1 port map( A1 => n11697, A2 => n11696, A3 => n11695, A4 => 
                           n11694, ZN => n11703);
   U1575 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_19_port, B1 => 
                           n12150, B2 => REGISTERS_31_19_port, ZN => n11701);
   U1576 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_19_port, B1 => 
                           n12149, B2 => REGISTERS_23_19_port, ZN => n11700);
   U1577 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_19_port, B1 => 
                           n12157, B2 => REGISTERS_24_19_port, ZN => n11699);
   U1578 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_19_port, B1 => 
                           n11941, B2 => REGISTERS_19_19_port, ZN => n11698);
   U1579 : NAND4_X1 port map( A1 => n11701, A2 => n11700, A3 => n11699, A4 => 
                           n11698, ZN => n11702);
   U1580 : NOR2_X1 port map( A1 => n11703, A2 => n11702, ZN => n11715);
   U1581 : CLKBUF_X1 port map( A => n12193, Z => n12036);
   U1582 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_19_port, B1 => 
                           n12077, B2 => REGISTERS_4_19_port, ZN => n11707);
   U1583 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_19_port, B1 => 
                           n12127, B2 => REGISTERS_0_19_port, ZN => n11706);
   U1584 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_19_port, B1 => 
                           n12049, B2 => REGISTERS_7_19_port, ZN => n11705);
   U1585 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_19_port, B1 => 
                           n11887, B2 => REGISTERS_3_19_port, ZN => n11704);
   U1586 : NAND4_X1 port map( A1 => n11707, A2 => n11706, A3 => n11705, A4 => 
                           n11704, ZN => n11713);
   U1587 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_19_port, B1 => 
                           n12182, B2 => REGISTERS_10_19_port, ZN => n11711);
   U1588 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_19_port, B1 => 
                           n12127, B2 => REGISTERS_8_19_port, ZN => n11710);
   U1589 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_15_19_port, B1 => 
                           n12184, B2 => REGISTERS_11_19_port, ZN => n11709);
   U1590 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_19_port, B1 => 
                           n12183, B2 => REGISTERS_12_19_port, ZN => n11708);
   U1591 : NAND4_X1 port map( A1 => n11711, A2 => n11710, A3 => n11709, A4 => 
                           n11708, ZN => n11712);
   U1592 : AOI22_X1 port map( A1 => n12036, A2 => n11713, B1 => n12034, B2 => 
                           n11712, ZN => n11714);
   U1593 : OAI21_X1 port map( B1 => n12196, B2 => n11715, A => n11714, ZN => 
                           N436);
   U1594 : AOI22_X1 port map( A1 => n12163, A2 => REGISTERS_28_18_port, B1 => 
                           n11826, B2 => REGISTERS_18_18_port, ZN => n11719);
   U1595 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_18_port, B1 => 
                           n12159, B2 => REGISTERS_25_18_port, ZN => n11718);
   U1596 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_18_port, B1 => 
                           n12149, B2 => REGISTERS_23_18_port, ZN => n11717);
   U1597 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_18_port, B1 => 
                           n12147, B2 => REGISTERS_27_18_port, ZN => n11716);
   U1598 : NAND4_X1 port map( A1 => n11719, A2 => n11718, A3 => n11717, A4 => 
                           n11716, ZN => n11725);
   U1599 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_18_port, B1 => 
                           n11941, B2 => REGISTERS_19_18_port, ZN => n11723);
   U1600 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_18_port, B1 => 
                           n11900, B2 => REGISTERS_20_18_port, ZN => n11722);
   U1601 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_18_port, B1 => 
                           n12158, B2 => REGISTERS_16_18_port, ZN => n11721);
   U1602 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_18_port, B1 => 
                           n12157, B2 => REGISTERS_24_18_port, ZN => n11720);
   U1603 : NAND4_X1 port map( A1 => n11723, A2 => n11722, A3 => n11721, A4 => 
                           n11720, ZN => n11724);
   U1604 : NOR2_X1 port map( A1 => n11725, A2 => n11724, ZN => n11737);
   U1605 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_18_port, B1 => 
                           n12099, B2 => REGISTERS_3_18_port, ZN => n11729);
   U1606 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_4_18_port, B1 => 
                           n12049, B2 => REGISTERS_7_18_port, ZN => n11728);
   U1607 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_6_18_port, B1 => 
                           n12173, B2 => REGISTERS_2_18_port, ZN => n11727);
   U1608 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_18_port, B1 => 
                           n12180, B2 => REGISTERS_0_18_port, ZN => n11726);
   U1609 : NAND4_X1 port map( A1 => n11729, A2 => n11728, A3 => n11727, A4 => 
                           n11726, ZN => n11735);
   U1610 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_15_18_port, B1 => 
                           n11887, B2 => REGISTERS_11_18_port, ZN => n11733);
   U1611 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_18_port, B1 => 
                           n12127, B2 => REGISTERS_8_18_port, ZN => n11732);
   U1612 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_12_18_port, B1 => 
                           n12054, B2 => REGISTERS_9_18_port, ZN => n11731);
   U1613 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_18_port, B1 => 
                           n12182, B2 => REGISTERS_10_18_port, ZN => n11730);
   U1614 : NAND4_X1 port map( A1 => n11733, A2 => n11732, A3 => n11731, A4 => 
                           n11730, ZN => n11734);
   U1615 : AOI22_X1 port map( A1 => n12036, A2 => n11735, B1 => n12034, B2 => 
                           n11734, ZN => n11736);
   U1616 : OAI21_X1 port map( B1 => n12196, B2 => n11737, A => n11736, ZN => 
                           N435);
   U1617 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_17_port, B1 => 
                           n12161, B2 => REGISTERS_18_17_port, ZN => n11741);
   U1618 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_17_port, B1 => 
                           n12157, B2 => REGISTERS_24_17_port, ZN => n11740);
   U1619 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_17_port, B1 => 
                           n12147, B2 => REGISTERS_27_17_port, ZN => n11739);
   U1620 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_17_port, B1 => 
                           n12150, B2 => REGISTERS_31_17_port, ZN => n11738);
   U1621 : NAND4_X1 port map( A1 => n11741, A2 => n11740, A3 => n11739, A4 => 
                           n11738, ZN => n11747);
   U1622 : AOI22_X1 port map( A1 => n12112, A2 => REGISTERS_26_17_port, B1 => 
                           n12119, B2 => REGISTERS_28_17_port, ZN => n11745);
   U1623 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_17_port, B1 => 
                           n11941, B2 => REGISTERS_19_17_port, ZN => n11744);
   U1624 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_17_port, B1 => 
                           n12159, B2 => REGISTERS_25_17_port, ZN => n11743);
   U1625 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_17_port, B1 => 
                           n12149, B2 => REGISTERS_23_17_port, ZN => n11742);
   U1626 : NAND4_X1 port map( A1 => n11745, A2 => n11744, A3 => n11743, A4 => 
                           n11742, ZN => n11746);
   U1627 : NOR2_X1 port map( A1 => n11747, A2 => n11746, ZN => n11759);
   U1628 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_17_port, B1 => 
                           n12180, B2 => REGISTERS_0_17_port, ZN => n11751);
   U1629 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_17_port, B1 => 
                           n12173, B2 => REGISTERS_2_17_port, ZN => n11750);
   U1630 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_17_port, B1 => 
                           n11887, B2 => REGISTERS_3_17_port, ZN => n11749);
   U1631 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_17_port, B1 => 
                           n12172, B2 => REGISTERS_7_17_port, ZN => n11748);
   U1632 : NAND4_X1 port map( A1 => n11751, A2 => n11750, A3 => n11749, A4 => 
                           n11748, ZN => n11757);
   U1633 : AOI22_X1 port map( A1 => n12173, A2 => REGISTERS_10_17_port, B1 => 
                           n12127, B2 => REGISTERS_8_17_port, ZN => n11755);
   U1634 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_17_port, B1 => 
                           n12049, B2 => REGISTERS_15_17_port, ZN => n11754);
   U1635 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_17_port, B1 => 
                           n12184, B2 => REGISTERS_11_17_port, ZN => n11753);
   U1636 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_17_port, B1 => 
                           n12097, B2 => REGISTERS_12_17_port, ZN => n11752);
   U1637 : NAND4_X1 port map( A1 => n11755, A2 => n11754, A3 => n11753, A4 => 
                           n11752, ZN => n11756);
   U1638 : AOI22_X1 port map( A1 => n12036, A2 => n11757, B1 => n12034, B2 => 
                           n11756, ZN => n11758);
   U1639 : OAI21_X1 port map( B1 => n12196, B2 => n11759, A => n11758, ZN => 
                           N434);
   U1640 : AOI22_X1 port map( A1 => n11853, A2 => REGISTERS_25_16_port, B1 => 
                           n12157, B2 => REGISTERS_24_16_port, ZN => n11763);
   U1641 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_16_port, B1 => 
                           n12146, B2 => REGISTERS_30_16_port, ZN => n11762);
   U1642 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_16_port, B1 => 
                           n11941, B2 => REGISTERS_19_16_port, ZN => n11761);
   U1643 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_16_port, B1 => 
                           n12150, B2 => REGISTERS_31_16_port, ZN => n11760);
   U1644 : NAND4_X1 port map( A1 => n11763, A2 => n11762, A3 => n11761, A4 => 
                           n11760, ZN => n11769);
   U1645 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_16_port, B1 => 
                           n12149, B2 => REGISTERS_23_16_port, ZN => n11767);
   U1646 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_16_port, B1 => 
                           n12147, B2 => REGISTERS_27_16_port, ZN => n11766);
   U1647 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_16_port, B1 => 
                           n12018, B2 => REGISTERS_17_16_port, ZN => n11765);
   U1648 : AOI22_X1 port map( A1 => n12112, A2 => REGISTERS_26_16_port, B1 => 
                           n12158, B2 => REGISTERS_16_16_port, ZN => n11764);
   U1649 : NAND4_X1 port map( A1 => n11767, A2 => n11766, A3 => n11765, A4 => 
                           n11764, ZN => n11768);
   U1650 : NOR2_X1 port map( A1 => n11769, A2 => n11768, ZN => n11781);
   U1651 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_16_port, B1 => 
                           n12077, B2 => REGISTERS_4_16_port, ZN => n11773);
   U1652 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_16_port, B1 => 
                           n12178, B2 => REGISTERS_7_16_port, ZN => n11772);
   U1653 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_16_port, B1 => 
                           n12180, B2 => REGISTERS_0_16_port, ZN => n11771);
   U1654 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_16_port, B1 => 
                           n12099, B2 => REGISTERS_3_16_port, ZN => n11770);
   U1655 : NAND4_X1 port map( A1 => n11773, A2 => n11772, A3 => n11771, A4 => 
                           n11770, ZN => n11779);
   U1656 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_14_16_port, B1 => 
                           n12097, B2 => REGISTERS_12_16_port, ZN => n11777);
   U1657 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_16_port, B1 => 
                           n12172, B2 => REGISTERS_15_16_port, ZN => n11776);
   U1658 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_16_port, B1 => 
                           n12135, B2 => REGISTERS_9_16_port, ZN => n11775);
   U1659 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_16_port, B1 => 
                           n12184, B2 => REGISTERS_11_16_port, ZN => n11774);
   U1660 : NAND4_X1 port map( A1 => n11777, A2 => n11776, A3 => n11775, A4 => 
                           n11774, ZN => n11778);
   U1661 : AOI22_X1 port map( A1 => n12036, A2 => n11779, B1 => n12034, B2 => 
                           n11778, ZN => n11780);
   U1662 : OAI21_X1 port map( B1 => n12196, B2 => n11781, A => n11780, ZN => 
                           N433);
   U1663 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_15_port, B1 => 
                           n12149, B2 => REGISTERS_23_15_port, ZN => n11785);
   U1664 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_15_port, B1 => 
                           n11941, B2 => REGISTERS_19_15_port, ZN => n11784);
   U1665 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_15_port, B1 => 
                           n12159, B2 => REGISTERS_25_15_port, ZN => n11783);
   U1666 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_15_port, B1 => 
                           n12119, B2 => REGISTERS_28_15_port, ZN => n11782);
   U1667 : NAND4_X1 port map( A1 => n11785, A2 => n11784, A3 => n11783, A4 => 
                           n11782, ZN => n11791);
   U1668 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_15_port, B1 => 
                           n12157, B2 => REGISTERS_24_15_port, ZN => n11789);
   U1669 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_15_port, B1 => 
                           n12114, B2 => REGISTERS_31_15_port, ZN => n11788);
   U1670 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_15_port, B1 => 
                           n11970, B2 => REGISTERS_22_15_port, ZN => n11787);
   U1671 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_15_port, B1 => 
                           n12147, B2 => REGISTERS_27_15_port, ZN => n11786);
   U1672 : NAND4_X1 port map( A1 => n11789, A2 => n11788, A3 => n11787, A4 => 
                           n11786, ZN => n11790);
   U1673 : NOR2_X1 port map( A1 => n11791, A2 => n11790, ZN => n11803);
   U1674 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_15_port, B1 => 
                           n12077, B2 => REGISTERS_4_15_port, ZN => n11795);
   U1675 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_15_port, B1 => 
                           n12127, B2 => REGISTERS_0_15_port, ZN => n11794);
   U1676 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_15_port, B1 => 
                           n12049, B2 => REGISTERS_7_15_port, ZN => n11793);
   U1677 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_15_port, B1 => 
                           n11887, B2 => REGISTERS_3_15_port, ZN => n11792);
   U1678 : NAND4_X1 port map( A1 => n11795, A2 => n11794, A3 => n11793, A4 => 
                           n11792, ZN => n11801);
   U1679 : AOI22_X1 port map( A1 => n12182, A2 => REGISTERS_10_15_port, B1 => 
                           n12172, B2 => REGISTERS_15_15_port, ZN => n11799);
   U1680 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_15_port, B1 => 
                           n12184, B2 => REGISTERS_11_15_port, ZN => n11798);
   U1681 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_15_port, B1 => 
                           n12054, B2 => REGISTERS_9_15_port, ZN => n11797);
   U1682 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_15_port, B1 => 
                           n12127, B2 => REGISTERS_8_15_port, ZN => n11796);
   U1683 : NAND4_X1 port map( A1 => n11799, A2 => n11798, A3 => n11797, A4 => 
                           n11796, ZN => n11800);
   U1684 : AOI22_X1 port map( A1 => n12036, A2 => n11801, B1 => n12034, B2 => 
                           n11800, ZN => n11802);
   U1685 : OAI21_X1 port map( B1 => n12144, B2 => n11803, A => n11802, ZN => 
                           N432);
   U1686 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_14_port, B1 => 
                           n12119, B2 => REGISTERS_28_14_port, ZN => n11807);
   U1687 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_14_port, B1 => 
                           n12146, B2 => REGISTERS_30_14_port, ZN => n11806);
   U1688 : AOI22_X1 port map( A1 => n12147, A2 => REGISTERS_27_14_port, B1 => 
                           n11941, B2 => REGISTERS_19_14_port, ZN => n11805);
   U1689 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_14_port, B1 => 
                           n12018, B2 => REGISTERS_17_14_port, ZN => n11804);
   U1690 : NAND4_X1 port map( A1 => n11807, A2 => n11806, A3 => n11805, A4 => 
                           n11804, ZN => n11813);
   U1691 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_14_port, B1 => 
                           n12114, B2 => REGISTERS_31_14_port, ZN => n11811);
   U1692 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_14_port, B1 => 
                           n12157, B2 => REGISTERS_24_14_port, ZN => n11810);
   U1693 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_14_port, B1 => 
                           n12159, B2 => REGISTERS_25_14_port, ZN => n11809);
   U1694 : AOI22_X1 port map( A1 => n11826, A2 => REGISTERS_18_14_port, B1 => 
                           n12149, B2 => REGISTERS_23_14_port, ZN => n11808);
   U1695 : NAND4_X1 port map( A1 => n11811, A2 => n11810, A3 => n11809, A4 => 
                           n11808, ZN => n11812);
   U1696 : NOR2_X1 port map( A1 => n11813, A2 => n11812, ZN => n11825);
   U1697 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_14_port, B1 => 
                           n12134, B2 => REGISTERS_0_14_port, ZN => n11817);
   U1698 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_4_14_port, B1 => 
                           n12099, B2 => REGISTERS_3_14_port, ZN => n11816);
   U1699 : AOI22_X1 port map( A1 => n12182, A2 => REGISTERS_2_14_port, B1 => 
                           n12049, B2 => REGISTERS_7_14_port, ZN => n11815);
   U1700 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_6_14_port, B1 => 
                           n12054, B2 => REGISTERS_1_14_port, ZN => n11814);
   U1701 : NAND4_X1 port map( A1 => n11817, A2 => n11816, A3 => n11815, A4 => 
                           n11814, ZN => n11823);
   U1702 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_14_14_port, B1 => 
                           n12097, B2 => REGISTERS_12_14_port, ZN => n11821);
   U1703 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_14_port, B1 => 
                           n12127, B2 => REGISTERS_8_14_port, ZN => n11820);
   U1704 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_14_port, B1 => 
                           n12181, B2 => REGISTERS_9_14_port, ZN => n11819);
   U1705 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_15_14_port, B1 => 
                           n12099, B2 => REGISTERS_11_14_port, ZN => n11818);
   U1706 : NAND4_X1 port map( A1 => n11821, A2 => n11820, A3 => n11819, A4 => 
                           n11818, ZN => n11822);
   U1707 : AOI22_X1 port map( A1 => n12036, A2 => n11823, B1 => n12034, B2 => 
                           n11822, ZN => n11824);
   U1708 : OAI21_X1 port map( B1 => n12196, B2 => n11825, A => n11824, ZN => 
                           N431);
   U1709 : AOI22_X1 port map( A1 => n11826, A2 => REGISTERS_18_13_port, B1 => 
                           n12147, B2 => REGISTERS_27_13_port, ZN => n11830);
   U1710 : AOI22_X1 port map( A1 => n11970, A2 => REGISTERS_22_13_port, B1 => 
                           n12018, B2 => REGISTERS_17_13_port, ZN => n11829);
   U1711 : AOI22_X1 port map( A1 => n12159, A2 => REGISTERS_25_13_port, B1 => 
                           n12157, B2 => REGISTERS_24_13_port, ZN => n11828);
   U1712 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_13_port, B1 => 
                           n12149, B2 => REGISTERS_23_13_port, ZN => n11827);
   U1713 : NAND4_X1 port map( A1 => n11830, A2 => n11829, A3 => n11828, A4 => 
                           n11827, ZN => n11836);
   U1714 : AOI22_X1 port map( A1 => n11900, A2 => REGISTERS_20_13_port, B1 => 
                           n12158, B2 => REGISTERS_16_13_port, ZN => n11834);
   U1715 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_13_port, B1 => 
                           n12119, B2 => REGISTERS_28_13_port, ZN => n11833);
   U1716 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_13_port, B1 => 
                           n12146, B2 => REGISTERS_30_13_port, ZN => n11832);
   U1717 : AOI22_X1 port map( A1 => n12150, A2 => REGISTERS_31_13_port, B1 => 
                           n11941, B2 => REGISTERS_19_13_port, ZN => n11831);
   U1718 : NAND4_X1 port map( A1 => n11834, A2 => n11833, A3 => n11832, A4 => 
                           n11831, ZN => n11835);
   U1719 : NOR2_X1 port map( A1 => n11836, A2 => n11835, ZN => n11848);
   U1720 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_13_port, B1 => 
                           n12049, B2 => REGISTERS_7_13_port, ZN => n11840);
   U1721 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_5_13_port, B1 => 
                           n12182, B2 => REGISTERS_2_13_port, ZN => n11839);
   U1722 : AOI22_X1 port map( A1 => n12180, A2 => REGISTERS_0_13_port, B1 => 
                           n11887, B2 => REGISTERS_3_13_port, ZN => n11838);
   U1723 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_13_port, B1 => 
                           n12054, B2 => REGISTERS_1_13_port, ZN => n11837);
   U1724 : NAND4_X1 port map( A1 => n11840, A2 => n11839, A3 => n11838, A4 => 
                           n11837, ZN => n11846);
   U1725 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_13_port, B1 => 
                           n12172, B2 => REGISTERS_15_13_port, ZN => n11844);
   U1726 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_13_port, B1 => 
                           n12077, B2 => REGISTERS_12_13_port, ZN => n11843);
   U1727 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_13_port, B1 => 
                           n12184, B2 => REGISTERS_11_13_port, ZN => n11842);
   U1728 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_13_port, B1 => 
                           n12134, B2 => REGISTERS_8_13_port, ZN => n11841);
   U1729 : NAND4_X1 port map( A1 => n11844, A2 => n11843, A3 => n11842, A4 => 
                           n11841, ZN => n11845);
   U1730 : AOI22_X1 port map( A1 => n12036, A2 => n11846, B1 => n12034, B2 => 
                           n11845, ZN => n11847);
   U1731 : OAI21_X1 port map( B1 => n12144, B2 => n11848, A => n11847, ZN => 
                           N430);
   U1732 : AOI22_X1 port map( A1 => n11970, A2 => REGISTERS_22_12_port, B1 => 
                           n12147, B2 => REGISTERS_27_12_port, ZN => n11852);
   U1733 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_12_port, B1 => 
                           n12157, B2 => REGISTERS_24_12_port, ZN => n11851);
   U1734 : AOI22_X1 port map( A1 => n12018, A2 => REGISTERS_17_12_port, B1 => 
                           n12114, B2 => REGISTERS_31_12_port, ZN => n11850);
   U1735 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_12_port, B1 => 
                           n12119, B2 => REGISTERS_28_12_port, ZN => n11849);
   U1736 : NAND4_X1 port map( A1 => n11852, A2 => n11851, A3 => n11850, A4 => 
                           n11849, ZN => n11859);
   U1737 : AOI22_X1 port map( A1 => n11900, A2 => REGISTERS_20_12_port, B1 => 
                           n12161, B2 => REGISTERS_18_12_port, ZN => n11857);
   U1738 : AOI22_X1 port map( A1 => n12086, A2 => REGISTERS_16_12_port, B1 => 
                           n12149, B2 => REGISTERS_23_12_port, ZN => n11856);
   U1739 : AOI22_X1 port map( A1 => n11853, A2 => REGISTERS_25_12_port, B1 => 
                           n11941, B2 => REGISTERS_19_12_port, ZN => n11855);
   U1740 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_12_port, B1 => 
                           n12146, B2 => REGISTERS_30_12_port, ZN => n11854);
   U1741 : NAND4_X1 port map( A1 => n11857, A2 => n11856, A3 => n11855, A4 => 
                           n11854, ZN => n11858);
   U1742 : NOR2_X1 port map( A1 => n11859, A2 => n11858, ZN => n11871);
   U1743 : AOI22_X1 port map( A1 => n12054, A2 => REGISTERS_1_12_port, B1 => 
                           n12178, B2 => REGISTERS_7_12_port, ZN => n11863);
   U1744 : AOI22_X1 port map( A1 => n12182, A2 => REGISTERS_2_12_port, B1 => 
                           n12134, B2 => REGISTERS_0_12_port, ZN => n11862);
   U1745 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_12_port, B1 => 
                           n12097, B2 => REGISTERS_4_12_port, ZN => n11861);
   U1746 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_12_port, B1 => 
                           n12099, B2 => REGISTERS_3_12_port, ZN => n11860);
   U1747 : NAND4_X1 port map( A1 => n11863, A2 => n11862, A3 => n11861, A4 => 
                           n11860, ZN => n11869);
   U1748 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_12_port, B1 => 
                           n12178, B2 => REGISTERS_15_12_port, ZN => n11867);
   U1749 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_12_port, B1 => 
                           n12135, B2 => REGISTERS_9_12_port, ZN => n11866);
   U1750 : AOI22_X1 port map( A1 => n12182, A2 => REGISTERS_10_12_port, B1 => 
                           n12180, B2 => REGISTERS_8_12_port, ZN => n11865);
   U1751 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_12_port, B1 => 
                           n12099, B2 => REGISTERS_11_12_port, ZN => n11864);
   U1752 : NAND4_X1 port map( A1 => n11867, A2 => n11866, A3 => n11865, A4 => 
                           n11864, ZN => n11868);
   U1753 : AOI22_X1 port map( A1 => n12036, A2 => n11869, B1 => n12034, B2 => 
                           n11868, ZN => n11870);
   U1754 : OAI21_X1 port map( B1 => n12196, B2 => n11871, A => n11870, ZN => 
                           N429);
   U1755 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_11_port, B1 => 
                           n12114, B2 => REGISTERS_31_11_port, ZN => n11875);
   U1756 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_11_port, B1 => 
                           n11941, B2 => REGISTERS_19_11_port, ZN => n11874);
   U1757 : AOI22_X1 port map( A1 => n12120, A2 => REGISTERS_21_11_port, B1 => 
                           n11970, B2 => REGISTERS_22_11_port, ZN => n11873);
   U1758 : AOI22_X1 port map( A1 => n11989, A2 => REGISTERS_24_11_port, B1 => 
                           n12147, B2 => REGISTERS_27_11_port, ZN => n11872);
   U1759 : NAND4_X1 port map( A1 => n11875, A2 => n11874, A3 => n11873, A4 => 
                           n11872, ZN => n11881);
   U1760 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_11_port, B1 => 
                           n12159, B2 => REGISTERS_25_11_port, ZN => n11879);
   U1761 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_11_port, B1 => 
                           n11900, B2 => REGISTERS_20_11_port, ZN => n11878);
   U1762 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_11_port, B1 => 
                           n12161, B2 => REGISTERS_18_11_port, ZN => n11877);
   U1763 : AOI22_X1 port map( A1 => n12018, A2 => REGISTERS_17_11_port, B1 => 
                           n12149, B2 => REGISTERS_23_11_port, ZN => n11876);
   U1764 : NAND4_X1 port map( A1 => n11879, A2 => n11878, A3 => n11877, A4 => 
                           n11876, ZN => n11880);
   U1765 : NOR2_X1 port map( A1 => n11881, A2 => n11880, ZN => n11895);
   U1766 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_11_port, B1 => 
                           n12173, B2 => REGISTERS_2_11_port, ZN => n11885);
   U1767 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_4_11_port, B1 => 
                           n12135, B2 => REGISTERS_1_11_port, ZN => n11884);
   U1768 : AOI22_X1 port map( A1 => n12127, A2 => REGISTERS_0_11_port, B1 => 
                           n12049, B2 => REGISTERS_7_11_port, ZN => n11883);
   U1769 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_6_11_port, B1 => 
                           n12099, B2 => REGISTERS_3_11_port, ZN => n11882);
   U1770 : NAND4_X1 port map( A1 => n11885, A2 => n11884, A3 => n11883, A4 => 
                           n11882, ZN => n11893);
   U1771 : AOI22_X1 port map( A1 => n11886, A2 => REGISTERS_13_11_port, B1 => 
                           n12132, B2 => REGISTERS_10_11_port, ZN => n11891);
   U1772 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_14_11_port, B1 => 
                           n12054, B2 => REGISTERS_9_11_port, ZN => n11890);
   U1773 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_11_port, B1 => 
                           n11887, B2 => REGISTERS_11_11_port, ZN => n11889);
   U1774 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_11_port, B1 => 
                           n12172, B2 => REGISTERS_15_11_port, ZN => n11888);
   U1775 : NAND4_X1 port map( A1 => n11891, A2 => n11890, A3 => n11889, A4 => 
                           n11888, ZN => n11892);
   U1776 : AOI22_X1 port map( A1 => n12036, A2 => n11893, B1 => n12034, B2 => 
                           n11892, ZN => n11894);
   U1777 : OAI21_X1 port map( B1 => n12196, B2 => n11895, A => n11894, ZN => 
                           N428);
   U1778 : AOI22_X1 port map( A1 => n12163, A2 => REGISTERS_28_10_port, B1 => 
                           n12159, B2 => REGISTERS_25_10_port, ZN => n11899);
   U1779 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_10_port, B1 => 
                           n12157, B2 => REGISTERS_24_10_port, ZN => n11898);
   U1780 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_10_port, B1 => 
                           n12149, B2 => REGISTERS_23_10_port, ZN => n11897);
   U1781 : AOI22_X1 port map( A1 => n12113, A2 => REGISTERS_30_10_port, B1 => 
                           n12151, B2 => REGISTERS_26_10_port, ZN => n11896);
   U1782 : NAND4_X1 port map( A1 => n11899, A2 => n11898, A3 => n11897, A4 => 
                           n11896, ZN => n11906);
   U1783 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_10_port, B1 => 
                           n12161, B2 => REGISTERS_18_10_port, ZN => n11904);
   U1784 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_10_port, B1 => 
                           n11941, B2 => REGISTERS_19_10_port, ZN => n11903);
   U1785 : AOI22_X1 port map( A1 => n11900, A2 => REGISTERS_20_10_port, B1 => 
                           n12147, B2 => REGISTERS_27_10_port, ZN => n11902);
   U1786 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_10_port, B1 => 
                           n12114, B2 => REGISTERS_31_10_port, ZN => n11901);
   U1787 : NAND4_X1 port map( A1 => n11904, A2 => n11903, A3 => n11902, A4 => 
                           n11901, ZN => n11905);
   U1788 : NOR2_X1 port map( A1 => n11906, A2 => n11905, ZN => n11918);
   U1789 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_10_port, B1 => 
                           n12182, B2 => REGISTERS_2_10_port, ZN => n11910);
   U1790 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_0_10_port, B1 => 
                           n12178, B2 => REGISTERS_7_10_port, ZN => n11909);
   U1791 : AOI22_X1 port map( A1 => n12135, A2 => REGISTERS_1_10_port, B1 => 
                           n12184, B2 => REGISTERS_3_10_port, ZN => n11908);
   U1792 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_10_port, B1 => 
                           n12077, B2 => REGISTERS_4_10_port, ZN => n11907);
   U1793 : NAND4_X1 port map( A1 => n11910, A2 => n11909, A3 => n11908, A4 => 
                           n11907, ZN => n11916);
   U1794 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_10_port, B1 => 
                           n12099, B2 => REGISTERS_11_10_port, ZN => n11914);
   U1795 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_12_10_port, B1 => 
                           n12134, B2 => REGISTERS_8_10_port, ZN => n11913);
   U1796 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_10_port, B1 => 
                           n12132, B2 => REGISTERS_10_10_port, ZN => n11912);
   U1797 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_10_port, B1 => 
                           n12172, B2 => REGISTERS_15_10_port, ZN => n11911);
   U1798 : NAND4_X1 port map( A1 => n11914, A2 => n11913, A3 => n11912, A4 => 
                           n11911, ZN => n11915);
   U1799 : AOI22_X1 port map( A1 => n12036, A2 => n11916, B1 => n12034, B2 => 
                           n11915, ZN => n11917);
   U1800 : OAI21_X1 port map( B1 => n12196, B2 => n11918, A => n11917, ZN => 
                           N427);
   U1801 : AOI22_X1 port map( A1 => n12163, A2 => REGISTERS_28_9_port, B1 => 
                           n12147, B2 => REGISTERS_27_9_port, ZN => n11922);
   U1802 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_9_port, B1 => 
                           n12086, B2 => REGISTERS_16_9_port, ZN => n11921);
   U1803 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_9_port, B1 => 
                           n11941, B2 => REGISTERS_19_9_port, ZN => n11920);
   U1804 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_9_port, B1 => 
                           n12112, B2 => REGISTERS_26_9_port, ZN => n11919);
   U1805 : NAND4_X1 port map( A1 => n11922, A2 => n11921, A3 => n11920, A4 => 
                           n11919, ZN => n11928);
   U1806 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_9_port, B1 => 
                           n12159, B2 => REGISTERS_25_9_port, ZN => n11926);
   U1807 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_9_port, B1 => 
                           n12149, B2 => REGISTERS_23_9_port, ZN => n11925);
   U1808 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_9_port, B1 => 
                           n12157, B2 => REGISTERS_24_9_port, ZN => n11924);
   U1809 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_9_port, B1 => 
                           n12114, B2 => REGISTERS_31_9_port, ZN => n11923);
   U1810 : NAND4_X1 port map( A1 => n11926, A2 => n11925, A3 => n11924, A4 => 
                           n11923, ZN => n11927);
   U1811 : NOR2_X1 port map( A1 => n11928, A2 => n11927, ZN => n11940);
   U1812 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_9_port, B1 => 
                           n12097, B2 => REGISTERS_4_9_port, ZN => n11932);
   U1813 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_9_port, B1 => 
                           n12132, B2 => REGISTERS_2_9_port, ZN => n11931);
   U1814 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_7_9_port, B1 => 
                           n12184, B2 => REGISTERS_3_9_port, ZN => n11930);
   U1815 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_9_port, B1 => 
                           n12127, B2 => REGISTERS_0_9_port, ZN => n11929);
   U1816 : NAND4_X1 port map( A1 => n11932, A2 => n11931, A3 => n11930, A4 => 
                           n11929, ZN => n11938);
   U1817 : AOI22_X1 port map( A1 => n12180, A2 => REGISTERS_8_9_port, B1 => 
                           n12049, B2 => REGISTERS_15_9_port, ZN => n11936);
   U1818 : AOI22_X1 port map( A1 => n12097, A2 => REGISTERS_12_9_port, B1 => 
                           n12135, B2 => REGISTERS_9_9_port, ZN => n11935);
   U1819 : AOI22_X1 port map( A1 => n12182, A2 => REGISTERS_10_9_port, B1 => 
                           n12099, B2 => REGISTERS_11_9_port, ZN => n11934);
   U1820 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_9_port, B1 => 
                           n12133, B2 => REGISTERS_14_9_port, ZN => n11933);
   U1821 : NAND4_X1 port map( A1 => n11936, A2 => n11935, A3 => n11934, A4 => 
                           n11933, ZN => n11937);
   U1822 : AOI22_X1 port map( A1 => n12036, A2 => n11938, B1 => n12034, B2 => 
                           n11937, ZN => n11939);
   U1823 : OAI21_X1 port map( B1 => n12144, B2 => n11940, A => n11939, ZN => 
                           N426);
   U1824 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_8_port, B1 => 
                           n11941, B2 => REGISTERS_19_8_port, ZN => n11945);
   U1825 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_8_port, B1 => 
                           n12147, B2 => REGISTERS_27_8_port, ZN => n11944);
   U1826 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_8_port, B1 => 
                           n11970, B2 => REGISTERS_22_8_port, ZN => n11943);
   U1827 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_8_port, B1 => 
                           n12159, B2 => REGISTERS_25_8_port, ZN => n11942);
   U1828 : NAND4_X1 port map( A1 => n11945, A2 => n11944, A3 => n11943, A4 => 
                           n11942, ZN => n11952);
   U1829 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_8_port, B1 => 
                           n12146, B2 => REGISTERS_30_8_port, ZN => n11950);
   U1830 : AOI22_X1 port map( A1 => n12013, A2 => REGISTERS_23_8_port, B1 => 
                           n12157, B2 => REGISTERS_24_8_port, ZN => n11949);
   U1831 : AOI22_X1 port map( A1 => n11946, A2 => REGISTERS_29_8_port, B1 => 
                           n12114, B2 => REGISTERS_31_8_port, ZN => n11948);
   U1832 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_8_port, B1 => 
                           n12161, B2 => REGISTERS_18_8_port, ZN => n11947);
   U1833 : NAND4_X1 port map( A1 => n11950, A2 => n11949, A3 => n11948, A4 => 
                           n11947, ZN => n11951);
   U1834 : NOR2_X1 port map( A1 => n11952, A2 => n11951, ZN => n11964);
   U1835 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_8_port, B1 => 
                           n12184, B2 => REGISTERS_3_8_port, ZN => n11956);
   U1836 : AOI22_X1 port map( A1 => n12127, A2 => REGISTERS_0_8_port, B1 => 
                           n12178, B2 => REGISTERS_7_8_port, ZN => n11955);
   U1837 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_8_port, B1 => 
                           n12054, B2 => REGISTERS_1_8_port, ZN => n11954);
   U1838 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_8_port, B1 => 
                           n12097, B2 => REGISTERS_4_8_port, ZN => n11953);
   U1839 : NAND4_X1 port map( A1 => n11956, A2 => n11955, A3 => n11954, A4 => 
                           n11953, ZN => n11962);
   U1840 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_8_port, B1 => 
                           n12182, B2 => REGISTERS_10_8_port, ZN => n11960);
   U1841 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_8_port, B1 => 
                           n12099, B2 => REGISTERS_11_8_port, ZN => n11959);
   U1842 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_13_8_port, B1 => 
                           n12180, B2 => REGISTERS_8_8_port, ZN => n11958);
   U1843 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_8_port, B1 => 
                           n12172, B2 => REGISTERS_15_8_port, ZN => n11957);
   U1844 : NAND4_X1 port map( A1 => n11960, A2 => n11959, A3 => n11958, A4 => 
                           n11957, ZN => n11961);
   U1845 : AOI22_X1 port map( A1 => n12036, A2 => n11962, B1 => n12034, B2 => 
                           n11961, ZN => n11963);
   U1846 : OAI21_X1 port map( B1 => n12196, B2 => n11964, A => n11963, ZN => 
                           N425);
   U1847 : AOI22_X1 port map( A1 => n12013, A2 => REGISTERS_23_7_port, B1 => 
                           n12159, B2 => REGISTERS_25_7_port, ZN => n11969);
   U1848 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_7_port, B1 => 
                           n12161, B2 => REGISTERS_18_7_port, ZN => n11968);
   U1849 : AOI22_X1 port map( A1 => n11965, A2 => REGISTERS_27_7_port, B1 => 
                           n12145, B2 => REGISTERS_19_7_port, ZN => n11967);
   U1850 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_7_port, B1 => 
                           n12157, B2 => REGISTERS_24_7_port, ZN => n11966);
   U1851 : NAND4_X1 port map( A1 => n11969, A2 => n11968, A3 => n11967, A4 => 
                           n11966, ZN => n11976);
   U1852 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_7_port, B1 => 
                           n12018, B2 => REGISTERS_17_7_port, ZN => n11974);
   U1853 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_7_port, B1 => 
                           n12086, B2 => REGISTERS_16_7_port, ZN => n11973);
   U1854 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_7_port, B1 => 
                           n11970, B2 => REGISTERS_22_7_port, ZN => n11972);
   U1855 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_7_port, B1 => 
                           n12113, B2 => REGISTERS_30_7_port, ZN => n11971);
   U1856 : NAND4_X1 port map( A1 => n11974, A2 => n11973, A3 => n11972, A4 => 
                           n11971, ZN => n11975);
   U1857 : NOR2_X1 port map( A1 => n11976, A2 => n11975, ZN => n11988);
   U1858 : AOI22_X1 port map( A1 => n12077, A2 => REGISTERS_4_7_port, B1 => 
                           n12173, B2 => REGISTERS_2_7_port, ZN => n11980);
   U1859 : AOI22_X1 port map( A1 => n12133, A2 => REGISTERS_6_7_port, B1 => 
                           n12049, B2 => REGISTERS_7_7_port, ZN => n11979);
   U1860 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_7_port, B1 => 
                           n12135, B2 => REGISTERS_1_7_port, ZN => n11978);
   U1861 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_0_7_port, B1 => 
                           n12099, B2 => REGISTERS_3_7_port, ZN => n11977);
   U1862 : NAND4_X1 port map( A1 => n11980, A2 => n11979, A3 => n11978, A4 => 
                           n11977, ZN => n11986);
   U1863 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_7_port, B1 => 
                           n12180, B2 => REGISTERS_8_7_port, ZN => n11984);
   U1864 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_7_port, B1 => 
                           n12135, B2 => REGISTERS_9_7_port, ZN => n11983);
   U1865 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_7_port, B1 => 
                           n12132, B2 => REGISTERS_10_7_port, ZN => n11982);
   U1866 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_15_7_port, B1 => 
                           n12184, B2 => REGISTERS_11_7_port, ZN => n11981);
   U1867 : NAND4_X1 port map( A1 => n11984, A2 => n11983, A3 => n11982, A4 => 
                           n11981, ZN => n11985);
   U1868 : AOI22_X1 port map( A1 => n12036, A2 => n11986, B1 => n12034, B2 => 
                           n11985, ZN => n11987);
   U1869 : OAI21_X1 port map( B1 => n12144, B2 => n11988, A => n11987, ZN => 
                           N424);
   U1870 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_6_port, B1 => 
                           n12149, B2 => REGISTERS_23_6_port, ZN => n11993);
   U1871 : AOI22_X1 port map( A1 => n11989, A2 => REGISTERS_24_6_port, B1 => 
                           n12145, B2 => REGISTERS_19_6_port, ZN => n11992);
   U1872 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_6_port, B1 => 
                           n12147, B2 => REGISTERS_27_6_port, ZN => n11991);
   U1873 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_6_port, B1 => 
                           n12113, B2 => REGISTERS_30_6_port, ZN => n11990);
   U1874 : NAND4_X1 port map( A1 => n11993, A2 => n11992, A3 => n11991, A4 => 
                           n11990, ZN => n11999);
   U1875 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_6_port, B1 => 
                           n12086, B2 => REGISTERS_16_6_port, ZN => n11997);
   U1876 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_6_port, B1 => 
                           n12112, B2 => REGISTERS_26_6_port, ZN => n11996);
   U1877 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_6_port, B1 => 
                           n12161, B2 => REGISTERS_18_6_port, ZN => n11995);
   U1878 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_6_port, B1 => 
                           n12159, B2 => REGISTERS_25_6_port, ZN => n11994);
   U1879 : NAND4_X1 port map( A1 => n11997, A2 => n11996, A3 => n11995, A4 => 
                           n11994, ZN => n11998);
   U1880 : NOR2_X1 port map( A1 => n11999, A2 => n11998, ZN => n12012);
   U1881 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_6_port, B1 => 
                           n12185, B2 => REGISTERS_6_6_port, ZN => n12003);
   U1882 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_6_port, B1 => 
                           n12127, B2 => REGISTERS_0_6_port, ZN => n12002);
   U1883 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_6_port, B1 => 
                           n12172, B2 => REGISTERS_7_6_port, ZN => n12001);
   U1884 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_6_port, B1 => 
                           n12099, B2 => REGISTERS_3_6_port, ZN => n12000);
   U1885 : NAND4_X1 port map( A1 => n12003, A2 => n12002, A3 => n12001, A4 => 
                           n12000, ZN => n12009);
   U1886 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_6_port, B1 => 
                           n12049, B2 => REGISTERS_15_6_port, ZN => n12007);
   U1887 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_6_port, B1 => 
                           n12184, B2 => REGISTERS_11_6_port, ZN => n12006);
   U1888 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_6_port, B1 => 
                           n12173, B2 => REGISTERS_10_6_port, ZN => n12005);
   U1889 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_6_port, B1 => 
                           n12127, B2 => REGISTERS_8_6_port, ZN => n12004);
   U1890 : NAND4_X1 port map( A1 => n12007, A2 => n12006, A3 => n12005, A4 => 
                           n12004, ZN => n12008);
   U1891 : AOI22_X1 port map( A1 => n12010, A2 => n12009, B1 => n12034, B2 => 
                           n12008, ZN => n12011);
   U1892 : OAI21_X1 port map( B1 => n12196, B2 => n12012, A => n12011, ZN => 
                           N423);
   U1893 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_5_port, B1 => 
                           n12112, B2 => REGISTERS_26_5_port, ZN => n12017);
   U1894 : AOI22_X1 port map( A1 => n12013, A2 => REGISTERS_23_5_port, B1 => 
                           n12145, B2 => REGISTERS_19_5_port, ZN => n12016);
   U1895 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_5_port, B1 => 
                           n12114, B2 => REGISTERS_31_5_port, ZN => n12015);
   U1896 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_5_port, B1 => 
                           n12157, B2 => REGISTERS_24_5_port, ZN => n12014);
   U1897 : NAND4_X1 port map( A1 => n12017, A2 => n12016, A3 => n12015, A4 => 
                           n12014, ZN => n12024);
   U1898 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_5_port, B1 => 
                           n12161, B2 => REGISTERS_18_5_port, ZN => n12022);
   U1899 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_5_port, B1 => 
                           n12159, B2 => REGISTERS_25_5_port, ZN => n12021);
   U1900 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_5_port, B1 => 
                           n12018, B2 => REGISTERS_17_5_port, ZN => n12020);
   U1901 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_5_port, B1 => 
                           n12147, B2 => REGISTERS_27_5_port, ZN => n12019);
   U1902 : NAND4_X1 port map( A1 => n12022, A2 => n12021, A3 => n12020, A4 => 
                           n12019, ZN => n12023);
   U1903 : NOR2_X1 port map( A1 => n12024, A2 => n12023, ZN => n12038);
   U1904 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_5_port, B1 => 
                           n12182, B2 => REGISTERS_2_5_port, ZN => n12028);
   U1905 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_5_port, B1 => 
                           n12178, B2 => REGISTERS_7_5_port, ZN => n12027);
   U1906 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_5_port, B1 => 
                           n12134, B2 => REGISTERS_0_5_port, ZN => n12026);
   U1907 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_5_port, B1 => 
                           n12099, B2 => REGISTERS_3_5_port, ZN => n12025);
   U1908 : NAND4_X1 port map( A1 => n12028, A2 => n12027, A3 => n12026, A4 => 
                           n12025, ZN => n12035);
   U1909 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_5_port, B1 => 
                           n12127, B2 => REGISTERS_8_5_port, ZN => n12032);
   U1910 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_5_port, B1 => 
                           n12172, B2 => REGISTERS_15_5_port, ZN => n12031);
   U1911 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_5_port, B1 => 
                           n12054, B2 => REGISTERS_9_5_port, ZN => n12030);
   U1912 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_5_port, B1 => 
                           n12184, B2 => REGISTERS_11_5_port, ZN => n12029);
   U1913 : NAND4_X1 port map( A1 => n12032, A2 => n12031, A3 => n12030, A4 => 
                           n12029, ZN => n12033);
   U1914 : AOI22_X1 port map( A1 => n12036, A2 => n12035, B1 => n12034, B2 => 
                           n12033, ZN => n12037);
   U1915 : OAI21_X1 port map( B1 => n12144, B2 => n12038, A => n12037, ZN => 
                           N422);
   U1916 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_4_port, B1 => 
                           n12149, B2 => REGISTERS_23_4_port, ZN => n12042);
   U1917 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_4_port, B1 => 
                           n12112, B2 => REGISTERS_26_4_port, ZN => n12041);
   U1918 : AOI22_X1 port map( A1 => n12159, A2 => REGISTERS_25_4_port, B1 => 
                           n12157, B2 => REGISTERS_24_4_port, ZN => n12040);
   U1919 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_4_port, B1 => 
                           n12145, B2 => REGISTERS_19_4_port, ZN => n12039);
   U1920 : NAND4_X1 port map( A1 => n12042, A2 => n12041, A3 => n12040, A4 => 
                           n12039, ZN => n12048);
   U1921 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_4_port, B1 => 
                           n12147, B2 => REGISTERS_27_4_port, ZN => n12046);
   U1922 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_4_port, B1 => 
                           n12114, B2 => REGISTERS_31_4_port, ZN => n12045);
   U1923 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_4_port, B1 => 
                           n12086, B2 => REGISTERS_16_4_port, ZN => n12044);
   U1924 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_4_port, B1 => 
                           n12161, B2 => REGISTERS_18_4_port, ZN => n12043);
   U1925 : NAND4_X1 port map( A1 => n12046, A2 => n12045, A3 => n12044, A4 => 
                           n12043, ZN => n12047);
   U1926 : NOR2_X1 port map( A1 => n12048, A2 => n12047, ZN => n12062);
   U1927 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_4_port, B1 => 
                           n12099, B2 => REGISTERS_3_4_port, ZN => n12053);
   U1928 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_4_port, B1 => 
                           n12182, B2 => REGISTERS_2_4_port, ZN => n12052);
   U1929 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_4_port, B1 => 
                           n12049, B2 => REGISTERS_7_4_port, ZN => n12051);
   U1930 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_4_port, B1 => 
                           n12134, B2 => REGISTERS_0_4_port, ZN => n12050);
   U1931 : NAND4_X1 port map( A1 => n12053, A2 => n12052, A3 => n12051, A4 => 
                           n12050, ZN => n12060);
   U1932 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_4_port, B1 => 
                           n12054, B2 => REGISTERS_9_4_port, ZN => n12058);
   U1933 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_4_port, B1 => 
                           n12184, B2 => REGISTERS_11_4_port, ZN => n12057);
   U1934 : AOI22_X1 port map( A1 => n12173, A2 => REGISTERS_10_4_port, B1 => 
                           n12178, B2 => REGISTERS_15_4_port, ZN => n12056);
   U1935 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_4_port, B1 => 
                           n12127, B2 => REGISTERS_8_4_port, ZN => n12055);
   U1936 : NAND4_X1 port map( A1 => n12058, A2 => n12057, A3 => n12056, A4 => 
                           n12055, ZN => n12059);
   U1937 : AOI22_X1 port map( A1 => n12193, A2 => n12060, B1 => n12191, B2 => 
                           n12059, ZN => n12061);
   U1938 : OAI21_X1 port map( B1 => n12196, B2 => n12062, A => n12061, ZN => 
                           N421);
   U1939 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_3_port, B1 => 
                           n12147, B2 => REGISTERS_27_3_port, ZN => n12066);
   U1940 : AOI22_X1 port map( A1 => n12149, A2 => REGISTERS_23_3_port, B1 => 
                           n12145, B2 => REGISTERS_19_3_port, ZN => n12065);
   U1941 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_3_port, B1 => 
                           n12157, B2 => REGISTERS_24_3_port, ZN => n12064);
   U1942 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_3_port, B1 => 
                           n12086, B2 => REGISTERS_16_3_port, ZN => n12063);
   U1943 : NAND4_X1 port map( A1 => n12066, A2 => n12065, A3 => n12064, A4 => 
                           n12063, ZN => n12072);
   U1944 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_3_port, B1 => 
                           n12113, B2 => REGISTERS_30_3_port, ZN => n12070);
   U1945 : AOI22_X1 port map( A1 => n12114, A2 => REGISTERS_31_3_port, B1 => 
                           n12161, B2 => REGISTERS_18_3_port, ZN => n12069);
   U1946 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_3_port, B1 => 
                           n12119, B2 => REGISTERS_28_3_port, ZN => n12068);
   U1947 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_3_port, B1 => 
                           n12159, B2 => REGISTERS_25_3_port, ZN => n12067);
   U1948 : NAND4_X1 port map( A1 => n12070, A2 => n12069, A3 => n12068, A4 => 
                           n12067, ZN => n12071);
   U1949 : NOR2_X1 port map( A1 => n12072, A2 => n12071, ZN => n12085);
   U1950 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_3_port, B1 => 
                           n12172, B2 => REGISTERS_7_3_port, ZN => n12076);
   U1951 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_3_port, B1 => 
                           n12097, B2 => REGISTERS_4_3_port, ZN => n12075);
   U1952 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_3_port, B1 => 
                           n12099, B2 => REGISTERS_3_3_port, ZN => n12074);
   U1953 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_3_port, B1 => 
                           n12127, B2 => REGISTERS_0_3_port, ZN => n12073);
   U1954 : NAND4_X1 port map( A1 => n12076, A2 => n12075, A3 => n12074, A4 => 
                           n12073, ZN => n12083);
   U1955 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_3_port, B1 => 
                           n12077, B2 => REGISTERS_12_3_port, ZN => n12081);
   U1956 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_3_port, B1 => 
                           n12172, B2 => REGISTERS_15_3_port, ZN => n12080);
   U1957 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_3_port, B1 => 
                           n12135, B2 => REGISTERS_9_3_port, ZN => n12079);
   U1958 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_3_port, B1 => 
                           n12184, B2 => REGISTERS_11_3_port, ZN => n12078);
   U1959 : NAND4_X1 port map( A1 => n12081, A2 => n12080, A3 => n12079, A4 => 
                           n12078, ZN => n12082);
   U1960 : AOI22_X1 port map( A1 => n12193, A2 => n12083, B1 => n12191, B2 => 
                           n12082, ZN => n12084);
   U1961 : OAI21_X1 port map( B1 => n12144, B2 => n12085, A => n12084, ZN => 
                           N420);
   U1962 : AOI22_X1 port map( A1 => n12151, A2 => REGISTERS_26_2_port, B1 => 
                           n12086, B2 => REGISTERS_16_2_port, ZN => n12090);
   U1963 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_2_port, B1 => 
                           n12113, B2 => REGISTERS_30_2_port, ZN => n12089);
   U1964 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_2_port, B1 => 
                           n12147, B2 => REGISTERS_27_2_port, ZN => n12088);
   U1965 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_2_port, B1 => 
                           n12157, B2 => REGISTERS_24_2_port, ZN => n12087);
   U1966 : NAND4_X1 port map( A1 => n12090, A2 => n12089, A3 => n12088, A4 => 
                           n12087, ZN => n12096);
   U1967 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_2_port, B1 => 
                           n12159, B2 => REGISTERS_25_2_port, ZN => n12094);
   U1968 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_2_port, B1 => 
                           n12149, B2 => REGISTERS_23_2_port, ZN => n12093);
   U1969 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_2_port, B1 => 
                           n12145, B2 => REGISTERS_19_2_port, ZN => n12092);
   U1970 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_2_port, B1 => 
                           n12114, B2 => REGISTERS_31_2_port, ZN => n12091);
   U1971 : NAND4_X1 port map( A1 => n12094, A2 => n12093, A3 => n12092, A4 => 
                           n12091, ZN => n12095);
   U1972 : NOR2_X1 port map( A1 => n12096, A2 => n12095, ZN => n12111);
   U1973 : AOI22_X1 port map( A1 => n12098, A2 => REGISTERS_5_2_port, B1 => 
                           n12097, B2 => REGISTERS_4_2_port, ZN => n12103);
   U1974 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_2_port, B1 => 
                           n12180, B2 => REGISTERS_0_2_port, ZN => n12102);
   U1975 : AOI22_X1 port map( A1 => n12172, A2 => REGISTERS_7_2_port, B1 => 
                           n12099, B2 => REGISTERS_3_2_port, ZN => n12101);
   U1976 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_2_port, B1 => 
                           n12173, B2 => REGISTERS_2_2_port, ZN => n12100);
   U1977 : NAND4_X1 port map( A1 => n12103, A2 => n12102, A3 => n12101, A4 => 
                           n12100, ZN => n12109);
   U1978 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_2_port, B1 => 
                           n12180, B2 => REGISTERS_8_2_port, ZN => n12107);
   U1979 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_2_port, B1 => 
                           n12173, B2 => REGISTERS_10_2_port, ZN => n12106);
   U1980 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_14_2_port, B1 => 
                           n12184, B2 => REGISTERS_11_2_port, ZN => n12105);
   U1981 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_2_port, B1 => 
                           n12172, B2 => REGISTERS_15_2_port, ZN => n12104);
   U1982 : NAND4_X1 port map( A1 => n12107, A2 => n12106, A3 => n12105, A4 => 
                           n12104, ZN => n12108);
   U1983 : AOI22_X1 port map( A1 => n12193, A2 => n12109, B1 => n12191, B2 => 
                           n12108, ZN => n12110);
   U1984 : OAI21_X1 port map( B1 => n12196, B2 => n12111, A => n12110, ZN => 
                           N419);
   U1985 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_1_port, B1 => 
                           n12112, B2 => REGISTERS_26_1_port, ZN => n12118);
   U1986 : AOI22_X1 port map( A1 => n12149, A2 => REGISTERS_23_1_port, B1 => 
                           n12145, B2 => REGISTERS_19_1_port, ZN => n12117);
   U1987 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_1_port, B1 => 
                           n12113, B2 => REGISTERS_30_1_port, ZN => n12116);
   U1988 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_1_port, B1 => 
                           n12114, B2 => REGISTERS_31_1_port, ZN => n12115);
   U1989 : NAND4_X1 port map( A1 => n12118, A2 => n12117, A3 => n12116, A4 => 
                           n12115, ZN => n12126);
   U1990 : AOI22_X1 port map( A1 => n12119, A2 => REGISTERS_28_1_port, B1 => 
                           n12147, B2 => REGISTERS_27_1_port, ZN => n12124);
   U1991 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_1_port, B1 => 
                           n12120, B2 => REGISTERS_21_1_port, ZN => n12123);
   U1992 : AOI22_X1 port map( A1 => n12161, A2 => REGISTERS_18_1_port, B1 => 
                           n12159, B2 => REGISTERS_25_1_port, ZN => n12122);
   U1993 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_1_port, B1 => 
                           n12157, B2 => REGISTERS_24_1_port, ZN => n12121);
   U1994 : NAND4_X1 port map( A1 => n12124, A2 => n12123, A3 => n12122, A4 => 
                           n12121, ZN => n12125);
   U1995 : NOR2_X1 port map( A1 => n12126, A2 => n12125, ZN => n12143);
   U1996 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_2_1_port, B1 => 
                           n12172, B2 => REGISTERS_7_1_port, ZN => n12131);
   U1997 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_1_port, B1 => 
                           n12184, B2 => REGISTERS_3_1_port, ZN => n12130);
   U1998 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_1_port, B1 => 
                           n12127, B2 => REGISTERS_0_1_port, ZN => n12129);
   U1999 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_1_port, B1 => 
                           n12135, B2 => REGISTERS_1_1_port, ZN => n12128);
   U2000 : NAND4_X1 port map( A1 => n12131, A2 => n12130, A3 => n12129, A4 => 
                           n12128, ZN => n12141);
   U2001 : AOI22_X1 port map( A1 => n12132, A2 => REGISTERS_10_1_port, B1 => 
                           n12178, B2 => REGISTERS_15_1_port, ZN => n12139);
   U2002 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_1_port, B1 => 
                           n12133, B2 => REGISTERS_14_1_port, ZN => n12138);
   U2003 : AOI22_X1 port map( A1 => n12134, A2 => REGISTERS_8_1_port, B1 => 
                           n12184, B2 => REGISTERS_11_1_port, ZN => n12137);
   U2004 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_1_port, B1 => 
                           n12135, B2 => REGISTERS_9_1_port, ZN => n12136);
   U2005 : NAND4_X1 port map( A1 => n12139, A2 => n12138, A3 => n12137, A4 => 
                           n12136, ZN => n12140);
   U2006 : AOI22_X1 port map( A1 => n12193, A2 => n12141, B1 => n12191, B2 => 
                           n12140, ZN => n12142);
   U2007 : OAI21_X1 port map( B1 => n12144, B2 => n12143, A => n12142, ZN => 
                           N418);
   U2008 : AOI22_X1 port map( A1 => n12146, A2 => REGISTERS_30_0_port, B1 => 
                           n12145, B2 => REGISTERS_19_0_port, ZN => n12156);
   U2009 : AOI22_X1 port map( A1 => n12148, A2 => REGISTERS_22_0_port, B1 => 
                           n12147, B2 => REGISTERS_27_0_port, ZN => n12155);
   U2010 : AOI22_X1 port map( A1 => n12150, A2 => REGISTERS_31_0_port, B1 => 
                           n12149, B2 => REGISTERS_23_0_port, ZN => n12154);
   U2011 : AOI22_X1 port map( A1 => n12152, A2 => REGISTERS_20_0_port, B1 => 
                           n12151, B2 => REGISTERS_26_0_port, ZN => n12153);
   U2012 : NAND4_X1 port map( A1 => n12156, A2 => n12155, A3 => n12154, A4 => 
                           n12153, ZN => n12170);
   U2013 : AOI22_X1 port map( A1 => n12158, A2 => REGISTERS_16_0_port, B1 => 
                           n12157, B2 => REGISTERS_24_0_port, ZN => n12168);
   U2014 : AOI22_X1 port map( A1 => n12160, A2 => REGISTERS_21_0_port, B1 => 
                           n12159, B2 => REGISTERS_25_0_port, ZN => n12167);
   U2015 : AOI22_X1 port map( A1 => n12162, A2 => REGISTERS_17_0_port, B1 => 
                           n12161, B2 => REGISTERS_18_0_port, ZN => n12166);
   U2016 : AOI22_X1 port map( A1 => n12164, A2 => REGISTERS_29_0_port, B1 => 
                           n12163, B2 => REGISTERS_28_0_port, ZN => n12165);
   U2017 : NAND4_X1 port map( A1 => n12168, A2 => n12167, A3 => n12166, A4 => 
                           n12165, ZN => n12169);
   U2018 : NOR2_X1 port map( A1 => n12170, A2 => n12169, ZN => n12195);
   U2019 : AOI22_X1 port map( A1 => n12171, A2 => REGISTERS_6_0_port, B1 => 
                           n12180, B2 => REGISTERS_0_0_port, ZN => n12177);
   U2020 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_4_0_port, B1 => 
                           n12172, B2 => REGISTERS_7_0_port, ZN => n12176);
   U2021 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_1_0_port, B1 => 
                           n12173, B2 => REGISTERS_2_0_port, ZN => n12175);
   U2022 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_5_0_port, B1 => 
                           n12184, B2 => REGISTERS_3_0_port, ZN => n12174);
   U2023 : NAND4_X1 port map( A1 => n12177, A2 => n12176, A3 => n12175, A4 => 
                           n12174, ZN => n12192);
   U2024 : AOI22_X1 port map( A1 => n12179, A2 => REGISTERS_13_0_port, B1 => 
                           n12178, B2 => REGISTERS_15_0_port, ZN => n12189);
   U2025 : AOI22_X1 port map( A1 => n12181, A2 => REGISTERS_9_0_port, B1 => 
                           n12180, B2 => REGISTERS_8_0_port, ZN => n12188);
   U2026 : AOI22_X1 port map( A1 => n12183, A2 => REGISTERS_12_0_port, B1 => 
                           n12182, B2 => REGISTERS_10_0_port, ZN => n12187);
   U2027 : AOI22_X1 port map( A1 => n12185, A2 => REGISTERS_14_0_port, B1 => 
                           n12184, B2 => REGISTERS_11_0_port, ZN => n12186);
   U2028 : NAND4_X1 port map( A1 => n12189, A2 => n12188, A3 => n12187, A4 => 
                           n12186, ZN => n12190);
   U2029 : AOI22_X1 port map( A1 => n12193, A2 => n12192, B1 => n12191, B2 => 
                           n12190, ZN => n12194);
   U2030 : OAI21_X1 port map( B1 => n12196, B2 => n12195, A => n12194, ZN => 
                           N417);
   U2031 : NAND3_X1 port map( A1 => n11229, A2 => ENABLE, A3 => RD1, ZN => 
                           n12978);
   U2032 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n12205)
                           ;
   U2033 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n12198);
   U2034 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => n12198, ZN => n12214);
   U2035 : NOR2_X1 port map( A1 => n12205, A2 => n12214, ZN => n12867);
   U2036 : CLKBUF_X1 port map( A => n12867, Z => n12926);
   U2037 : INV_X1 port map( A => ADD_RD1(2), ZN => n12204);
   U2038 : INV_X1 port map( A => ADD_RD1(0), ZN => n12203);
   U2039 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => n12204, A3 => n12203, ZN 
                           => n12220);
   U2040 : INV_X1 port map( A => ADD_RD1(3), ZN => n12225);
   U2041 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n12225, ZN => n12206);
   U2042 : NOR2_X1 port map( A1 => n12220, A2 => n12206, ZN => n12874);
   U2043 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n12926, B1 => 
                           REGISTERS_18_31_port, B2 => n12874, ZN => n12202);
   U2044 : INV_X1 port map( A => ADD_RD1(1), ZN => n12197);
   U2045 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => n12197,
                           ZN => n12215);
   U2046 : NOR2_X1 port map( A1 => n12205, A2 => n12215, ZN => n12843);
   U2047 : CLKBUF_X1 port map( A => n12843, Z => n12930);
   U2048 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n12204, A3 => n12197, ZN 
                           => n12219);
   U2049 : NOR2_X1 port map( A1 => n12206, A2 => n12219, ZN => n12939);
   U2050 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n12930, B1 => 
                           REGISTERS_17_31_port, B2 => n12939, ZN => n12201);
   U2051 : NOR2_X1 port map( A1 => n12206, A2 => n12215, ZN => n12940);
   U2052 : CLKBUF_X1 port map( A => n12940, Z => n12902);
   U2053 : NAND2_X1 port map( A1 => n12198, A2 => n12204, ZN => n12213);
   U2054 : NOR2_X1 port map( A1 => n12205, A2 => n12213, ZN => n12613);
   U2055 : CLKBUF_X1 port map( A => n12613, Z => n12942);
   U2056 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n12902, B1 => 
                           REGISTERS_24_31_port, B2 => n12942, ZN => n12200);
   U2057 : NOR2_X1 port map( A1 => n12206, A2 => n12214, ZN => n12771);
   U2058 : CLKBUF_X1 port map( A => n12771, Z => n12931);
   U2059 : NOR2_X1 port map( A1 => n12206, A2 => n12213, ZN => n12865);
   U2060 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n12931, B1 => 
                           REGISTERS_16_31_port, B2 => n12865, ZN => n12199);
   U2061 : NAND4_X1 port map( A1 => n12202, A2 => n12201, A3 => n12200, A4 => 
                           n12199, ZN => n12212);
   U2062 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n12203,
                           ZN => n12216);
   U2063 : NOR2_X1 port map( A1 => n12206, A2 => n12216, ZN => n12844);
   U2064 : CLKBUF_X1 port map( A => n12844, Z => n12944);
   U2065 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), A3 => 
                           ADD_RD1(0), ZN => n12218);
   U2066 : NOR2_X1 port map( A1 => n12206, A2 => n12218, ZN => n12658);
   U2067 : CLKBUF_X1 port map( A => n12658, Z => n12927);
   U2068 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n12944, B1 => 
                           REGISTERS_23_31_port, B2 => n12927, ZN => n12210);
   U2069 : NOR2_X1 port map( A1 => n12205, A2 => n12220, ZN => n12929);
   U2070 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => n12204,
                           ZN => n12217);
   U2071 : NOR2_X1 port map( A1 => n12205, A2 => n12217, ZN => n12872);
   U2072 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n12929, B1 => 
                           REGISTERS_27_31_port, B2 => n12872, ZN => n12209);
   U2073 : NOR2_X1 port map( A1 => n12205, A2 => n12216, ZN => n12678);
   U2074 : CLKBUF_X1 port map( A => n12678, Z => n12941);
   U2075 : NOR2_X1 port map( A1 => n12205, A2 => n12219, ZN => n12586);
   U2076 : CLKBUF_X1 port map( A => n12586, Z => n12938);
   U2077 : AOI22_X1 port map( A1 => REGISTERS_30_31_port, A2 => n12941, B1 => 
                           REGISTERS_25_31_port, B2 => n12938, ZN => n12208);
   U2078 : NOR2_X1 port map( A1 => n12205, A2 => n12218, ZN => n12838);
   U2079 : CLKBUF_X1 port map( A => n12838, Z => n12943);
   U2080 : NOR2_X1 port map( A1 => n12217, A2 => n12206, ZN => n12677);
   U2081 : CLKBUF_X1 port map( A => n12677, Z => n12925);
   U2082 : AOI22_X1 port map( A1 => REGISTERS_31_31_port, A2 => n12943, B1 => 
                           REGISTERS_19_31_port, B2 => n12925, ZN => n12207);
   U2083 : NAND4_X1 port map( A1 => n12210, A2 => n12209, A3 => n12208, A4 => 
                           n12207, ZN => n12211);
   U2084 : NOR2_X1 port map( A1 => n12212, A2 => n12211, ZN => n12233);
   U2085 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n12924, 
                           ZN => n12975);
   U2086 : CLKBUF_X1 port map( A => n12975, Z => n12788);
   U2087 : INV_X1 port map( A => n12213, ZN => n12915);
   U2088 : CLKBUF_X1 port map( A => n12915, Z => n12955);
   U2089 : INV_X1 port map( A => n12214, ZN => n12965);
   U2090 : CLKBUF_X1 port map( A => n12965, Z => n12913);
   U2091 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n12955, B1 => 
                           REGISTERS_4_31_port, B2 => n12913, ZN => n12224);
   U2092 : INV_X1 port map( A => n12215, ZN => n12805);
   U2093 : CLKBUF_X1 port map( A => n12805, Z => n12963);
   U2094 : INV_X1 port map( A => n12216, ZN => n12889);
   U2095 : CLKBUF_X1 port map( A => n12889, Z => n12883);
   U2096 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n12963, B1 => 
                           REGISTERS_6_31_port, B2 => n12883, ZN => n12223);
   U2097 : INV_X1 port map( A => n12217, ZN => n12852);
   U2098 : CLKBUF_X1 port map( A => n12852, Z => n12914);
   U2099 : INV_X1 port map( A => n12218, ZN => n12851);
   U2100 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n12914, B1 => 
                           REGISTERS_7_31_port, B2 => n12851, ZN => n12222);
   U2101 : INV_X1 port map( A => n12219, ZN => n12884);
   U2102 : CLKBUF_X1 port map( A => n12884, Z => n12967);
   U2103 : INV_X1 port map( A => n12220, ZN => n12966);
   U2104 : CLKBUF_X1 port map( A => n12966, Z => n12881);
   U2105 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n12967, B1 => 
                           REGISTERS_2_31_port, B2 => n12881, ZN => n12221);
   U2106 : NAND4_X1 port map( A1 => n12224, A2 => n12223, A3 => n12222, A4 => 
                           n12221, ZN => n12231);
   U2107 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n12225, A3 => n12924, ZN 
                           => n12973);
   U2108 : CLKBUF_X1 port map( A => n12973, Z => n12811);
   U2109 : CLKBUF_X1 port map( A => n12805, Z => n12951);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_10_31_port, A2 => n12966, B1 => 
                           REGISTERS_13_31_port, B2 => n12951, ZN => n12229);
   U2111 : CLKBUF_X1 port map( A => n12915, Z => n12962);
   U2112 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n12884, B1 => 
                           REGISTERS_8_31_port, B2 => n12962, ZN => n12228);
   U2113 : CLKBUF_X1 port map( A => n12889, Z => n12964);
   U2114 : CLKBUF_X1 port map( A => n12851, Z => n12961);
   U2115 : AOI22_X1 port map( A1 => REGISTERS_14_31_port, A2 => n12964, B1 => 
                           REGISTERS_15_31_port, B2 => n12961, ZN => n12227);
   U2116 : CLKBUF_X1 port map( A => n12965, Z => n12882);
   U2117 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n12882, B1 => 
                           REGISTERS_11_31_port, B2 => n12852, ZN => n12226);
   U2118 : NAND4_X1 port map( A1 => n12229, A2 => n12228, A3 => n12227, A4 => 
                           n12226, ZN => n12230);
   U2119 : AOI22_X1 port map( A1 => n12788, A2 => n12231, B1 => n12811, B2 => 
                           n12230, ZN => n12232);
   U2120 : OAI21_X1 port map( B1 => n12924, B2 => n12233, A => n12232, ZN => 
                           N416);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n12867, B1 => 
                           REGISTERS_25_30_port, B2 => n12586, ZN => n12237);
   U2122 : CLKBUF_X1 port map( A => n12872, Z => n12932);
   U2123 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n12932, B1 => 
                           REGISTERS_16_30_port, B2 => n12865, ZN => n12236);
   U2124 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n12942, B1 => 
                           REGISTERS_26_30_port, B2 => n12929, ZN => n12235);
   U2125 : CLKBUF_X1 port map( A => n12939, Z => n12873);
   U2126 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n12873, B1 => 
                           REGISTERS_29_30_port, B2 => n12843, ZN => n12234);
   U2127 : NAND4_X1 port map( A1 => n12237, A2 => n12236, A3 => n12235, A4 => 
                           n12234, ZN => n12243);
   U2128 : AOI22_X1 port map( A1 => REGISTERS_22_30_port, A2 => n12944, B1 => 
                           REGISTERS_23_30_port, B2 => n12658, ZN => n12241);
   U2129 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n12902, B1 => 
                           REGISTERS_31_30_port, B2 => n12943, ZN => n12240);
   U2130 : AOI22_X1 port map( A1 => REGISTERS_19_30_port, A2 => n12925, B1 => 
                           REGISTERS_18_30_port, B2 => n12874, ZN => n12239);
   U2131 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n12931, B1 => 
                           REGISTERS_30_30_port, B2 => n12941, ZN => n12238);
   U2132 : NAND4_X1 port map( A1 => n12241, A2 => n12240, A3 => n12239, A4 => 
                           n12238, ZN => n12242);
   U2133 : NOR2_X1 port map( A1 => n12243, A2 => n12242, ZN => n12255);
   U2134 : CLKBUF_X1 port map( A => n12884, Z => n12952);
   U2135 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n12805, B1 => 
                           REGISTERS_1_30_port, B2 => n12952, ZN => n12247);
   U2136 : CLKBUF_X1 port map( A => n12852, Z => n12960);
   U2137 : AOI22_X1 port map( A1 => REGISTERS_6_30_port, A2 => n12964, B1 => 
                           REGISTERS_3_30_port, B2 => n12960, ZN => n12246);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n12882, B1 => 
                           REGISTERS_0_30_port, B2 => n12962, ZN => n12245);
   U2139 : CLKBUF_X1 port map( A => n12851, Z => n12953);
   U2140 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n12953, B1 => 
                           REGISTERS_2_30_port, B2 => n12881, ZN => n12244);
   U2141 : NAND4_X1 port map( A1 => n12247, A2 => n12246, A3 => n12245, A4 => 
                           n12244, ZN => n12253);
   U2142 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n12955, B1 => 
                           REGISTERS_9_30_port, B2 => n12952, ZN => n12251);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_11_30_port, A2 => n12914, B1 => 
                           REGISTERS_10_30_port, B2 => n12881, ZN => n12250);
   U2144 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n12953, B1 => 
                           REGISTERS_13_30_port, B2 => n12951, ZN => n12249);
   U2145 : AOI22_X1 port map( A1 => REGISTERS_14_30_port, A2 => n12964, B1 => 
                           REGISTERS_12_30_port, B2 => n12913, ZN => n12248);
   U2146 : NAND4_X1 port map( A1 => n12251, A2 => n12250, A3 => n12249, A4 => 
                           n12248, ZN => n12252);
   U2147 : AOI22_X1 port map( A1 => n12788, A2 => n12253, B1 => n12811, B2 => 
                           n12252, ZN => n12254);
   U2148 : OAI21_X1 port map( B1 => n12924, B2 => n12255, A => n12254, ZN => 
                           N415);
   U2149 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n12931, B1 => 
                           REGISTERS_21_29_port, B2 => n12940, ZN => n12259);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_22_29_port, A2 => n12944, B1 => 
                           REGISTERS_24_29_port, B2 => n12942, ZN => n12258);
   U2151 : AOI22_X1 port map( A1 => REGISTERS_31_29_port, A2 => n12943, B1 => 
                           REGISTERS_17_29_port, B2 => n12939, ZN => n12257);
   U2152 : CLKBUF_X1 port map( A => n12929, Z => n12866);
   U2153 : AOI22_X1 port map( A1 => REGISTERS_26_29_port, A2 => n12866, B1 => 
                           REGISTERS_18_29_port, B2 => n12874, ZN => n12256);
   U2154 : NAND4_X1 port map( A1 => n12259, A2 => n12258, A3 => n12257, A4 => 
                           n12256, ZN => n12265);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_30_29_port, A2 => n12941, B1 => 
                           REGISTERS_27_29_port, B2 => n12872, ZN => n12263);
   U2156 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n12938, B1 => 
                           REGISTERS_28_29_port, B2 => n12867, ZN => n12262);
   U2157 : CLKBUF_X1 port map( A => n12865, Z => n12928);
   U2158 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n12928, B1 => 
                           REGISTERS_19_29_port, B2 => n12677, ZN => n12261);
   U2159 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n12930, B1 => 
                           REGISTERS_23_29_port, B2 => n12658, ZN => n12260);
   U2160 : NAND4_X1 port map( A1 => n12263, A2 => n12262, A3 => n12261, A4 => 
                           n12260, ZN => n12264);
   U2161 : NOR2_X1 port map( A1 => n12265, A2 => n12264, ZN => n12277);
   U2162 : AOI22_X1 port map( A1 => REGISTERS_2_29_port, A2 => n12881, B1 => 
                           REGISTERS_6_29_port, B2 => n12883, ZN => n12269);
   U2163 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n12951, B1 => 
                           REGISTERS_7_29_port, B2 => n12961, ZN => n12268);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n12955, B1 => 
                           REGISTERS_4_29_port, B2 => n12913, ZN => n12267);
   U2165 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n12914, B1 => 
                           REGISTERS_1_29_port, B2 => n12884, ZN => n12266);
   U2166 : NAND4_X1 port map( A1 => n12269, A2 => n12268, A3 => n12267, A4 => 
                           n12266, ZN => n12275);
   U2167 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n12952, B1 => 
                           REGISTERS_10_29_port, B2 => n12966, ZN => n12273);
   U2168 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n12955, B1 => 
                           REGISTERS_15_29_port, B2 => n12961, ZN => n12272);
   U2169 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n12963, B1 => 
                           REGISTERS_14_29_port, B2 => n12883, ZN => n12271);
   U2170 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n12914, B1 => 
                           REGISTERS_12_29_port, B2 => n12913, ZN => n12270);
   U2171 : NAND4_X1 port map( A1 => n12273, A2 => n12272, A3 => n12271, A4 => 
                           n12270, ZN => n12274);
   U2172 : AOI22_X1 port map( A1 => n12788, A2 => n12275, B1 => n12811, B2 => 
                           n12274, ZN => n12276);
   U2173 : OAI21_X1 port map( B1 => n12924, B2 => n12277, A => n12276, ZN => 
                           N414);
   U2174 : AOI22_X1 port map( A1 => REGISTERS_22_28_port, A2 => n12944, B1 => 
                           REGISTERS_24_28_port, B2 => n12613, ZN => n12281);
   U2175 : AOI22_X1 port map( A1 => REGISTERS_31_28_port, A2 => n12943, B1 => 
                           REGISTERS_28_28_port, B2 => n12867, ZN => n12280);
   U2176 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n12932, B1 => 
                           REGISTERS_30_28_port, B2 => n12678, ZN => n12279);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n12931, B1 => 
                           REGISTERS_23_28_port, B2 => n12658, ZN => n12278);
   U2178 : NAND4_X1 port map( A1 => n12281, A2 => n12280, A3 => n12279, A4 => 
                           n12278, ZN => n12287);
   U2179 : CLKBUF_X1 port map( A => n12874, Z => n12937);
   U2180 : AOI22_X1 port map( A1 => REGISTERS_18_28_port, A2 => n12937, B1 => 
                           REGISTERS_29_28_port, B2 => n12843, ZN => n12285);
   U2181 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n12902, B1 => 
                           REGISTERS_19_28_port, B2 => n12677, ZN => n12284);
   U2182 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n12873, B1 => 
                           REGISTERS_16_28_port, B2 => n12865, ZN => n12283);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_26_28_port, A2 => n12866, B1 => 
                           REGISTERS_25_28_port, B2 => n12586, ZN => n12282);
   U2184 : NAND4_X1 port map( A1 => n12285, A2 => n12284, A3 => n12283, A4 => 
                           n12282, ZN => n12286);
   U2185 : NOR2_X1 port map( A1 => n12287, A2 => n12286, ZN => n12299);
   U2186 : AOI22_X1 port map( A1 => REGISTERS_7_28_port, A2 => n12953, B1 => 
                           REGISTERS_5_28_port, B2 => n12805, ZN => n12291);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n12955, B1 => 
                           REGISTERS_2_28_port, B2 => n12881, ZN => n12290);
   U2188 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n12882, B1 => 
                           REGISTERS_1_28_port, B2 => n12952, ZN => n12289);
   U2189 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n12914, B1 => 
                           REGISTERS_6_28_port, B2 => n12883, ZN => n12288);
   U2190 : NAND4_X1 port map( A1 => n12291, A2 => n12290, A3 => n12289, A4 => 
                           n12288, ZN => n12297);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n12967, B1 => 
                           REGISTERS_8_28_port, B2 => n12962, ZN => n12295);
   U2192 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n12914, B1 => 
                           REGISTERS_13_28_port, B2 => n12951, ZN => n12294);
   U2193 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n12882, B1 => 
                           REGISTERS_10_28_port, B2 => n12966, ZN => n12293);
   U2194 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n12953, B1 => 
                           REGISTERS_14_28_port, B2 => n12883, ZN => n12292);
   U2195 : NAND4_X1 port map( A1 => n12295, A2 => n12294, A3 => n12293, A4 => 
                           n12292, ZN => n12296);
   U2196 : AOI22_X1 port map( A1 => n12788, A2 => n12297, B1 => n12811, B2 => 
                           n12296, ZN => n12298);
   U2197 : OAI21_X1 port map( B1 => n12924, B2 => n12299, A => n12298, ZN => 
                           N413);
   U2198 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n12942, B1 => 
                           REGISTERS_25_27_port, B2 => n12586, ZN => n12303);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_26_27_port, A2 => n12866, B1 => 
                           REGISTERS_20_27_port, B2 => n12931, ZN => n12302);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_18_27_port, A2 => n12937, B1 => 
                           REGISTERS_22_27_port, B2 => n12944, ZN => n12301);
   U2201 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n12867, B1 => 
                           REGISTERS_23_27_port, B2 => n12658, ZN => n12300);
   U2202 : NAND4_X1 port map( A1 => n12303, A2 => n12302, A3 => n12301, A4 => 
                           n12300, ZN => n12309);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n12872, B1 => 
                           REGISTERS_30_27_port, B2 => n12678, ZN => n12307);
   U2204 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n12930, B1 => 
                           REGISTERS_21_27_port, B2 => n12940, ZN => n12306);
   U2205 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n12928, B1 => 
                           REGISTERS_17_27_port, B2 => n12939, ZN => n12305);
   U2206 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n12943, B1 => 
                           REGISTERS_19_27_port, B2 => n12677, ZN => n12304);
   U2207 : NAND4_X1 port map( A1 => n12307, A2 => n12306, A3 => n12305, A4 => 
                           n12304, ZN => n12308);
   U2208 : NOR2_X1 port map( A1 => n12309, A2 => n12308, ZN => n12321);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_2_27_port, A2 => n12966, B1 => 
                           REGISTERS_6_27_port, B2 => n12883, ZN => n12313);
   U2210 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n12967, B1 => 
                           REGISTERS_4_27_port, B2 => n12913, ZN => n12312);
   U2211 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n12805, B1 => 
                           REGISTERS_3_27_port, B2 => n12960, ZN => n12311);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n12953, B1 => 
                           REGISTERS_0_27_port, B2 => n12962, ZN => n12310);
   U2213 : NAND4_X1 port map( A1 => n12313, A2 => n12312, A3 => n12311, A4 => 
                           n12310, ZN => n12319);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_10_27_port, A2 => n12966, B1 => 
                           REGISTERS_9_27_port, B2 => n12884, ZN => n12317);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n12955, B1 => 
                           REGISTERS_15_27_port, B2 => n12961, ZN => n12316);
   U2216 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n12914, B1 => 
                           REGISTERS_14_27_port, B2 => n12889, ZN => n12315);
   U2217 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n12882, B1 => 
                           REGISTERS_13_27_port, B2 => n12951, ZN => n12314);
   U2218 : NAND4_X1 port map( A1 => n12317, A2 => n12316, A3 => n12315, A4 => 
                           n12314, ZN => n12318);
   U2219 : AOI22_X1 port map( A1 => n12788, A2 => n12319, B1 => n12811, B2 => 
                           n12318, ZN => n12320);
   U2220 : OAI21_X1 port map( B1 => n12924, B2 => n12321, A => n12320, ZN => 
                           N412);
   U2221 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n12931, B1 => 
                           REGISTERS_25_26_port, B2 => n12586, ZN => n12325);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_22_26_port, A2 => n12944, B1 => 
                           REGISTERS_30_26_port, B2 => n12678, ZN => n12324);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n12902, B1 => 
                           REGISTERS_18_26_port, B2 => n12937, ZN => n12323);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n12925, B1 => 
                           REGISTERS_26_26_port, B2 => n12929, ZN => n12322);
   U2225 : NAND4_X1 port map( A1 => n12325, A2 => n12324, A3 => n12323, A4 => 
                           n12322, ZN => n12331);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n12928, B1 => 
                           REGISTERS_23_26_port, B2 => n12658, ZN => n12329);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_31_26_port, A2 => n12943, B1 => 
                           REGISTERS_24_26_port, B2 => n12613, ZN => n12328);
   U2228 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n12873, B1 => 
                           REGISTERS_27_26_port, B2 => n12932, ZN => n12327);
   U2229 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n12926, B1 => 
                           REGISTERS_29_26_port, B2 => n12843, ZN => n12326);
   U2230 : NAND4_X1 port map( A1 => n12329, A2 => n12328, A3 => n12327, A4 => 
                           n12326, ZN => n12330);
   U2231 : NOR2_X1 port map( A1 => n12331, A2 => n12330, ZN => n12343);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n12914, B1 => 
                           REGISTERS_6_26_port, B2 => n12883, ZN => n12335);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n12955, B1 => 
                           REGISTERS_1_26_port, B2 => n12952, ZN => n12334);
   U2234 : CLKBUF_X1 port map( A => n12966, Z => n12954);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_2_26_port, A2 => n12954, B1 => 
                           REGISTERS_4_26_port, B2 => n12913, ZN => n12333);
   U2236 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n12953, B1 => 
                           REGISTERS_5_26_port, B2 => n12805, ZN => n12332);
   U2237 : NAND4_X1 port map( A1 => n12335, A2 => n12334, A3 => n12333, A4 => 
                           n12332, ZN => n12341);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n12952, B1 => 
                           REGISTERS_10_26_port, B2 => n12881, ZN => n12339);
   U2239 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n12953, B1 => 
                           REGISTERS_12_26_port, B2 => n12965, ZN => n12338);
   U2240 : AOI22_X1 port map( A1 => REGISTERS_14_26_port, A2 => n12964, B1 => 
                           REGISTERS_8_26_port, B2 => n12962, ZN => n12337);
   U2241 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n12914, B1 => 
                           REGISTERS_13_26_port, B2 => n12951, ZN => n12336);
   U2242 : NAND4_X1 port map( A1 => n12339, A2 => n12338, A3 => n12337, A4 => 
                           n12336, ZN => n12340);
   U2243 : AOI22_X1 port map( A1 => n12788, A2 => n12341, B1 => n12811, B2 => 
                           n12340, ZN => n12342);
   U2244 : OAI21_X1 port map( B1 => n12924, B2 => n12343, A => n12342, ZN => 
                           N411);
   U2245 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n12872, B1 => 
                           REGISTERS_24_25_port, B2 => n12613, ZN => n12347);
   U2246 : AOI22_X1 port map( A1 => REGISTERS_30_25_port, A2 => n12941, B1 => 
                           REGISTERS_23_25_port, B2 => n12658, ZN => n12346);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n12902, B1 => 
                           REGISTERS_22_25_port, B2 => n12844, ZN => n12345);
   U2248 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n12925, B1 => 
                           REGISTERS_18_25_port, B2 => n12937, ZN => n12344);
   U2249 : NAND4_X1 port map( A1 => n12347, A2 => n12346, A3 => n12345, A4 => 
                           n12344, ZN => n12353);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n12928, B1 => 
                           REGISTERS_29_25_port, B2 => n12843, ZN => n12351);
   U2251 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n12943, B1 => 
                           REGISTERS_28_25_port, B2 => n12867, ZN => n12350);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n12938, B1 => 
                           REGISTERS_20_25_port, B2 => n12771, ZN => n12349);
   U2253 : AOI22_X1 port map( A1 => REGISTERS_26_25_port, A2 => n12866, B1 => 
                           REGISTERS_17_25_port, B2 => n12939, ZN => n12348);
   U2254 : NAND4_X1 port map( A1 => n12351, A2 => n12350, A3 => n12349, A4 => 
                           n12348, ZN => n12352);
   U2255 : NOR2_X1 port map( A1 => n12353, A2 => n12352, ZN => n12365);
   U2256 : AOI22_X1 port map( A1 => REGISTERS_2_25_port, A2 => n12881, B1 => 
                           REGISTERS_3_25_port, B2 => n12960, ZN => n12357);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n12884, B1 => 
                           REGISTERS_4_25_port, B2 => n12913, ZN => n12356);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n12963, B1 => 
                           REGISTERS_7_25_port, B2 => n12961, ZN => n12355);
   U2259 : AOI22_X1 port map( A1 => REGISTERS_6_25_port, A2 => n12964, B1 => 
                           REGISTERS_0_25_port, B2 => n12962, ZN => n12354);
   U2260 : NAND4_X1 port map( A1 => n12357, A2 => n12356, A3 => n12355, A4 => 
                           n12354, ZN => n12363);
   U2261 : AOI22_X1 port map( A1 => REGISTERS_10_25_port, A2 => n12881, B1 => 
                           REGISTERS_11_25_port, B2 => n12960, ZN => n12361);
   U2262 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n12851, B1 => 
                           REGISTERS_8_25_port, B2 => n12915, ZN => n12360);
   U2263 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n12805, B1 => 
                           REGISTERS_14_25_port, B2 => n12889, ZN => n12359);
   U2264 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n12882, B1 => 
                           REGISTERS_9_25_port, B2 => n12884, ZN => n12358);
   U2265 : NAND4_X1 port map( A1 => n12361, A2 => n12360, A3 => n12359, A4 => 
                           n12358, ZN => n12362);
   U2266 : AOI22_X1 port map( A1 => n12788, A2 => n12363, B1 => n12811, B2 => 
                           n12362, ZN => n12364);
   U2267 : OAI21_X1 port map( B1 => n12924, B2 => n12365, A => n12364, ZN => 
                           N410);
   U2268 : AOI22_X1 port map( A1 => REGISTERS_19_24_port, A2 => n12925, B1 => 
                           REGISTERS_27_24_port, B2 => n12932, ZN => n12369);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n12874, B1 => 
                           REGISTERS_22_24_port, B2 => n12844, ZN => n12368);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n12927, B1 => 
                           REGISTERS_21_24_port, B2 => n12940, ZN => n12367);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n12930, B1 => 
                           REGISTERS_25_24_port, B2 => n12586, ZN => n12366);
   U2272 : NAND4_X1 port map( A1 => n12369, A2 => n12368, A3 => n12367, A4 => 
                           n12366, ZN => n12375);
   U2273 : AOI22_X1 port map( A1 => REGISTERS_26_24_port, A2 => n12929, B1 => 
                           REGISTERS_20_24_port, B2 => n12771, ZN => n12373);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n12873, B1 => 
                           REGISTERS_30_24_port, B2 => n12678, ZN => n12372);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n12867, B1 => 
                           REGISTERS_24_24_port, B2 => n12613, ZN => n12371);
   U2276 : AOI22_X1 port map( A1 => REGISTERS_31_24_port, A2 => n12943, B1 => 
                           REGISTERS_16_24_port, B2 => n12928, ZN => n12370);
   U2277 : NAND4_X1 port map( A1 => n12373, A2 => n12372, A3 => n12371, A4 => 
                           n12370, ZN => n12374);
   U2278 : NOR2_X1 port map( A1 => n12375, A2 => n12374, ZN => n12387);
   U2279 : AOI22_X1 port map( A1 => REGISTERS_2_24_port, A2 => n12966, B1 => 
                           REGISTERS_3_24_port, B2 => n12960, ZN => n12379);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n12963, B1 => 
                           REGISTERS_1_24_port, B2 => n12884, ZN => n12378);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n12955, B1 => 
                           REGISTERS_7_24_port, B2 => n12851, ZN => n12377);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n12882, B1 => 
                           REGISTERS_6_24_port, B2 => n12883, ZN => n12376);
   U2283 : NAND4_X1 port map( A1 => n12379, A2 => n12378, A3 => n12377, A4 => 
                           n12376, ZN => n12385);
   U2284 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n12965, B1 => 
                           REGISTERS_11_24_port, B2 => n12852, ZN => n12383);
   U2285 : AOI22_X1 port map( A1 => REGISTERS_15_24_port, A2 => n12961, B1 => 
                           REGISTERS_10_24_port, B2 => n12954, ZN => n12382);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n12951, B1 => 
                           REGISTERS_9_24_port, B2 => n12952, ZN => n12381);
   U2287 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n12962, B1 => 
                           REGISTERS_14_24_port, B2 => n12889, ZN => n12380);
   U2288 : NAND4_X1 port map( A1 => n12383, A2 => n12382, A3 => n12381, A4 => 
                           n12380, ZN => n12384);
   U2289 : AOI22_X1 port map( A1 => n12788, A2 => n12385, B1 => n12811, B2 => 
                           n12384, ZN => n12386);
   U2290 : OAI21_X1 port map( B1 => n12924, B2 => n12387, A => n12386, ZN => 
                           N409);
   U2291 : AOI22_X1 port map( A1 => REGISTERS_23_23_port, A2 => n12927, B1 => 
                           REGISTERS_28_23_port, B2 => n12926, ZN => n12391);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n12873, B1 => 
                           REGISTERS_24_23_port, B2 => n12613, ZN => n12390);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_26_23_port, A2 => n12866, B1 => 
                           REGISTERS_29_23_port, B2 => n12930, ZN => n12389);
   U2294 : AOI22_X1 port map( A1 => REGISTERS_27_23_port, A2 => n12872, B1 => 
                           REGISTERS_22_23_port, B2 => n12944, ZN => n12388);
   U2295 : NAND4_X1 port map( A1 => n12391, A2 => n12390, A3 => n12389, A4 => 
                           n12388, ZN => n12397);
   U2296 : AOI22_X1 port map( A1 => REGISTERS_18_23_port, A2 => n12874, B1 => 
                           REGISTERS_20_23_port, B2 => n12771, ZN => n12395);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_30_23_port, A2 => n12941, B1 => 
                           REGISTERS_31_23_port, B2 => n12838, ZN => n12394);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n12928, B1 => 
                           REGISTERS_21_23_port, B2 => n12940, ZN => n12393);
   U2299 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n12938, B1 => 
                           REGISTERS_19_23_port, B2 => n12677, ZN => n12392);
   U2300 : NAND4_X1 port map( A1 => n12395, A2 => n12394, A3 => n12393, A4 => 
                           n12392, ZN => n12396);
   U2301 : NOR2_X1 port map( A1 => n12397, A2 => n12396, ZN => n12409);
   U2302 : AOI22_X1 port map( A1 => REGISTERS_2_23_port, A2 => n12966, B1 => 
                           REGISTERS_6_23_port, B2 => n12883, ZN => n12401);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n12915, B1 => 
                           REGISTERS_3_23_port, B2 => n12914, ZN => n12400);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n12805, B1 => 
                           REGISTERS_1_23_port, B2 => n12884, ZN => n12399);
   U2305 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n12882, B1 => 
                           REGISTERS_7_23_port, B2 => n12961, ZN => n12398);
   U2306 : NAND4_X1 port map( A1 => n12401, A2 => n12400, A3 => n12399, A4 => 
                           n12398, ZN => n12407);
   U2307 : AOI22_X1 port map( A1 => REGISTERS_14_23_port, A2 => n12964, B1 => 
                           REGISTERS_11_23_port, B2 => n12852, ZN => n12405);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n12955, B1 => 
                           REGISTERS_13_23_port, B2 => n12951, ZN => n12404);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n12953, B1 => 
                           REGISTERS_9_23_port, B2 => n12967, ZN => n12403);
   U2310 : AOI22_X1 port map( A1 => REGISTERS_10_23_port, A2 => n12966, B1 => 
                           REGISTERS_12_23_port, B2 => n12965, ZN => n12402);
   U2311 : NAND4_X1 port map( A1 => n12405, A2 => n12404, A3 => n12403, A4 => 
                           n12402, ZN => n12406);
   U2312 : AOI22_X1 port map( A1 => n12788, A2 => n12407, B1 => n12811, B2 => 
                           n12406, ZN => n12408);
   U2313 : OAI21_X1 port map( B1 => n12978, B2 => n12409, A => n12408, ZN => 
                           N408);
   U2314 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n12928, B1 => 
                           REGISTERS_19_22_port, B2 => n12677, ZN => n12413);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n12902, B1 => 
                           REGISTERS_17_22_port, B2 => n12873, ZN => n12412);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_22_22_port, A2 => n12944, B1 => 
                           REGISTERS_24_22_port, B2 => n12613, ZN => n12411);
   U2317 : AOI22_X1 port map( A1 => REGISTERS_27_22_port, A2 => n12932, B1 => 
                           REGISTERS_26_22_port, B2 => n12866, ZN => n12410);
   U2318 : NAND4_X1 port map( A1 => n12413, A2 => n12412, A3 => n12411, A4 => 
                           n12410, ZN => n12419);
   U2319 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n12930, B1 => 
                           REGISTERS_28_22_port, B2 => n12926, ZN => n12417);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_30_22_port, A2 => n12941, B1 => 
                           REGISTERS_25_22_port, B2 => n12586, ZN => n12416);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n12931, B1 => 
                           REGISTERS_31_22_port, B2 => n12838, ZN => n12415);
   U2322 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n12927, B1 => 
                           REGISTERS_18_22_port, B2 => n12874, ZN => n12414);
   U2323 : NAND4_X1 port map( A1 => n12417, A2 => n12416, A3 => n12415, A4 => 
                           n12414, ZN => n12418);
   U2324 : NOR2_X1 port map( A1 => n12419, A2 => n12418, ZN => n12431);
   U2325 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n12965, B1 => 
                           REGISTERS_3_22_port, B2 => n12960, ZN => n12423);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n12953, B1 => 
                           REGISTERS_6_22_port, B2 => n12889, ZN => n12422);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n12884, B1 => 
                           REGISTERS_0_22_port, B2 => n12962, ZN => n12421);
   U2328 : AOI22_X1 port map( A1 => REGISTERS_2_22_port, A2 => n12966, B1 => 
                           REGISTERS_5_22_port, B2 => n12963, ZN => n12420);
   U2329 : NAND4_X1 port map( A1 => n12423, A2 => n12422, A3 => n12421, A4 => 
                           n12420, ZN => n12429);
   U2330 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n12952, B1 => 
                           REGISTERS_14_22_port, B2 => n12883, ZN => n12427);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n12805, B1 => 
                           REGISTERS_10_22_port, B2 => n12881, ZN => n12426);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n12851, B1 => 
                           REGISTERS_8_22_port, B2 => n12915, ZN => n12425);
   U2333 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n12882, B1 => 
                           REGISTERS_11_22_port, B2 => n12852, ZN => n12424);
   U2334 : NAND4_X1 port map( A1 => n12427, A2 => n12426, A3 => n12425, A4 => 
                           n12424, ZN => n12428);
   U2335 : AOI22_X1 port map( A1 => n12788, A2 => n12429, B1 => n12811, B2 => 
                           n12428, ZN => n12430);
   U2336 : OAI21_X1 port map( B1 => n12978, B2 => n12431, A => n12430, ZN => 
                           N407);
   U2337 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n12942, B1 => 
                           REGISTERS_27_21_port, B2 => n12932, ZN => n12435);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_18_21_port, A2 => n12874, B1 => 
                           REGISTERS_21_21_port, B2 => n12902, ZN => n12434);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n12930, B1 => 
                           REGISTERS_31_21_port, B2 => n12838, ZN => n12433);
   U2340 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n12873, B1 => 
                           REGISTERS_16_21_port, B2 => n12928, ZN => n12432);
   U2341 : NAND4_X1 port map( A1 => n12435, A2 => n12434, A3 => n12433, A4 => 
                           n12432, ZN => n12441);
   U2342 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n12944, B1 => 
                           REGISTERS_28_21_port, B2 => n12926, ZN => n12439);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n12931, B1 => 
                           REGISTERS_30_21_port, B2 => n12678, ZN => n12438);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n12925, B1 => 
                           REGISTERS_26_21_port, B2 => n12866, ZN => n12437);
   U2345 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n12938, B1 => 
                           REGISTERS_23_21_port, B2 => n12658, ZN => n12436);
   U2346 : NAND4_X1 port map( A1 => n12439, A2 => n12438, A3 => n12437, A4 => 
                           n12436, ZN => n12440);
   U2347 : NOR2_X1 port map( A1 => n12441, A2 => n12440, ZN => n12453);
   U2348 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n12955, B1 => 
                           REGISTERS_6_21_port, B2 => n12889, ZN => n12445);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_3_21_port, A2 => n12914, B1 => 
                           REGISTERS_7_21_port, B2 => n12851, ZN => n12444);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n12963, B1 => 
                           REGISTERS_1_21_port, B2 => n12952, ZN => n12443);
   U2351 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n12882, B1 => 
                           REGISTERS_2_21_port, B2 => n12966, ZN => n12442);
   U2352 : NAND4_X1 port map( A1 => n12445, A2 => n12444, A3 => n12443, A4 => 
                           n12442, ZN => n12451);
   U2353 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n12915, B1 => 
                           REGISTERS_14_21_port, B2 => n12883, ZN => n12449);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n12951, B1 => 
                           REGISTERS_12_21_port, B2 => n12913, ZN => n12448);
   U2355 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n12953, B1 => 
                           REGISTERS_9_21_port, B2 => n12884, ZN => n12447);
   U2356 : AOI22_X1 port map( A1 => REGISTERS_10_21_port, A2 => n12954, B1 => 
                           REGISTERS_11_21_port, B2 => n12960, ZN => n12446);
   U2357 : NAND4_X1 port map( A1 => n12449, A2 => n12448, A3 => n12447, A4 => 
                           n12446, ZN => n12450);
   U2358 : AOI22_X1 port map( A1 => n12788, A2 => n12451, B1 => n12811, B2 => 
                           n12450, ZN => n12452);
   U2359 : OAI21_X1 port map( B1 => n12978, B2 => n12453, A => n12452, ZN => 
                           N406);
   U2360 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n12942, B1 => 
                           REGISTERS_30_20_port, B2 => n12678, ZN => n12457);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n12932, B1 => 
                           REGISTERS_18_20_port, B2 => n12937, ZN => n12456);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_31_20_port, A2 => n12838, B1 => 
                           REGISTERS_25_20_port, B2 => n12586, ZN => n12455);
   U2363 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n12902, B1 => 
                           REGISTERS_23_20_port, B2 => n12658, ZN => n12454);
   U2364 : NAND4_X1 port map( A1 => n12457, A2 => n12456, A3 => n12455, A4 => 
                           n12454, ZN => n12463);
   U2365 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n12930, B1 => 
                           REGISTERS_22_20_port, B2 => n12844, ZN => n12461);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_26_20_port, A2 => n12929, B1 => 
                           REGISTERS_16_20_port, B2 => n12928, ZN => n12460);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n12939, B1 => 
                           REGISTERS_28_20_port, B2 => n12926, ZN => n12459);
   U2368 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n12677, B1 => 
                           REGISTERS_20_20_port, B2 => n12771, ZN => n12458);
   U2369 : NAND4_X1 port map( A1 => n12461, A2 => n12460, A3 => n12459, A4 => 
                           n12458, ZN => n12462);
   U2370 : NOR2_X1 port map( A1 => n12463, A2 => n12462, ZN => n12475);
   U2371 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n12805, B1 => 
                           REGISTERS_1_20_port, B2 => n12967, ZN => n12467);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n12955, B1 => 
                           REGISTERS_4_20_port, B2 => n12965, ZN => n12466);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_2_20_port, A2 => n12966, B1 => 
                           REGISTERS_7_20_port, B2 => n12961, ZN => n12465);
   U2374 : AOI22_X1 port map( A1 => REGISTERS_3_20_port, A2 => n12852, B1 => 
                           REGISTERS_6_20_port, B2 => n12889, ZN => n12464);
   U2375 : NAND4_X1 port map( A1 => n12467, A2 => n12466, A3 => n12465, A4 => 
                           n12464, ZN => n12473);
   U2376 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n12914, B1 => 
                           REGISTERS_12_20_port, B2 => n12913, ZN => n12471);
   U2377 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n12951, B1 => 
                           REGISTERS_14_20_port, B2 => n12889, ZN => n12470);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_10_20_port, A2 => n12954, B1 => 
                           REGISTERS_15_20_port, B2 => n12851, ZN => n12469);
   U2379 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n12962, B1 => 
                           REGISTERS_9_20_port, B2 => n12952, ZN => n12468);
   U2380 : NAND4_X1 port map( A1 => n12471, A2 => n12470, A3 => n12469, A4 => 
                           n12468, ZN => n12472);
   U2381 : AOI22_X1 port map( A1 => n12788, A2 => n12473, B1 => n12973, B2 => 
                           n12472, ZN => n12474);
   U2382 : OAI21_X1 port map( B1 => n12978, B2 => n12475, A => n12474, ZN => 
                           N405);
   U2383 : AOI22_X1 port map( A1 => REGISTERS_31_19_port, A2 => n12943, B1 => 
                           REGISTERS_21_19_port, B2 => n12940, ZN => n12479);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n12930, B1 => 
                           REGISTERS_16_19_port, B2 => n12928, ZN => n12478);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n12927, B1 => 
                           REGISTERS_28_19_port, B2 => n12926, ZN => n12477);
   U2386 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n12942, B1 => 
                           REGISTERS_26_19_port, B2 => n12866, ZN => n12476);
   U2387 : NAND4_X1 port map( A1 => n12479, A2 => n12478, A3 => n12477, A4 => 
                           n12476, ZN => n12485);
   U2388 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n12939, B1 => 
                           REGISTERS_22_19_port, B2 => n12844, ZN => n12483);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_30_19_port, A2 => n12941, B1 => 
                           REGISTERS_27_19_port, B2 => n12932, ZN => n12482);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n12586, B1 => 
                           REGISTERS_18_19_port, B2 => n12937, ZN => n12481);
   U2391 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n12931, B1 => 
                           REGISTERS_19_19_port, B2 => n12677, ZN => n12480);
   U2392 : NAND4_X1 port map( A1 => n12483, A2 => n12482, A3 => n12481, A4 => 
                           n12480, ZN => n12484);
   U2393 : NOR2_X1 port map( A1 => n12485, A2 => n12484, ZN => n12497);
   U2394 : CLKBUF_X1 port map( A => n12975, Z => n12813);
   U2395 : AOI22_X1 port map( A1 => REGISTERS_6_19_port, A2 => n12883, B1 => 
                           REGISTERS_1_19_port, B2 => n12952, ZN => n12489);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n12963, B1 => 
                           REGISTERS_0_19_port, B2 => n12962, ZN => n12488);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n12851, B1 => 
                           REGISTERS_2_19_port, B2 => n12966, ZN => n12487);
   U2398 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n12882, B1 => 
                           REGISTERS_3_19_port, B2 => n12852, ZN => n12486);
   U2399 : NAND4_X1 port map( A1 => n12489, A2 => n12488, A3 => n12487, A4 => 
                           n12486, ZN => n12495);
   U2400 : AOI22_X1 port map( A1 => REGISTERS_10_19_port, A2 => n12881, B1 => 
                           REGISTERS_8_19_port, B2 => n12915, ZN => n12493);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n12852, B1 => 
                           REGISTERS_12_19_port, B2 => n12965, ZN => n12492);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n12967, B1 => 
                           REGISTERS_15_19_port, B2 => n12961, ZN => n12491);
   U2403 : AOI22_X1 port map( A1 => REGISTERS_14_19_port, A2 => n12964, B1 => 
                           REGISTERS_13_19_port, B2 => n12805, ZN => n12490);
   U2404 : NAND4_X1 port map( A1 => n12493, A2 => n12492, A3 => n12491, A4 => 
                           n12490, ZN => n12494);
   U2405 : AOI22_X1 port map( A1 => n12813, A2 => n12495, B1 => n12811, B2 => 
                           n12494, ZN => n12496);
   U2406 : OAI21_X1 port map( B1 => n12978, B2 => n12497, A => n12496, ZN => 
                           N404);
   U2407 : AOI22_X1 port map( A1 => REGISTERS_26_18_port, A2 => n12866, B1 => 
                           REGISTERS_22_18_port, B2 => n12844, ZN => n12501);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n12771, B1 => 
                           REGISTERS_21_18_port, B2 => n12902, ZN => n12500);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n12932, B1 => 
                           REGISTERS_23_18_port, B2 => n12927, ZN => n12499);
   U2410 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n12928, B1 => 
                           REGISTERS_31_18_port, B2 => n12838, ZN => n12498);
   U2411 : NAND4_X1 port map( A1 => n12501, A2 => n12500, A3 => n12499, A4 => 
                           n12498, ZN => n12507);
   U2412 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n12677, B1 => 
                           REGISTERS_28_18_port, B2 => n12926, ZN => n12505);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_30_18_port, A2 => n12941, B1 => 
                           REGISTERS_18_18_port, B2 => n12937, ZN => n12504);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n12613, B1 => 
                           REGISTERS_25_18_port, B2 => n12586, ZN => n12503);
   U2415 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n12930, B1 => 
                           REGISTERS_17_18_port, B2 => n12939, ZN => n12502);
   U2416 : NAND4_X1 port map( A1 => n12505, A2 => n12504, A3 => n12503, A4 => 
                           n12502, ZN => n12506);
   U2417 : NOR2_X1 port map( A1 => n12507, A2 => n12506, ZN => n12519);
   U2418 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n12961, B1 => 
                           REGISTERS_2_18_port, B2 => n12954, ZN => n12511);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n12805, B1 => 
                           REGISTERS_4_18_port, B2 => n12913, ZN => n12510);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n12914, B1 => 
                           REGISTERS_1_18_port, B2 => n12952, ZN => n12509);
   U2421 : AOI22_X1 port map( A1 => REGISTERS_6_18_port, A2 => n12964, B1 => 
                           REGISTERS_0_18_port, B2 => n12962, ZN => n12508);
   U2422 : NAND4_X1 port map( A1 => n12511, A2 => n12510, A3 => n12509, A4 => 
                           n12508, ZN => n12517);
   U2423 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n12951, B1 => 
                           REGISTERS_9_18_port, B2 => n12952, ZN => n12515);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n12913, B1 => 
                           REGISTERS_10_18_port, B2 => n12954, ZN => n12514);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n12953, B1 => 
                           REGISTERS_14_18_port, B2 => n12883, ZN => n12513);
   U2426 : AOI22_X1 port map( A1 => REGISTERS_11_18_port, A2 => n12960, B1 => 
                           REGISTERS_8_18_port, B2 => n12915, ZN => n12512);
   U2427 : NAND4_X1 port map( A1 => n12515, A2 => n12514, A3 => n12513, A4 => 
                           n12512, ZN => n12516);
   U2428 : AOI22_X1 port map( A1 => n12813, A2 => n12517, B1 => n12811, B2 => 
                           n12516, ZN => n12518);
   U2429 : OAI21_X1 port map( B1 => n12978, B2 => n12519, A => n12518, ZN => 
                           N403);
   U2430 : AOI22_X1 port map( A1 => REGISTERS_26_17_port, A2 => n12866, B1 => 
                           REGISTERS_27_17_port, B2 => n12932, ZN => n12523);
   U2431 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n12930, B1 => 
                           REGISTERS_17_17_port, B2 => n12873, ZN => n12522);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n12613, B1 => 
                           REGISTERS_18_17_port, B2 => n12937, ZN => n12521);
   U2433 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n12927, B1 => 
                           REGISTERS_31_17_port, B2 => n12838, ZN => n12520);
   U2434 : NAND4_X1 port map( A1 => n12523, A2 => n12522, A3 => n12521, A4 => 
                           n12520, ZN => n12529);
   U2435 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n12865, B1 => 
                           REGISTERS_21_17_port, B2 => n12902, ZN => n12527);
   U2436 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n12586, B1 => 
                           REGISTERS_22_17_port, B2 => n12844, ZN => n12526);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_30_17_port, A2 => n12941, B1 => 
                           REGISTERS_20_17_port, B2 => n12771, ZN => n12525);
   U2438 : AOI22_X1 port map( A1 => REGISTERS_19_17_port, A2 => n12925, B1 => 
                           REGISTERS_28_17_port, B2 => n12926, ZN => n12524);
   U2439 : NAND4_X1 port map( A1 => n12527, A2 => n12526, A3 => n12525, A4 => 
                           n12524, ZN => n12528);
   U2440 : NOR2_X1 port map( A1 => n12529, A2 => n12528, ZN => n12541);
   U2441 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n12955, B1 => 
                           REGISTERS_2_17_port, B2 => n12966, ZN => n12533);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n12889, B1 => 
                           REGISTERS_3_17_port, B2 => n12960, ZN => n12532);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n12913, B1 => 
                           REGISTERS_7_17_port, B2 => n12851, ZN => n12531);
   U2444 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n12963, B1 => 
                           REGISTERS_1_17_port, B2 => n12967, ZN => n12530);
   U2445 : NAND4_X1 port map( A1 => n12533, A2 => n12532, A3 => n12531, A4 => 
                           n12530, ZN => n12539);
   U2446 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n12881, B1 => 
                           REGISTERS_9_17_port, B2 => n12884, ZN => n12537);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n12851, B1 => 
                           REGISTERS_12_17_port, B2 => n12965, ZN => n12536);
   U2448 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n12915, B1 => 
                           REGISTERS_13_17_port, B2 => n12951, ZN => n12535);
   U2449 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n12960, B1 => 
                           REGISTERS_14_17_port, B2 => n12889, ZN => n12534);
   U2450 : NAND4_X1 port map( A1 => n12537, A2 => n12536, A3 => n12535, A4 => 
                           n12534, ZN => n12538);
   U2451 : AOI22_X1 port map( A1 => n12813, A2 => n12539, B1 => n12811, B2 => 
                           n12538, ZN => n12540);
   U2452 : OAI21_X1 port map( B1 => n12978, B2 => n12541, A => n12540, ZN => 
                           N402);
   U2453 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n12865, B1 => 
                           REGISTERS_22_16_port, B2 => n12844, ZN => n12545);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n12902, B1 => 
                           REGISTERS_24_16_port, B2 => n12613, ZN => n12544);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n12658, B1 => 
                           REGISTERS_31_16_port, B2 => n12838, ZN => n12543);
   U2456 : AOI22_X1 port map( A1 => REGISTERS_18_16_port, A2 => n12937, B1 => 
                           REGISTERS_17_16_port, B2 => n12873, ZN => n12542);
   U2457 : NAND4_X1 port map( A1 => n12545, A2 => n12544, A3 => n12543, A4 => 
                           n12542, ZN => n12551);
   U2458 : AOI22_X1 port map( A1 => REGISTERS_26_16_port, A2 => n12866, B1 => 
                           REGISTERS_29_16_port, B2 => n12843, ZN => n12549);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_30_16_port, A2 => n12678, B1 => 
                           REGISTERS_20_16_port, B2 => n12771, ZN => n12548);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n12932, B1 => 
                           REGISTERS_25_16_port, B2 => n12938, ZN => n12547);
   U2461 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n12926, B1 => 
                           REGISTERS_19_16_port, B2 => n12677, ZN => n12546);
   U2462 : NAND4_X1 port map( A1 => n12549, A2 => n12548, A3 => n12547, A4 => 
                           n12546, ZN => n12550);
   U2463 : NOR2_X1 port map( A1 => n12551, A2 => n12550, ZN => n12563);
   U2464 : AOI22_X1 port map( A1 => REGISTERS_2_16_port, A2 => n12954, B1 => 
                           REGISTERS_5_16_port, B2 => n12951, ZN => n12555);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n12884, B1 => 
                           REGISTERS_3_16_port, B2 => n12852, ZN => n12554);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n12882, B1 => 
                           REGISTERS_7_16_port, B2 => n12961, ZN => n12553);
   U2467 : AOI22_X1 port map( A1 => REGISTERS_6_16_port, A2 => n12883, B1 => 
                           REGISTERS_0_16_port, B2 => n12962, ZN => n12552);
   U2468 : NAND4_X1 port map( A1 => n12555, A2 => n12554, A3 => n12553, A4 => 
                           n12552, ZN => n12561);
   U2469 : AOI22_X1 port map( A1 => REGISTERS_14_16_port, A2 => n12964, B1 => 
                           REGISTERS_11_16_port, B2 => n12960, ZN => n12559);
   U2470 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n12966, B1 => 
                           REGISTERS_8_16_port, B2 => n12915, ZN => n12558);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n12913, B1 => 
                           REGISTERS_9_16_port, B2 => n12952, ZN => n12557);
   U2472 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n12961, B1 => 
                           REGISTERS_13_16_port, B2 => n12951, ZN => n12556);
   U2473 : NAND4_X1 port map( A1 => n12559, A2 => n12558, A3 => n12557, A4 => 
                           n12556, ZN => n12560);
   U2474 : AOI22_X1 port map( A1 => n12813, A2 => n12561, B1 => n12811, B2 => 
                           n12560, ZN => n12562);
   U2475 : OAI21_X1 port map( B1 => n12978, B2 => n12563, A => n12562, ZN => 
                           N401);
   U2476 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n12942, B1 => 
                           REGISTERS_28_15_port, B2 => n12926, ZN => n12567);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_30_15_port, A2 => n12678, B1 => 
                           REGISTERS_17_15_port, B2 => n12873, ZN => n12566);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n12865, B1 => 
                           REGISTERS_20_15_port, B2 => n12771, ZN => n12565);
   U2479 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n12838, B1 => 
                           REGISTERS_27_15_port, B2 => n12932, ZN => n12564);
   U2480 : NAND4_X1 port map( A1 => n12567, A2 => n12566, A3 => n12565, A4 => 
                           n12564, ZN => n12573);
   U2481 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n12843, B1 => 
                           REGISTERS_26_15_port, B2 => n12866, ZN => n12571);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n12940, B1 => 
                           REGISTERS_18_15_port, B2 => n12937, ZN => n12570);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n12925, B1 => 
                           REGISTERS_23_15_port, B2 => n12927, ZN => n12569);
   U2484 : AOI22_X1 port map( A1 => REGISTERS_22_15_port, A2 => n12844, B1 => 
                           REGISTERS_25_15_port, B2 => n12938, ZN => n12568);
   U2485 : NAND4_X1 port map( A1 => n12571, A2 => n12570, A3 => n12569, A4 => 
                           n12568, ZN => n12572);
   U2486 : NOR2_X1 port map( A1 => n12573, A2 => n12572, ZN => n12585);
   U2487 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n12851, B1 => 
                           REGISTERS_1_15_port, B2 => n12967, ZN => n12577);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_2_15_port, A2 => n12881, B1 => 
                           REGISTERS_3_15_port, B2 => n12852, ZN => n12576);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n12805, B1 => 
                           REGISTERS_0_15_port, B2 => n12962, ZN => n12575);
   U2490 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n12882, B1 => 
                           REGISTERS_6_15_port, B2 => n12883, ZN => n12574);
   U2491 : NAND4_X1 port map( A1 => n12577, A2 => n12576, A3 => n12575, A4 => 
                           n12574, ZN => n12583);
   U2492 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n12953, B1 => 
                           REGISTERS_11_15_port, B2 => n12852, ZN => n12581);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n12951, B1 => 
                           REGISTERS_8_15_port, B2 => n12915, ZN => n12580);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_14_15_port, A2 => n12883, B1 => 
                           REGISTERS_9_15_port, B2 => n12967, ZN => n12579);
   U2495 : AOI22_X1 port map( A1 => REGISTERS_10_15_port, A2 => n12954, B1 => 
                           REGISTERS_12_15_port, B2 => n12913, ZN => n12578);
   U2496 : NAND4_X1 port map( A1 => n12581, A2 => n12580, A3 => n12579, A4 => 
                           n12578, ZN => n12582);
   U2497 : AOI22_X1 port map( A1 => n12813, A2 => n12583, B1 => n12811, B2 => 
                           n12582, ZN => n12584);
   U2498 : OAI21_X1 port map( B1 => n12924, B2 => n12585, A => n12584, ZN => 
                           N400);
   U2499 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n12931, B1 => 
                           REGISTERS_21_14_port, B2 => n12902, ZN => n12590);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n12613, B1 => 
                           REGISTERS_31_14_port, B2 => n12838, ZN => n12589);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n12586, B1 => 
                           REGISTERS_28_14_port, B2 => n12926, ZN => n12588);
   U2502 : AOI22_X1 port map( A1 => REGISTERS_23_14_port, A2 => n12658, B1 => 
                           REGISTERS_22_14_port, B2 => n12844, ZN => n12587);
   U2503 : NAND4_X1 port map( A1 => n12590, A2 => n12589, A3 => n12588, A4 => 
                           n12587, ZN => n12596);
   U2504 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n12843, B1 => 
                           REGISTERS_27_14_port, B2 => n12932, ZN => n12594);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n12928, B1 => 
                           REGISTERS_17_14_port, B2 => n12873, ZN => n12593);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_30_14_port, A2 => n12678, B1 => 
                           REGISTERS_26_14_port, B2 => n12866, ZN => n12592);
   U2507 : AOI22_X1 port map( A1 => REGISTERS_18_14_port, A2 => n12937, B1 => 
                           REGISTERS_19_14_port, B2 => n12677, ZN => n12591);
   U2508 : NAND4_X1 port map( A1 => n12594, A2 => n12593, A3 => n12592, A4 => 
                           n12591, ZN => n12595);
   U2509 : NOR2_X1 port map( A1 => n12596, A2 => n12595, ZN => n12608);
   U2510 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n12955, B1 => 
                           REGISTERS_2_14_port, B2 => n12881, ZN => n12600);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n12851, B1 => 
                           REGISTERS_1_14_port, B2 => n12884, ZN => n12599);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n12963, B1 => 
                           REGISTERS_3_14_port, B2 => n12960, ZN => n12598);
   U2513 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n12965, B1 => 
                           REGISTERS_6_14_port, B2 => n12889, ZN => n12597);
   U2514 : NAND4_X1 port map( A1 => n12600, A2 => n12599, A3 => n12598, A4 => 
                           n12597, ZN => n12606);
   U2515 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n12913, B1 => 
                           REGISTERS_13_14_port, B2 => n12805, ZN => n12604);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_14_14_port, A2 => n12889, B1 => 
                           REGISTERS_15_14_port, B2 => n12851, ZN => n12603);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_10_14_port, A2 => n12966, B1 => 
                           REGISTERS_11_14_port, B2 => n12852, ZN => n12602);
   U2518 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n12962, B1 => 
                           REGISTERS_9_14_port, B2 => n12884, ZN => n12601);
   U2519 : NAND4_X1 port map( A1 => n12604, A2 => n12603, A3 => n12602, A4 => 
                           n12601, ZN => n12605);
   U2520 : AOI22_X1 port map( A1 => n12813, A2 => n12606, B1 => n12811, B2 => 
                           n12605, ZN => n12607);
   U2521 : OAI21_X1 port map( B1 => n12978, B2 => n12608, A => n12607, ZN => 
                           N399);
   U2522 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n12928, B1 => 
                           REGISTERS_26_13_port, B2 => n12866, ZN => n12612);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n12771, B1 => 
                           REGISTERS_23_13_port, B2 => n12927, ZN => n12611);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_30_13_port, A2 => n12941, B1 => 
                           REGISTERS_27_13_port, B2 => n12932, ZN => n12610);
   U2525 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n12940, B1 => 
                           REGISTERS_17_13_port, B2 => n12873, ZN => n12609);
   U2526 : NAND4_X1 port map( A1 => n12612, A2 => n12611, A3 => n12610, A4 => 
                           n12609, ZN => n12619);
   U2527 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n12926, B1 => 
                           REGISTERS_24_13_port, B2 => n12613, ZN => n12617);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n12925, B1 => 
                           REGISTERS_18_13_port, B2 => n12937, ZN => n12616);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_31_13_port, A2 => n12943, B1 => 
                           REGISTERS_25_13_port, B2 => n12938, ZN => n12615);
   U2530 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n12843, B1 => 
                           REGISTERS_22_13_port, B2 => n12944, ZN => n12614);
   U2531 : NAND4_X1 port map( A1 => n12617, A2 => n12616, A3 => n12615, A4 => 
                           n12614, ZN => n12618);
   U2532 : NOR2_X1 port map( A1 => n12619, A2 => n12618, ZN => n12631);
   U2533 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n12805, B1 => 
                           REGISTERS_3_13_port, B2 => n12960, ZN => n12623);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n12961, B1 => 
                           REGISTERS_4_13_port, B2 => n12965, ZN => n12622);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n12955, B1 => 
                           REGISTERS_6_13_port, B2 => n12883, ZN => n12621);
   U2536 : AOI22_X1 port map( A1 => REGISTERS_2_13_port, A2 => n12881, B1 => 
                           REGISTERS_1_13_port, B2 => n12884, ZN => n12620);
   U2537 : NAND4_X1 port map( A1 => n12623, A2 => n12622, A3 => n12621, A4 => 
                           n12620, ZN => n12629);
   U2538 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n12963, B1 => 
                           REGISTERS_11_13_port, B2 => n12852, ZN => n12627);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n12913, B1 => 
                           REGISTERS_8_13_port, B2 => n12915, ZN => n12626);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n12953, B1 => 
                           REGISTERS_10_13_port, B2 => n12966, ZN => n12625);
   U2541 : AOI22_X1 port map( A1 => REGISTERS_14_13_port, A2 => n12889, B1 => 
                           REGISTERS_9_13_port, B2 => n12967, ZN => n12624);
   U2542 : NAND4_X1 port map( A1 => n12627, A2 => n12626, A3 => n12625, A4 => 
                           n12624, ZN => n12628);
   U2543 : AOI22_X1 port map( A1 => n12813, A2 => n12629, B1 => n12811, B2 => 
                           n12628, ZN => n12630);
   U2544 : OAI21_X1 port map( B1 => n12924, B2 => n12631, A => n12630, ZN => 
                           N398);
   U2545 : AOI22_X1 port map( A1 => REGISTERS_23_12_port, A2 => n12927, B1 => 
                           REGISTERS_30_12_port, B2 => n12678, ZN => n12635);
   U2546 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n12939, B1 => 
                           REGISTERS_31_12_port, B2 => n12838, ZN => n12634);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n12938, B1 => 
                           REGISTERS_19_12_port, B2 => n12925, ZN => n12633);
   U2548 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n12926, B1 => 
                           REGISTERS_26_12_port, B2 => n12929, ZN => n12632);
   U2549 : NAND4_X1 port map( A1 => n12635, A2 => n12634, A3 => n12633, A4 => 
                           n12632, ZN => n12641);
   U2550 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n12928, B1 => 
                           REGISTERS_29_12_port, B2 => n12930, ZN => n12639);
   U2551 : AOI22_X1 port map( A1 => REGISTERS_18_12_port, A2 => n12937, B1 => 
                           REGISTERS_24_12_port, B2 => n12942, ZN => n12638);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n12902, B1 => 
                           REGISTERS_22_12_port, B2 => n12944, ZN => n12637);
   U2553 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n12931, B1 => 
                           REGISTERS_27_12_port, B2 => n12932, ZN => n12636);
   U2554 : NAND4_X1 port map( A1 => n12639, A2 => n12638, A3 => n12637, A4 => 
                           n12636, ZN => n12640);
   U2555 : NOR2_X1 port map( A1 => n12641, A2 => n12640, ZN => n12653);
   U2556 : AOI22_X1 port map( A1 => REGISTERS_2_12_port, A2 => n12954, B1 => 
                           REGISTERS_5_12_port, B2 => n12963, ZN => n12645);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n12967, B1 => 
                           REGISTERS_3_12_port, B2 => n12960, ZN => n12644);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n12851, B1 => 
                           REGISTERS_4_12_port, B2 => n12965, ZN => n12643);
   U2559 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n12962, B1 => 
                           REGISTERS_6_12_port, B2 => n12889, ZN => n12642);
   U2560 : NAND4_X1 port map( A1 => n12645, A2 => n12644, A3 => n12643, A4 => 
                           n12642, ZN => n12651);
   U2561 : AOI22_X1 port map( A1 => REGISTERS_10_12_port, A2 => n12966, B1 => 
                           REGISTERS_11_12_port, B2 => n12914, ZN => n12649);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n12882, B1 => 
                           REGISTERS_13_12_port, B2 => n12951, ZN => n12648);
   U2563 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n12851, B1 => 
                           REGISTERS_9_12_port, B2 => n12952, ZN => n12647);
   U2564 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n12889, B1 => 
                           REGISTERS_8_12_port, B2 => n12962, ZN => n12646);
   U2565 : NAND4_X1 port map( A1 => n12649, A2 => n12648, A3 => n12647, A4 => 
                           n12646, ZN => n12650);
   U2566 : AOI22_X1 port map( A1 => n12813, A2 => n12651, B1 => n12811, B2 => 
                           n12650, ZN => n12652);
   U2567 : OAI21_X1 port map( B1 => n12978, B2 => n12653, A => n12652, ZN => 
                           N397);
   U2568 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n12931, B1 => 
                           REGISTERS_28_11_port, B2 => n12926, ZN => n12657);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n12938, B1 => 
                           REGISTERS_22_11_port, B2 => n12944, ZN => n12656);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n12930, B1 => 
                           REGISTERS_31_11_port, B2 => n12943, ZN => n12655);
   U2571 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n12873, B1 => 
                           REGISTERS_21_11_port, B2 => n12902, ZN => n12654);
   U2572 : NAND4_X1 port map( A1 => n12657, A2 => n12656, A3 => n12655, A4 => 
                           n12654, ZN => n12664);
   U2573 : AOI22_X1 port map( A1 => REGISTERS_18_11_port, A2 => n12937, B1 => 
                           REGISTERS_19_11_port, B2 => n12925, ZN => n12662);
   U2574 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n12658, B1 => 
                           REGISTERS_26_11_port, B2 => n12866, ZN => n12661);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_30_11_port, A2 => n12941, B1 => 
                           REGISTERS_27_11_port, B2 => n12932, ZN => n12660);
   U2576 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n12928, B1 => 
                           REGISTERS_24_11_port, B2 => n12942, ZN => n12659);
   U2577 : NAND4_X1 port map( A1 => n12662, A2 => n12661, A3 => n12660, A4 => 
                           n12659, ZN => n12663);
   U2578 : NOR2_X1 port map( A1 => n12664, A2 => n12663, ZN => n12676);
   U2579 : AOI22_X1 port map( A1 => REGISTERS_2_11_port, A2 => n12881, B1 => 
                           REGISTERS_1_11_port, B2 => n12884, ZN => n12668);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n12965, B1 => 
                           REGISTERS_0_11_port, B2 => n12915, ZN => n12667);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n12851, B1 => 
                           REGISTERS_6_11_port, B2 => n12889, ZN => n12666);
   U2582 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n12963, B1 => 
                           REGISTERS_3_11_port, B2 => n12914, ZN => n12665);
   U2583 : NAND4_X1 port map( A1 => n12668, A2 => n12667, A3 => n12666, A4 => 
                           n12665, ZN => n12674);
   U2584 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n12963, B1 => 
                           REGISTERS_11_11_port, B2 => n12852, ZN => n12672);
   U2585 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n12954, B1 => 
                           REGISTERS_9_11_port, B2 => n12952, ZN => n12671);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n12882, B1 => 
                           REGISTERS_15_11_port, B2 => n12961, ZN => n12670);
   U2587 : AOI22_X1 port map( A1 => REGISTERS_14_11_port, A2 => n12883, B1 => 
                           REGISTERS_8_11_port, B2 => n12962, ZN => n12669);
   U2588 : NAND4_X1 port map( A1 => n12672, A2 => n12671, A3 => n12670, A4 => 
                           n12669, ZN => n12673);
   U2589 : AOI22_X1 port map( A1 => n12813, A2 => n12674, B1 => n12811, B2 => 
                           n12673, ZN => n12675);
   U2590 : OAI21_X1 port map( B1 => n12978, B2 => n12676, A => n12675, ZN => 
                           N396);
   U2591 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n12942, B1 => 
                           REGISTERS_28_10_port, B2 => n12867, ZN => n12682);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n12677, B1 => 
                           REGISTERS_20_10_port, B2 => n12771, ZN => n12681);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_18_10_port, A2 => n12937, B1 => 
                           REGISTERS_31_10_port, B2 => n12943, ZN => n12680);
   U2594 : AOI22_X1 port map( A1 => REGISTERS_26_10_port, A2 => n12866, B1 => 
                           REGISTERS_30_10_port, B2 => n12678, ZN => n12679);
   U2595 : NAND4_X1 port map( A1 => n12682, A2 => n12681, A3 => n12680, A4 => 
                           n12679, ZN => n12688);
   U2596 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n12928, B1 => 
                           REGISTERS_23_10_port, B2 => n12927, ZN => n12686);
   U2597 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n12873, B1 => 
                           REGISTERS_21_10_port, B2 => n12940, ZN => n12685);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n12932, B1 => 
                           REGISTERS_25_10_port, B2 => n12938, ZN => n12684);
   U2599 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n12930, B1 => 
                           REGISTERS_22_10_port, B2 => n12944, ZN => n12683);
   U2600 : NAND4_X1 port map( A1 => n12686, A2 => n12685, A3 => n12684, A4 => 
                           n12683, ZN => n12687);
   U2601 : NOR2_X1 port map( A1 => n12688, A2 => n12687, ZN => n12700);
   U2602 : AOI22_X1 port map( A1 => REGISTERS_2_10_port, A2 => n12966, B1 => 
                           REGISTERS_0_10_port, B2 => n12915, ZN => n12692);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n12851, B1 => 
                           REGISTERS_1_10_port, B2 => n12952, ZN => n12691);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_6_10_port, A2 => n12964, B1 => 
                           REGISTERS_4_10_port, B2 => n12913, ZN => n12690);
   U2605 : AOI22_X1 port map( A1 => REGISTERS_3_10_port, A2 => n12852, B1 => 
                           REGISTERS_5_10_port, B2 => n12805, ZN => n12689);
   U2606 : NAND4_X1 port map( A1 => n12692, A2 => n12691, A3 => n12690, A4 => 
                           n12689, ZN => n12698);
   U2607 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n12965, B1 => 
                           REGISTERS_14_10_port, B2 => n12889, ZN => n12696);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n12960, B1 => 
                           REGISTERS_8_10_port, B2 => n12915, ZN => n12695);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n12967, B1 => 
                           REGISTERS_15_10_port, B2 => n12851, ZN => n12694);
   U2610 : AOI22_X1 port map( A1 => REGISTERS_10_10_port, A2 => n12881, B1 => 
                           REGISTERS_13_10_port, B2 => n12805, ZN => n12693);
   U2611 : NAND4_X1 port map( A1 => n12696, A2 => n12695, A3 => n12694, A4 => 
                           n12693, ZN => n12697);
   U2612 : AOI22_X1 port map( A1 => n12813, A2 => n12698, B1 => n12811, B2 => 
                           n12697, ZN => n12699);
   U2613 : OAI21_X1 port map( B1 => n12978, B2 => n12700, A => n12699, ZN => 
                           N395);
   U2614 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n12926, B1 => 
                           REGISTERS_19_9_port, B2 => n12925, ZN => n12704);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n12927, B1 => 
                           REGISTERS_25_9_port, B2 => n12938, ZN => n12703);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_30_9_port, A2 => n12941, B1 => 
                           REGISTERS_24_9_port, B2 => n12942, ZN => n12702);
   U2617 : AOI22_X1 port map( A1 => REGISTERS_22_9_port, A2 => n12944, B1 => 
                           REGISTERS_18_9_port, B2 => n12937, ZN => n12701);
   U2618 : NAND4_X1 port map( A1 => n12704, A2 => n12703, A3 => n12702, A4 => 
                           n12701, ZN => n12710);
   U2619 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n12931, B1 => 
                           REGISTERS_27_9_port, B2 => n12872, ZN => n12708);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n12902, B1 => 
                           REGISTERS_26_9_port, B2 => n12929, ZN => n12707);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n12873, B1 => 
                           REGISTERS_29_9_port, B2 => n12843, ZN => n12706);
   U2622 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n12943, B1 => 
                           REGISTERS_16_9_port, B2 => n12865, ZN => n12705);
   U2623 : NAND4_X1 port map( A1 => n12708, A2 => n12707, A3 => n12706, A4 => 
                           n12705, ZN => n12709);
   U2624 : NOR2_X1 port map( A1 => n12710, A2 => n12709, ZN => n12722);
   U2625 : AOI22_X1 port map( A1 => REGISTERS_6_9_port, A2 => n12883, B1 => 
                           REGISTERS_7_9_port, B2 => n12961, ZN => n12714);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n12852, B1 => 
                           REGISTERS_1_9_port, B2 => n12884, ZN => n12713);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n12882, B1 => 
                           REGISTERS_2_9_port, B2 => n12881, ZN => n12712);
   U2628 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n12963, B1 => 
                           REGISTERS_0_9_port, B2 => n12955, ZN => n12711);
   U2629 : NAND4_X1 port map( A1 => n12714, A2 => n12713, A3 => n12712, A4 => 
                           n12711, ZN => n12720);
   U2630 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n12915, B1 => 
                           REGISTERS_9_9_port, B2 => n12952, ZN => n12718);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_10_9_port, A2 => n12954, B1 => 
                           REGISTERS_13_9_port, B2 => n12805, ZN => n12717);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n12965, B1 => 
                           REGISTERS_11_9_port, B2 => n12852, ZN => n12716);
   U2633 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n12961, B1 => 
                           REGISTERS_14_9_port, B2 => n12883, ZN => n12715);
   U2634 : NAND4_X1 port map( A1 => n12718, A2 => n12717, A3 => n12716, A4 => 
                           n12715, ZN => n12719);
   U2635 : AOI22_X1 port map( A1 => n12813, A2 => n12720, B1 => n12811, B2 => 
                           n12719, ZN => n12721);
   U2636 : OAI21_X1 port map( B1 => n12924, B2 => n12722, A => n12721, ZN => 
                           N394);
   U2637 : AOI22_X1 port map( A1 => REGISTERS_30_8_port, A2 => n12941, B1 => 
                           REGISTERS_28_8_port, B2 => n12867, ZN => n12726);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n12928, B1 => 
                           REGISTERS_26_8_port, B2 => n12929, ZN => n12725);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n12930, B1 => 
                           REGISTERS_20_8_port, B2 => n12931, ZN => n12724);
   U2640 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n12942, B1 => 
                           REGISTERS_31_8_port, B2 => n12943, ZN => n12723);
   U2641 : NAND4_X1 port map( A1 => n12726, A2 => n12725, A3 => n12724, A4 => 
                           n12723, ZN => n12732);
   U2642 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n12925, B1 => 
                           REGISTERS_21_8_port, B2 => n12940, ZN => n12730);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n12927, B1 => 
                           REGISTERS_25_8_port, B2 => n12938, ZN => n12729);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n12873, B1 => 
                           REGISTERS_22_8_port, B2 => n12944, ZN => n12728);
   U2645 : AOI22_X1 port map( A1 => REGISTERS_18_8_port, A2 => n12937, B1 => 
                           REGISTERS_27_8_port, B2 => n12872, ZN => n12727);
   U2646 : NAND4_X1 port map( A1 => n12730, A2 => n12729, A3 => n12728, A4 => 
                           n12727, ZN => n12731);
   U2647 : NOR2_X1 port map( A1 => n12732, A2 => n12731, ZN => n12744);
   U2648 : AOI22_X1 port map( A1 => REGISTERS_2_8_port, A2 => n12954, B1 => 
                           REGISTERS_3_8_port, B2 => n12960, ZN => n12736);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n12915, B1 => 
                           REGISTERS_4_8_port, B2 => n12913, ZN => n12735);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n12851, B1 => 
                           REGISTERS_1_8_port, B2 => n12884, ZN => n12734);
   U2651 : AOI22_X1 port map( A1 => REGISTERS_6_8_port, A2 => n12964, B1 => 
                           REGISTERS_5_8_port, B2 => n12805, ZN => n12733);
   U2652 : NAND4_X1 port map( A1 => n12736, A2 => n12735, A3 => n12734, A4 => 
                           n12733, ZN => n12742);
   U2653 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n12914, B1 => 
                           REGISTERS_8_8_port, B2 => n12962, ZN => n12740);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_14_8_port, A2 => n12889, B1 => 
                           REGISTERS_12_8_port, B2 => n12965, ZN => n12739);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_10_8_port, A2 => n12881, B1 => 
                           REGISTERS_15_8_port, B2 => n12953, ZN => n12738);
   U2656 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n12967, B1 => 
                           REGISTERS_13_8_port, B2 => n12805, ZN => n12737);
   U2657 : NAND4_X1 port map( A1 => n12740, A2 => n12739, A3 => n12738, A4 => 
                           n12737, ZN => n12741);
   U2658 : AOI22_X1 port map( A1 => n12813, A2 => n12742, B1 => n12811, B2 => 
                           n12741, ZN => n12743);
   U2659 : OAI21_X1 port map( B1 => n12978, B2 => n12744, A => n12743, ZN => 
                           N393);
   U2660 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n12930, B1 => 
                           REGISTERS_28_7_port, B2 => n12867, ZN => n12748);
   U2661 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n12931, B1 => 
                           REGISTERS_18_7_port, B2 => n12874, ZN => n12747);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_31_7_port, A2 => n12943, B1 => 
                           REGISTERS_24_7_port, B2 => n12942, ZN => n12746);
   U2663 : AOI22_X1 port map( A1 => REGISTERS_26_7_port, A2 => n12866, B1 => 
                           REGISTERS_27_7_port, B2 => n12872, ZN => n12745);
   U2664 : NAND4_X1 port map( A1 => n12748, A2 => n12747, A3 => n12746, A4 => 
                           n12745, ZN => n12754);
   U2665 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n12928, B1 => 
                           REGISTERS_19_7_port, B2 => n12925, ZN => n12752);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n12873, B1 => 
                           REGISTERS_25_7_port, B2 => n12938, ZN => n12751);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n12944, B1 => 
                           REGISTERS_21_7_port, B2 => n12940, ZN => n12750);
   U2668 : AOI22_X1 port map( A1 => REGISTERS_30_7_port, A2 => n12941, B1 => 
                           REGISTERS_23_7_port, B2 => n12927, ZN => n12749);
   U2669 : NAND4_X1 port map( A1 => n12752, A2 => n12751, A3 => n12750, A4 => 
                           n12749, ZN => n12753);
   U2670 : NOR2_X1 port map( A1 => n12754, A2 => n12753, ZN => n12766);
   U2671 : AOI22_X1 port map( A1 => REGISTERS_2_7_port, A2 => n12954, B1 => 
                           REGISTERS_6_7_port, B2 => n12964, ZN => n12758);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n12961, B1 => 
                           REGISTERS_5_7_port, B2 => n12805, ZN => n12757);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n12852, B1 => 
                           REGISTERS_0_7_port, B2 => n12915, ZN => n12756);
   U2674 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n12882, B1 => 
                           REGISTERS_1_7_port, B2 => n12952, ZN => n12755);
   U2675 : NAND4_X1 port map( A1 => n12758, A2 => n12757, A3 => n12756, A4 => 
                           n12755, ZN => n12764);
   U2676 : AOI22_X1 port map( A1 => REGISTERS_14_7_port, A2 => n12964, B1 => 
                           REGISTERS_12_7_port, B2 => n12913, ZN => n12762);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_15_7_port, A2 => n12961, B1 => 
                           REGISTERS_11_7_port, B2 => n12960, ZN => n12761);
   U2678 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n12967, B1 => 
                           REGISTERS_13_7_port, B2 => n12951, ZN => n12760);
   U2679 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n12915, B1 => 
                           REGISTERS_10_7_port, B2 => n12966, ZN => n12759);
   U2680 : NAND4_X1 port map( A1 => n12762, A2 => n12761, A3 => n12760, A4 => 
                           n12759, ZN => n12763);
   U2681 : AOI22_X1 port map( A1 => n12813, A2 => n12764, B1 => n12811, B2 => 
                           n12763, ZN => n12765);
   U2682 : OAI21_X1 port map( B1 => n12924, B2 => n12766, A => n12765, ZN => 
                           N392);
   U2683 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n12928, B1 => 
                           REGISTERS_27_6_port, B2 => n12872, ZN => n12770);
   U2684 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n12930, B1 => 
                           REGISTERS_18_6_port, B2 => n12874, ZN => n12769);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_26_6_port, A2 => n12866, B1 => 
                           REGISTERS_23_6_port, B2 => n12927, ZN => n12768);
   U2686 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n12938, B1 => 
                           REGISTERS_24_6_port, B2 => n12942, ZN => n12767);
   U2687 : NAND4_X1 port map( A1 => n12770, A2 => n12769, A3 => n12768, A4 => 
                           n12767, ZN => n12777);
   U2688 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n12902, B1 => 
                           REGISTERS_19_6_port, B2 => n12925, ZN => n12775);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n12771, B1 => 
                           REGISTERS_30_6_port, B2 => n12941, ZN => n12774);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_31_6_port, A2 => n12943, B1 => 
                           REGISTERS_17_6_port, B2 => n12939, ZN => n12773);
   U2691 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n12926, B1 => 
                           REGISTERS_22_6_port, B2 => n12944, ZN => n12772);
   U2692 : NAND4_X1 port map( A1 => n12775, A2 => n12774, A3 => n12773, A4 => 
                           n12772, ZN => n12776);
   U2693 : NOR2_X1 port map( A1 => n12777, A2 => n12776, ZN => n12790);
   U2694 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n12882, B1 => 
                           REGISTERS_0_6_port, B2 => n12955, ZN => n12781);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n12967, B1 => 
                           REGISTERS_7_6_port, B2 => n12851, ZN => n12780);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n12963, B1 => 
                           REGISTERS_3_6_port, B2 => n12914, ZN => n12779);
   U2697 : AOI22_X1 port map( A1 => REGISTERS_6_6_port, A2 => n12889, B1 => 
                           REGISTERS_2_6_port, B2 => n12881, ZN => n12778);
   U2698 : NAND4_X1 port map( A1 => n12781, A2 => n12780, A3 => n12779, A4 => 
                           n12778, ZN => n12787);
   U2699 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n12967, B1 => 
                           REGISTERS_14_6_port, B2 => n12883, ZN => n12785);
   U2700 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n12852, B1 => 
                           REGISTERS_13_6_port, B2 => n12951, ZN => n12784);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_10_6_port, A2 => n12954, B1 => 
                           REGISTERS_8_6_port, B2 => n12962, ZN => n12783);
   U2702 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n12953, B1 => 
                           REGISTERS_12_6_port, B2 => n12913, ZN => n12782);
   U2703 : NAND4_X1 port map( A1 => n12785, A2 => n12784, A3 => n12783, A4 => 
                           n12782, ZN => n12786);
   U2704 : AOI22_X1 port map( A1 => n12788, A2 => n12787, B1 => n12811, B2 => 
                           n12786, ZN => n12789);
   U2705 : OAI21_X1 port map( B1 => n12978, B2 => n12790, A => n12789, ZN => 
                           N391);
   U2706 : AOI22_X1 port map( A1 => REGISTERS_26_5_port, A2 => n12866, B1 => 
                           REGISTERS_16_5_port, B2 => n12865, ZN => n12794);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n12873, B1 => 
                           REGISTERS_31_5_port, B2 => n12943, ZN => n12793);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n12926, B1 => 
                           REGISTERS_19_5_port, B2 => n12925, ZN => n12792);
   U2709 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n12902, B1 => 
                           REGISTERS_20_5_port, B2 => n12931, ZN => n12791);
   U2710 : NAND4_X1 port map( A1 => n12794, A2 => n12793, A3 => n12792, A4 => 
                           n12791, ZN => n12800);
   U2711 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n12938, B1 => 
                           REGISTERS_24_5_port, B2 => n12942, ZN => n12798);
   U2712 : AOI22_X1 port map( A1 => REGISTERS_18_5_port, A2 => n12937, B1 => 
                           REGISTERS_23_5_port, B2 => n12927, ZN => n12797);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_30_5_port, A2 => n12941, B1 => 
                           REGISTERS_29_5_port, B2 => n12843, ZN => n12796);
   U2714 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n12932, B1 => 
                           REGISTERS_22_5_port, B2 => n12944, ZN => n12795);
   U2715 : NAND4_X1 port map( A1 => n12798, A2 => n12797, A3 => n12796, A4 => 
                           n12795, ZN => n12799);
   U2716 : NOR2_X1 port map( A1 => n12800, A2 => n12799, ZN => n12815);
   U2717 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n12962, B1 => 
                           REGISTERS_6_5_port, B2 => n12889, ZN => n12804);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n12953, B1 => 
                           REGISTERS_4_5_port, B2 => n12965, ZN => n12803);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n12963, B1 => 
                           REGISTERS_3_5_port, B2 => n12852, ZN => n12802);
   U2720 : AOI22_X1 port map( A1 => REGISTERS_2_5_port, A2 => n12954, B1 => 
                           REGISTERS_1_5_port, B2 => n12884, ZN => n12801);
   U2721 : NAND4_X1 port map( A1 => n12804, A2 => n12803, A3 => n12802, A4 => 
                           n12801, ZN => n12812);
   U2722 : AOI22_X1 port map( A1 => REGISTERS_14_5_port, A2 => n12964, B1 => 
                           REGISTERS_15_5_port, B2 => n12961, ZN => n12809);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n12955, B1 => 
                           REGISTERS_10_5_port, B2 => n12881, ZN => n12808);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n12967, B1 => 
                           REGISTERS_13_5_port, B2 => n12805, ZN => n12807);
   U2725 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n12965, B1 => 
                           REGISTERS_11_5_port, B2 => n12960, ZN => n12806);
   U2726 : NAND4_X1 port map( A1 => n12809, A2 => n12808, A3 => n12807, A4 => 
                           n12806, ZN => n12810);
   U2727 : AOI22_X1 port map( A1 => n12813, A2 => n12812, B1 => n12811, B2 => 
                           n12810, ZN => n12814);
   U2728 : OAI21_X1 port map( B1 => n12924, B2 => n12815, A => n12814, ZN => 
                           N390);
   U2729 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n12932, B1 => 
                           REGISTERS_28_4_port, B2 => n12867, ZN => n12819);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n12930, B1 => 
                           REGISTERS_16_4_port, B2 => n12865, ZN => n12818);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_26_4_port, A2 => n12866, B1 => 
                           REGISTERS_23_4_port, B2 => n12927, ZN => n12817);
   U2732 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n12902, B1 => 
                           REGISTERS_18_4_port, B2 => n12874, ZN => n12816);
   U2733 : NAND4_X1 port map( A1 => n12819, A2 => n12818, A3 => n12817, A4 => 
                           n12816, ZN => n12825);
   U2734 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n12873, B1 => 
                           REGISTERS_24_4_port, B2 => n12942, ZN => n12823);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_31_4_port, A2 => n12943, B1 => 
                           REGISTERS_30_4_port, B2 => n12941, ZN => n12822);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n12844, B1 => 
                           REGISTERS_20_4_port, B2 => n12931, ZN => n12821);
   U2737 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n12925, B1 => 
                           REGISTERS_25_4_port, B2 => n12938, ZN => n12820);
   U2738 : NAND4_X1 port map( A1 => n12823, A2 => n12822, A3 => n12821, A4 => 
                           n12820, ZN => n12824);
   U2739 : NOR2_X1 port map( A1 => n12825, A2 => n12824, ZN => n12837);
   U2740 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n12914, B1 => 
                           REGISTERS_4_4_port, B2 => n12882, ZN => n12829);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_2_4_port, A2 => n12954, B1 => 
                           REGISTERS_1_4_port, B2 => n12884, ZN => n12828);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n12961, B1 => 
                           REGISTERS_0_4_port, B2 => n12915, ZN => n12827);
   U2743 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n12963, B1 => 
                           REGISTERS_6_4_port, B2 => n12964, ZN => n12826);
   U2744 : NAND4_X1 port map( A1 => n12829, A2 => n12828, A3 => n12827, A4 => 
                           n12826, ZN => n12835);
   U2745 : AOI22_X1 port map( A1 => REGISTERS_10_4_port, A2 => n12954, B1 => 
                           REGISTERS_8_4_port, B2 => n12955, ZN => n12833);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n12963, B1 => 
                           REGISTERS_14_4_port, B2 => n12964, ZN => n12832);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n12967, B1 => 
                           REGISTERS_15_4_port, B2 => n12953, ZN => n12831);
   U2748 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n12960, B1 => 
                           REGISTERS_12_4_port, B2 => n12882, ZN => n12830);
   U2749 : NAND4_X1 port map( A1 => n12833, A2 => n12832, A3 => n12831, A4 => 
                           n12830, ZN => n12834);
   U2750 : AOI22_X1 port map( A1 => n12975, A2 => n12835, B1 => n12973, B2 => 
                           n12834, ZN => n12836);
   U2751 : OAI21_X1 port map( B1 => n12978, B2 => n12837, A => n12836, ZN => 
                           N389);
   U2752 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n12938, B1 => 
                           REGISTERS_23_3_port, B2 => n12927, ZN => n12842);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n12926, B1 => 
                           REGISTERS_16_3_port, B2 => n12865, ZN => n12841);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_31_3_port, A2 => n12838, B1 => 
                           REGISTERS_27_3_port, B2 => n12872, ZN => n12840);
   U2755 : AOI22_X1 port map( A1 => REGISTERS_18_3_port, A2 => n12937, B1 => 
                           REGISTERS_30_3_port, B2 => n12941, ZN => n12839);
   U2756 : NAND4_X1 port map( A1 => n12842, A2 => n12841, A3 => n12840, A4 => 
                           n12839, ZN => n12850);
   U2757 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n12902, B1 => 
                           REGISTERS_29_3_port, B2 => n12843, ZN => n12848);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n12925, B1 => 
                           REGISTERS_20_3_port, B2 => n12931, ZN => n12847);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_22_3_port, A2 => n12844, B1 => 
                           REGISTERS_24_3_port, B2 => n12942, ZN => n12846);
   U2760 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n12873, B1 => 
                           REGISTERS_26_3_port, B2 => n12929, ZN => n12845);
   U2761 : NAND4_X1 port map( A1 => n12848, A2 => n12847, A3 => n12846, A4 => 
                           n12845, ZN => n12849);
   U2762 : NOR2_X1 port map( A1 => n12850, A2 => n12849, ZN => n12864);
   U2763 : AOI22_X1 port map( A1 => REGISTERS_6_3_port, A2 => n12964, B1 => 
                           REGISTERS_0_3_port, B2 => n12955, ZN => n12856);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n12954, B1 => 
                           REGISTERS_5_3_port, B2 => n12951, ZN => n12855);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_7_3_port, A2 => n12851, B1 => 
                           REGISTERS_4_3_port, B2 => n12965, ZN => n12854);
   U2766 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n12967, B1 => 
                           REGISTERS_3_3_port, B2 => n12852, ZN => n12853);
   U2767 : NAND4_X1 port map( A1 => n12856, A2 => n12855, A3 => n12854, A4 => 
                           n12853, ZN => n12862);
   U2768 : AOI22_X1 port map( A1 => REGISTERS_14_3_port, A2 => n12964, B1 => 
                           REGISTERS_8_3_port, B2 => n12962, ZN => n12860);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n12967, B1 => 
                           REGISTERS_11_3_port, B2 => n12960, ZN => n12859);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_15_3_port, A2 => n12953, B1 => 
                           REGISTERS_10_3_port, B2 => n12881, ZN => n12858);
   U2771 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n12963, B1 => 
                           REGISTERS_12_3_port, B2 => n12882, ZN => n12857);
   U2772 : NAND4_X1 port map( A1 => n12860, A2 => n12859, A3 => n12858, A4 => 
                           n12857, ZN => n12861);
   U2773 : AOI22_X1 port map( A1 => n12975, A2 => n12862, B1 => n12973, B2 => 
                           n12861, ZN => n12863);
   U2774 : OAI21_X1 port map( B1 => n12924, B2 => n12864, A => n12863, ZN => 
                           N388);
   U2775 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n12930, B1 => 
                           REGISTERS_30_2_port, B2 => n12941, ZN => n12871);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_26_2_port, A2 => n12866, B1 => 
                           REGISTERS_16_2_port, B2 => n12865, ZN => n12870);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n12927, B1 => 
                           REGISTERS_19_2_port, B2 => n12925, ZN => n12869);
   U2778 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n12943, B1 => 
                           REGISTERS_28_2_port, B2 => n12867, ZN => n12868);
   U2779 : NAND4_X1 port map( A1 => n12871, A2 => n12870, A3 => n12869, A4 => 
                           n12868, ZN => n12880);
   U2780 : AOI22_X1 port map( A1 => REGISTERS_22_2_port, A2 => n12944, B1 => 
                           REGISTERS_25_2_port, B2 => n12938, ZN => n12878);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n12902, B1 => 
                           REGISTERS_27_2_port, B2 => n12872, ZN => n12877);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n12873, B1 => 
                           REGISTERS_20_2_port, B2 => n12931, ZN => n12876);
   U2783 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n12942, B1 => 
                           REGISTERS_18_2_port, B2 => n12874, ZN => n12875);
   U2784 : NAND4_X1 port map( A1 => n12878, A2 => n12877, A3 => n12876, A4 => 
                           n12875, ZN => n12879);
   U2785 : NOR2_X1 port map( A1 => n12880, A2 => n12879, ZN => n12897);
   U2786 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n12955, B1 => 
                           REGISTERS_2_2_port, B2 => n12881, ZN => n12888);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n12882, B1 => 
                           REGISTERS_3_2_port, B2 => n12914, ZN => n12887);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n12961, B1 => 
                           REGISTERS_6_2_port, B2 => n12883, ZN => n12886);
   U2789 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n12963, B1 => 
                           REGISTERS_1_2_port, B2 => n12884, ZN => n12885);
   U2790 : NAND4_X1 port map( A1 => n12888, A2 => n12887, A3 => n12886, A4 => 
                           n12885, ZN => n12895);
   U2791 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n12963, B1 => 
                           REGISTERS_15_2_port, B2 => n12953, ZN => n12893);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n12955, B1 => 
                           REGISTERS_11_2_port, B2 => n12914, ZN => n12892);
   U2793 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n12967, B1 => 
                           REGISTERS_12_2_port, B2 => n12965, ZN => n12891);
   U2794 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n12954, B1 => 
                           REGISTERS_14_2_port, B2 => n12889, ZN => n12890);
   U2795 : NAND4_X1 port map( A1 => n12893, A2 => n12892, A3 => n12891, A4 => 
                           n12890, ZN => n12894);
   U2796 : AOI22_X1 port map( A1 => n12975, A2 => n12895, B1 => n12973, B2 => 
                           n12894, ZN => n12896);
   U2797 : OAI21_X1 port map( B1 => n12978, B2 => n12897, A => n12896, ZN => 
                           N387);
   U2798 : AOI22_X1 port map( A1 => REGISTERS_27_1_port, A2 => n12932, B1 => 
                           REGISTERS_25_1_port, B2 => n12938, ZN => n12901);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n12928, B1 => 
                           REGISTERS_31_1_port, B2 => n12943, ZN => n12900);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n12930, B1 => 
                           REGISTERS_22_1_port, B2 => n12944, ZN => n12899);
   U2801 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n12931, B1 => 
                           REGISTERS_30_1_port, B2 => n12941, ZN => n12898);
   U2802 : NAND4_X1 port map( A1 => n12901, A2 => n12900, A3 => n12899, A4 => 
                           n12898, ZN => n12908);
   U2803 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n12925, B1 => 
                           REGISTERS_17_1_port, B2 => n12939, ZN => n12906);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n12926, B1 => 
                           REGISTERS_24_1_port, B2 => n12942, ZN => n12905);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n12937, B1 => 
                           REGISTERS_26_1_port, B2 => n12929, ZN => n12904);
   U2806 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n12902, B1 => 
                           REGISTERS_23_1_port, B2 => n12927, ZN => n12903);
   U2807 : NAND4_X1 port map( A1 => n12906, A2 => n12905, A3 => n12904, A4 => 
                           n12903, ZN => n12907);
   U2808 : NOR2_X1 port map( A1 => n12908, A2 => n12907, ZN => n12923);
   U2809 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n12964, B1 => 
                           REGISTERS_1_1_port, B2 => n12952, ZN => n12912);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_3_1_port, A2 => n12914, B1 => 
                           REGISTERS_0_1_port, B2 => n12915, ZN => n12911);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n12953, B1 => 
                           REGISTERS_4_1_port, B2 => n12913, ZN => n12910);
   U2812 : AOI22_X1 port map( A1 => REGISTERS_2_1_port, A2 => n12954, B1 => 
                           REGISTERS_5_1_port, B2 => n12951, ZN => n12909);
   U2813 : NAND4_X1 port map( A1 => n12912, A2 => n12911, A3 => n12910, A4 => 
                           n12909, ZN => n12921);
   U2814 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n12914, B1 => 
                           REGISTERS_12_1_port, B2 => n12913, ZN => n12919);
   U2815 : AOI22_X1 port map( A1 => REGISTERS_10_1_port, A2 => n12954, B1 => 
                           REGISTERS_13_1_port, B2 => n12951, ZN => n12918);
   U2816 : AOI22_X1 port map( A1 => REGISTERS_14_1_port, A2 => n12964, B1 => 
                           REGISTERS_9_1_port, B2 => n12952, ZN => n12917);
   U2817 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n12953, B1 => 
                           REGISTERS_8_1_port, B2 => n12915, ZN => n12916);
   U2818 : NAND4_X1 port map( A1 => n12919, A2 => n12918, A3 => n12917, A4 => 
                           n12916, ZN => n12920);
   U2819 : AOI22_X1 port map( A1 => n12975, A2 => n12921, B1 => n12973, B2 => 
                           n12920, ZN => n12922);
   U2820 : OAI21_X1 port map( B1 => n12924, B2 => n12923, A => n12922, ZN => 
                           N386);
   U2821 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n12926, B1 => 
                           REGISTERS_19_0_port, B2 => n12925, ZN => n12936);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n12928, B1 => 
                           REGISTERS_23_0_port, B2 => n12927, ZN => n12935);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n12930, B1 => 
                           REGISTERS_26_0_port, B2 => n12929, ZN => n12934);
   U2824 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n12932, B1 => 
                           REGISTERS_20_0_port, B2 => n12931, ZN => n12933);
   U2825 : NAND4_X1 port map( A1 => n12936, A2 => n12935, A3 => n12934, A4 => 
                           n12933, ZN => n12950);
   U2826 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n12938, B1 => 
                           REGISTERS_18_0_port, B2 => n12937, ZN => n12948);
   U2827 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n12940, B1 => 
                           REGISTERS_17_0_port, B2 => n12939, ZN => n12947);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n12942, B1 => 
                           REGISTERS_30_0_port, B2 => n12941, ZN => n12946);
   U2829 : AOI22_X1 port map( A1 => REGISTERS_22_0_port, A2 => n12944, B1 => 
                           REGISTERS_31_0_port, B2 => n12943, ZN => n12945);
   U2830 : NAND4_X1 port map( A1 => n12948, A2 => n12947, A3 => n12946, A4 => 
                           n12945, ZN => n12949);
   U2831 : NOR2_X1 port map( A1 => n12950, A2 => n12949, ZN => n12977);
   U2832 : AOI22_X1 port map( A1 => REGISTERS_6_0_port, A2 => n12964, B1 => 
                           REGISTERS_5_0_port, B2 => n12951, ZN => n12959);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n12953, B1 => 
                           REGISTERS_1_0_port, B2 => n12952, ZN => n12958);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n12954, B1 => 
                           REGISTERS_3_0_port, B2 => n12960, ZN => n12957);
   U2835 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n12955, B1 => 
                           REGISTERS_4_0_port, B2 => n12965, ZN => n12956);
   U2836 : NAND4_X1 port map( A1 => n12959, A2 => n12958, A3 => n12957, A4 => 
                           n12956, ZN => n12974);
   U2837 : AOI22_X1 port map( A1 => REGISTERS_15_0_port, A2 => n12961, B1 => 
                           REGISTERS_11_0_port, B2 => n12960, ZN => n12971);
   U2838 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n12963, B1 => 
                           REGISTERS_8_0_port, B2 => n12962, ZN => n12970);
   U2839 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n12965, B1 => 
                           REGISTERS_14_0_port, B2 => n12964, ZN => n12969);
   U2840 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n12967, B1 => 
                           REGISTERS_10_0_port, B2 => n12966, ZN => n12968);
   U2841 : NAND4_X1 port map( A1 => n12971, A2 => n12970, A3 => n12969, A4 => 
                           n12968, ZN => n12972);
   U2842 : AOI22_X1 port map( A1 => n12975, A2 => n12974, B1 => n12973, B2 => 
                           n12972, ZN => n12976);
   U2843 : OAI21_X1 port map( B1 => n12978, B2 => n12977, A => n12976, ZN => 
                           N385);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ENABLE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_28_port, 
      curr_instruction_to_cu_i_27_port, curr_instruction_to_cu_i_26_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_5_port, curr_instruction_to_cu_i_4_port, 
      curr_instruction_to_cu_i_3_port, curr_instruction_to_cu_i_2_port, 
      curr_instruction_to_cu_i_1_port, curr_instruction_to_cu_i_0_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n131, cu_i_n127, 
      cu_i_n126, cu_i_n125, cu_i_n124, cu_i_n123, cu_i_n210, cu_i_n209, 
      cu_i_n145, cu_i_n26, cu_i_n25, cu_i_n23, cu_i_cw1_i_4_port, 
      cu_i_cw1_i_7_port, cu_i_cw1_i_8_port, cu_i_cw3_6_port, cu_i_cw2_5_port, 
      cu_i_cw2_6_port, cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_0_port, 
      cu_i_cw1_1_port, cu_i_cw1_2_port, cu_i_cw1_3_port, cu_i_cw1_4_port, 
      cu_i_cw1_5_port, cu_i_cw1_6_port, cu_i_cw1_7_port, cu_i_cw1_8_port, 
      cu_i_cw1_10_port, cu_i_cw1_11_port, cu_i_cw1_12_port, cu_i_N279, 
      cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, 
      cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, 
      cu_i_cmd_word_4_port, cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, 
      cu_i_cmd_word_8_port, cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n78, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_n12, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n309, n311, n691, n697, n699,
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n737, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n756, 
      n758, n759, n760, n761, n762, n763, n764, n1152, n2319, n2704, n2705, 
      n2706, n2707, n2708, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, 
      DRAM_ENABLE_port, n3109, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => n3088, QN => cu_i_n125);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => n_1413, QN => cu_i_n123);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n12, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n43, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1414, mul_exeception => 
                           n_1415, FUNC(0) => n2704, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1416, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n3107, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n3107, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n3107, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n3107, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n309, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n3107, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n3107, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n3107, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n309, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n3107, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n3107, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n3107, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n3107, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n309, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n3107, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n3107, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n3107, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n309, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n3107, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n3107, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n309, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n3107, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n309, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n309, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n309, Z =>
                           DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n309, Z =>
                           DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n3107, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n3107, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n3107, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n3107, Z 
                           => DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n3109, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n3109, Z =>
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n3109, Z =>
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n3109, Z =>
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n3109, Z =>
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n3109, Z =>
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n3109, Z =>
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n3109, Z =>
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n3109, Z =>
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n3109, Z =>
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n3109, Z =>
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n3109, Z =>
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => n3109, Z =>
                           DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => n3109, Z =>
                           DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => n3109, Z =>
                           DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => n3109, Z =>
                           DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => n3109, Z =>
                           DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1417);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n3105, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n3106, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n3105, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n3106, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n3105, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n3106, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n3106, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n3104, D => datapath_i_n18, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n3104, D => datapath_i_n17, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n3104, D => datapath_i_n16, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n3104, D => datapath_i_n15, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n3104, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n3104, D => 
                           curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n3104, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n3104, D => datapath_i_n12, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n3104, D => datapath_i_n11, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n3104, D => datapath_i_n10, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n3104, D => datapath_i_n9, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n2712, CK => CLK, RN => RST
                           , Q => cu_i_cw3_6_port, QN => n_1418);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n131, CK => CLK, RN =>
                           RST, Q => n_1419, QN => n699);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1420);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1421);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1422);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n126, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n3103);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => n_1423, QN => n756);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n3106, CK => CLK, RN => RST
                           , Q => n_1424, QN => n2319);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1425)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1426)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1427)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1428);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1429);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n311, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1430);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1431);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => n1152, CK => CLK, RN => RST,
                           Q => cu_i_cw1_4_port, QN => n_1432);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1433);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1434);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1435);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1436);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1437);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1438);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1439);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1440);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1441);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1442);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1443);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1444);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1445);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1446);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1447);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1448);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1449);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1450);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1451);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1452);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1453);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1454);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1455);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1456);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1457);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1458);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1459);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1460);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1461);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1462);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1463);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1464);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1465);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1466);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1467);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1468)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1469)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1470)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1471)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1472)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1473)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1474)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1475)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1476)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1477)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1478)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1479)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1480)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1481)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1482)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1483)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1484)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1485)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1486)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1487)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1488)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1489)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1490);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1491);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1492);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1493);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1494);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1495);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1496);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1497);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1498);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1499);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1500);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1501);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1502);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1503);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1504);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1505);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1506);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1507);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1508);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1509);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1510);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1511);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1512);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1513);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1514);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1515);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1516);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1517);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1518);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1519);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1520);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1521);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1522);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1523);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1524);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1525);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1526);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1527);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1528);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1529);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1530);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1531);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1532);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1533);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1534);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1535);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1536);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1537);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1538);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1539);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1540);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1541);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1542);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1543);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1544);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1545);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1546);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1547);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1548);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1549);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1550);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1551);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1552);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1553);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1554);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1555);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1556);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1557);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1558);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1559);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1560);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1561);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1562);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1563);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1564, QN => n703);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1565, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1566, QN => n726);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1567, QN => n725);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1568, QN => n724);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1569, QN => n691);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1570, QN => n723);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1571, QN => n722);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1572, QN => n721);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1573, QN => n720);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1574, QN => n719);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1575, QN => n718);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1576, QN => n717);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1577, QN => n716);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1578, QN => n715);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1579, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1580, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1581, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1582, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1583, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1584, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1585, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1586, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1587, QN => n706);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1588, QN => n705);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1589, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1590, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1591, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1592, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1593, QN => n728);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1594, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1595, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1596);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1597);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1598);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1599);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1600);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1601);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1602);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1603);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1604);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1605);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1606);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1607);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1608);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1609);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1610);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1611);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1612);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1613);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1614);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1615);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1616);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1617);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1618);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1619);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1620);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1621);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1622);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1623);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1624);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1625);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1626);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1627);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n3104, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1628);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1629);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1630);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1631);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1632);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1633);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1634);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1635);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1636);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1637);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1638);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1639);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1640);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1641);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1642);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1643);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1644);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1645);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1646);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1647);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1648);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1649);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1650);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1651);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1652);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1653);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1654);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n764);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n763);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n762);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n761);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n760);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n759);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n758);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1655);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1656);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1657);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1658);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1659);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1660);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1661);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1662);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1663);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1664);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1665);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1666);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1667);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1668);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1669);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1670);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1671);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1672);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1673);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1674);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1675);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1676);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1677);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1678);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1679);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1680);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1681);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1682);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1683);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1684);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1685);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1686);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1687);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1688);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1689);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1690);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1691);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1692);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1693);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1694);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1695);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1696);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1697);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1698);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1699);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1700);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1701);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1702);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1703);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1704);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1705);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1706);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1707);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1708);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1709);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1710);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1711);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1712);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1713);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1714);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1715);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1716);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1717);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1718);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1719);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1720);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1721);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => n2708, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1722);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => n2707, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1723);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1724);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => n2706, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1725);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n2705, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1726);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n3101);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n3089);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => n3100, QN => n737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n3085);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n3091);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n3086);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1727);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1728);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1729);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1730);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1731);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1732);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1733);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n697);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1734);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1735);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1736);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1738);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1741);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1742);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1743);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1744);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n_1745);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n3090);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n3098);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n3094);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n3097);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n_1746);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1747
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1748
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1749
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1750
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1751
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1752
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1753
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1754
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1755
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1756
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1757
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1758
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1759
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1760
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1761
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1762
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1763
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1764
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1765
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1766
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1767
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1768
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1769)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1770)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1771)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1772)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1773)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1774)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1775)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1776)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1777)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1778)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1779);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_30_port, QN => 
                           n_1780);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n753);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_28_port, QN => 
                           n_1781);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n751);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_26_port, QN => 
                           n_1782);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n750);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_24_port, QN => 
                           n_1783);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n749);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_22_port, QN => 
                           n_1784);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n748);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_20_port, QN => 
                           n_1785);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n747);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_18_port, QN => 
                           n_1786);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n746);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_16_port, QN => 
                           n_1787);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n745);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_14_port, QN => 
                           n_1788);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n752);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_12_port, QN => 
                           n_1789);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n744);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_10_port, QN => 
                           n_1790);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n743
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_8_port, QN => 
                           n_1791);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n742
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_6_port, QN => 
                           n_1792);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n741
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_1793);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_1794);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_1795);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1796);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1797);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => n3087, QN => n3092);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1798);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => n3095, QN => cu_i_n26);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => n3102, QN => cu_i_n25);
   U2604 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(0), ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   U2605 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(10), ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U2606 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(11), ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U2607 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(12), ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U2608 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(13), ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U2609 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(14), ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U2610 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(15), ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U2611 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U2612 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U2613 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U2614 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U2615 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U2616 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U2617 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(21), ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U2618 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(22), ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U2619 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(23), ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U2620 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(24), ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U2621 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(25), ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U2622 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(26), ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U2623 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(27), ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U2624 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(28), ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U2625 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(29), ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U2626 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U2627 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(30), ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U2628 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(31), ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U2629 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U2630 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U2631 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U2632 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U2633 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U2634 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(8), ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U2635 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => n3096, QN => cu_i_n124);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => n3099, QN => cu_i_n23);
   cu_i_stall_reg : DFFR_X2 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n704, QN => n3093);
   U2636 : NAND2_X1 port map( A1 => n2742, A2 => n3096, ZN => n2843);
   U2637 : AOI21_X1 port map( B1 => n2975, B2 => n2974, A => cu_i_cw3_6_port, 
                           ZN => n2976);
   U2638 : OAI21_X1 port map( B1 => n2843, B2 => n2844, A => n699, ZN => 
                           write_rf_i);
   U2639 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_0_port, B1
                           => cu_i_cw1_0_port, B2 => n3093, ZN => n2799);
   U2640 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_2_port, B1
                           => cu_i_cw1_2_port, B2 => n3093, ZN => n2807);
   U2641 : NAND2_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, ZN => n2742);
   U2642 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U2643 : AOI211_X1 port map( C1 => n2792, C2 => n2851, A => 
                           cu_i_cmd_word_4_port, B => cu_i_cmd_word_7_port, ZN 
                           => n2794);
   U2644 : NOR2_X1 port map( A1 => cu_i_n123, A2 => n3099, ZN => n2792);
   U2645 : CLKBUF_X1 port map( A => n3084, Z => n3073);
   U2646 : CLKBUF_X1 port map( A => n2920, Z => n2969);
   U2647 : AOI21_X1 port map( B1 => n2785, B2 => n2796, A => n2849, ZN => n2972
                           );
   U2648 : NOR4_X1 port map( A1 => n2824, A2 => n2809, A3 => n3094, A4 => n3090
                           , ZN => n2796);
   U2649 : OR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n3091
                           , A3 => n3017, ZN => n3015);
   U2650 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           curr_instruction_to_cu_i_30_port, A3 => n2713, ZN =>
                           cu_i_cmd_word_4_port);
   U2651 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           curr_instruction_to_cu_i_31_port, A3 => n2792, A4 =>
                           curr_instruction_to_cu_i_26_port, ZN => n2713);
   U2652 : OAI22_X1 port map( A1 => n3093, A2 => cu_i_cmd_word_4_port, B1 => 
                           cu_i_cw2_8_port, B2 => n704, ZN => n309);
   U2653 : INV_X1 port map( A => n309, ZN => DRAM_ENABLE_port);
   U2654 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n3107);
   U2655 : INV_X1 port map( A => cu_i_cmd_word_4_port, ZN => n2970);
   U2656 : NOR2_X1 port map( A1 => n3100, A2 => n2970, ZN => 
                           cu_i_cmd_word_3_port);
   U2657 : OAI22_X1 port map( A1 => n3093, A2 => cu_i_cmd_word_3_port, B1 => 
                           cu_i_cw2_7_port, B2 => n704, ZN => n2797);
   U2658 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n2797, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U2659 : CLKBUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n3109);
   U2660 : NAND2_X2 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n3092, ZN => n2963);
   U2661 : INV_X1 port map( A => n3092, ZN => n2961);
   U2662 : NOR2_X1 port map( A1 => n3087, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n2960);
   U2663 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_29_port, ZN => 
                           n2714);
   U2664 : OAI21_X1 port map( B1 => n726, B2 => n2963, A => n2714, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U2665 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_27_port, ZN => 
                           n2715);
   U2666 : OAI21_X1 port map( B1 => n724, B2 => n2963, A => n2715, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U2667 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_25_port, ZN => 
                           n2716);
   U2668 : OAI21_X1 port map( B1 => n723, B2 => n2963, A => n2716, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U2669 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_23_port, ZN => 
                           n2717);
   U2670 : OAI21_X1 port map( B1 => n721, B2 => n2963, A => n2717, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U2671 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_21_port, ZN => 
                           n2718);
   U2672 : OAI21_X1 port map( B1 => n719, B2 => n2963, A => n2718, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U2673 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_19_port, ZN => 
                           n2719);
   U2674 : OAI21_X1 port map( B1 => n717, B2 => n2963, A => n2719, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U2675 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_17_port, ZN => 
                           n2720);
   U2676 : OAI21_X1 port map( B1 => n715, B2 => n2963, A => n2720, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U2677 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_15_port, ZN => 
                           n2721);
   U2678 : OAI21_X1 port map( B1 => n713, B2 => n2963, A => n2721, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U2679 : CLKBUF_X1 port map( A => n2960, Z => n2954);
   U2680 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_13_port, ZN => 
                           n2722);
   U2681 : OAI21_X1 port map( B1 => n711, B2 => n2963, A => n2722, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U2682 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_11_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_11_port, ZN => 
                           n2723);
   U2683 : OAI21_X1 port map( B1 => n709, B2 => n2963, A => n2723, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U2684 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_9_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_9_port, ZN => 
                           n2724);
   U2685 : OAI21_X1 port map( B1 => n707, B2 => n2963, A => n2724, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U2686 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_7_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_7_port, ZN => 
                           n2725);
   U2687 : OAI21_X1 port map( B1 => n705, B2 => n2963, A => n2725, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U2688 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_5_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_5_port, ZN => 
                           n2726);
   U2689 : OAI21_X1 port map( B1 => n731, B2 => n2963, A => n2726, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U2690 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_4_port, ZN => 
                           n2727);
   U2691 : OAI21_X1 port map( B1 => n730, B2 => n2963, A => n2727, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U2692 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_2_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_2_port, ZN => 
                           n2728);
   U2693 : OAI21_X1 port map( B1 => n728, B2 => n2963, A => n2728, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U2694 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_3_port, ZN => 
                           n2729);
   U2695 : OAI21_X1 port map( B1 => n729, B2 => n2963, A => n2729, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U2696 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_6_port, ZN => 
                           n2730);
   U2697 : OAI21_X1 port map( B1 => n732, B2 => n2963, A => n2730, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U2698 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_8_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_8_port, ZN => 
                           n2731);
   U2699 : OAI21_X1 port map( B1 => n706, B2 => n2963, A => n2731, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U2700 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_10_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_10_port, ZN => 
                           n2732);
   U2701 : OAI21_X1 port map( B1 => n708, B2 => n2963, A => n2732, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U2702 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_12_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_12_port, ZN => 
                           n2733);
   U2703 : OAI21_X1 port map( B1 => n710, B2 => n2963, A => n2733, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U2704 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_14_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_14_port, ZN => 
                           n2734);
   U2705 : OAI21_X1 port map( B1 => n712, B2 => n2963, A => n2734, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U2706 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_16_port, B1 => n2960, B2
                           => datapath_i_new_pc_value_decode_16_port, ZN => 
                           n2735);
   U2707 : OAI21_X1 port map( B1 => n714, B2 => n2963, A => n2735, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U2708 : AOI22_X1 port map( A1 => n3087, A2 => 
                           datapath_i_alu_output_val_i_18_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_18_port, ZN => 
                           n2736);
   U2709 : OAI21_X1 port map( B1 => n716, B2 => n2963, A => n2736, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U2710 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_20_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_20_port, ZN => 
                           n2737);
   U2711 : OAI21_X1 port map( B1 => n718, B2 => n2963, A => n2737, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U2712 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_22_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_22_port, ZN => 
                           n2738);
   U2713 : OAI21_X1 port map( B1 => n720, B2 => n2963, A => n2738, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U2714 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_24_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_24_port, ZN => 
                           n2739);
   U2715 : OAI21_X1 port map( B1 => n722, B2 => n2963, A => n2739, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U2716 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_26_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_26_port, ZN => 
                           n2740);
   U2717 : OAI21_X1 port map( B1 => n691, B2 => n2963, A => n2740, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U2718 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_28_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_28_port, ZN => 
                           n2741);
   U2719 : OAI21_X1 port map( B1 => n725, B2 => n2963, A => n2741, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U2720 : NAND4_X1 port map( A1 => n737, A2 => n2792, A3 => n3101, A4 => n3089
                           , ZN => n3017);
   U2721 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n3091, ZN => n2833);
   U2722 : OAI21_X1 port map( B1 => n3017, B2 => n2833, A => n3015, ZN => n1152
                           );
   U2723 : NAND4_X1 port map( A1 => cu_i_n26, A2 => cu_i_n25, A3 => n3088, A4 
                           => n3096, ZN => cu_i_n145);
   U2724 : NAND2_X1 port map( A1 => cu_i_n145, A2 => n2843, ZN => n2785);
   U2725 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_5_port, A2 => 
                           curr_instruction_to_cu_i_1_port, ZN => n2824);
   U2726 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_0_port, ZN => n2809);
   U2727 : NAND3_X1 port map( A1 => n737, A2 => n3101, A3 => n3086, ZN => n2784
                           );
   U2728 : NOR4_X2 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           curr_instruction_to_cu_i_28_port, A3 => 
                           curr_instruction_to_cu_i_30_port, A4 => n2784, ZN =>
                           n2856);
   U2729 : NAND2_X1 port map( A1 => n2796, A2 => n2856, ZN => n2816);
   U2730 : OAI21_X1 port map( B1 => n2785, B2 => n2816, A => n2792, ZN => n2743
                           );
   U2731 : NAND2_X1 port map( A1 => cu_i_n123, A2 => n3099, ZN => n2860);
   U2732 : AOI21_X1 port map( B1 => n2743, B2 => n2860, A => n704, ZN => 
                           IRAM_ENABLE_port);
   U2733 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, 
                           ZN => n2744);
   U2734 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, 
                           ZN => n2747);
   U2735 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, 
                           ZN => n2750);
   U2736 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, 
                           ZN => n2753);
   U2737 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, 
                           ZN => n2756);
   U2738 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, 
                           ZN => n2759);
   U2739 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, 
                           ZN => n2762);
   U2740 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, 
                           ZN => n2765);
   U2741 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, 
                           ZN => n2768);
   U2742 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, 
                           ZN => n2771);
   U2743 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN
                           => n2774);
   U2744 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN
                           => n2777);
   U2745 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN
                           => n2780);
   U2746 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_3_port, ZN =>
                           n2875);
   U2747 : NOR2_X1 port map( A1 => n2780, A2 => n2875, ZN => n2882);
   U2748 : NAND2_X1 port map( A1 => n2882, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n2881);
   U2749 : NOR2_X1 port map( A1 => n2777, A2 => n2881, ZN => n2888);
   U2750 : NAND2_X1 port map( A1 => n2888, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n2887);
   U2751 : NOR2_X1 port map( A1 => n2774, A2 => n2887, ZN => n2894);
   U2752 : NAND2_X1 port map( A1 => n2894, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n2893);
   U2753 : NOR2_X1 port map( A1 => n2771, A2 => n2893, ZN => n2900);
   U2754 : NAND2_X1 port map( A1 => n2900, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n2899);
   U2755 : NOR2_X1 port map( A1 => n2768, A2 => n2899, ZN => n2906);
   U2756 : NAND2_X1 port map( A1 => n2906, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n2905);
   U2757 : NOR2_X1 port map( A1 => n2765, A2 => n2905, ZN => n2912);
   U2758 : NAND2_X1 port map( A1 => n2912, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n2911);
   U2759 : NOR2_X1 port map( A1 => n2762, A2 => n2911, ZN => n2918);
   U2760 : NAND2_X1 port map( A1 => n2918, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n2917);
   U2761 : NOR2_X1 port map( A1 => n2759, A2 => n2917, ZN => n2925);
   U2762 : NAND2_X1 port map( A1 => n2925, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n2924);
   U2763 : NOR2_X1 port map( A1 => n2756, A2 => n2924, ZN => n2931);
   U2764 : NAND2_X1 port map( A1 => n2931, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n2930);
   U2765 : NOR2_X1 port map( A1 => n2753, A2 => n2930, ZN => n2937);
   U2766 : NAND2_X1 port map( A1 => n2937, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n2936);
   U2767 : NOR2_X1 port map( A1 => n2750, A2 => n2936, ZN => n2943);
   U2768 : NAND2_X1 port map( A1 => n2943, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n2942);
   U2769 : NOR2_X1 port map( A1 => n2747, A2 => n2942, ZN => n2949);
   U2770 : NAND2_X1 port map( A1 => n2949, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n2948);
   U2771 : INV_X1 port map( A => n1152, ZN => n2861);
   U2772 : OAI221_X1 port map( B1 => n3093, B2 => n2861, C1 => n704, C2 => n756
                           , A => n3092, ZN => n2872);
   U2773 : INV_X1 port map( A => n2872, ZN => n2920);
   U2774 : NOR2_X1 port map( A1 => n2744, A2 => n2948, ZN => n2956);
   U2775 : AOI211_X1 port map( C1 => n2744, C2 => n2948, A => n2920, B => n2956
                           , ZN => n2746);
   U2776 : NAND2_X1 port map( A1 => IRAM_ENABLE_port, A2 => IRAM_ADDRESS_2_port
                           , ZN => n2869);
   U2777 : INV_X1 port map( A => n2869, ZN => n2871);
   U2778 : AND2_X1 port map( A1 => n2871, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n2878);
   U2779 : NAND2_X1 port map( A1 => n2878, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n2877);
   U2780 : NOR2_X1 port map( A1 => n741, A2 => n2877, ZN => n2884);
   U2781 : NAND2_X1 port map( A1 => n2884, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n2883);
   U2782 : NOR2_X1 port map( A1 => n742, A2 => n2883, ZN => n2890);
   U2783 : NAND2_X1 port map( A1 => n2890, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n2889);
   U2784 : NOR2_X1 port map( A1 => n743, A2 => n2889, ZN => n2896);
   U2785 : NAND2_X1 port map( A1 => n2896, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n2895);
   U2786 : NOR2_X1 port map( A1 => n744, A2 => n2895, ZN => n2902);
   U2787 : NAND2_X1 port map( A1 => n2902, A2 => IRAM_ADDRESS_12_port, ZN => 
                           n2901);
   U2788 : NOR2_X1 port map( A1 => n752, A2 => n2901, ZN => n2908);
   U2789 : NAND2_X1 port map( A1 => n2908, A2 => IRAM_ADDRESS_14_port, ZN => 
                           n2907);
   U2790 : NOR2_X1 port map( A1 => n745, A2 => n2907, ZN => n2914);
   U2791 : NAND2_X1 port map( A1 => n2914, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n2913);
   U2792 : NOR2_X1 port map( A1 => n746, A2 => n2913, ZN => n2921);
   U2793 : NAND2_X1 port map( A1 => n2921, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n2919);
   U2794 : NOR2_X1 port map( A1 => n747, A2 => n2919, ZN => n2927);
   U2795 : NAND2_X1 port map( A1 => n2927, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n2926);
   U2796 : NOR2_X1 port map( A1 => n748, A2 => n2926, ZN => n2933);
   U2797 : NAND2_X1 port map( A1 => n2933, A2 => IRAM_ADDRESS_22_port, ZN => 
                           n2932);
   U2798 : NOR2_X1 port map( A1 => n749, A2 => n2932, ZN => n2939);
   U2799 : NAND2_X1 port map( A1 => n2939, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n2938);
   U2800 : NOR2_X1 port map( A1 => n750, A2 => n2938, ZN => n2945);
   U2801 : NAND2_X1 port map( A1 => n2945, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n2944);
   U2802 : NOR2_X1 port map( A1 => n751, A2 => n2944, ZN => n2951);
   U2803 : NAND2_X1 port map( A1 => n2951, A2 => IRAM_ADDRESS_28_port, ZN => 
                           n2950);
   U2804 : NOR2_X1 port map( A1 => n753, A2 => n2950, ZN => n2957);
   U2805 : AOI211_X1 port map( C1 => n753, C2 => n2950, A => n2957, B => n2872,
                           ZN => n2745);
   U2806 : OR2_X1 port map( A1 => n2746, A2 => n2745, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U2807 : AOI211_X1 port map( C1 => n2747, C2 => n2942, A => n2969, B => n2949
                           , ZN => n2749);
   U2808 : AOI211_X1 port map( C1 => n751, C2 => n2944, A => n2951, B => n2872,
                           ZN => n2748);
   U2809 : OR2_X1 port map( A1 => n2749, A2 => n2748, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U2810 : AOI211_X1 port map( C1 => n2750, C2 => n2936, A => n2920, B => n2943
                           , ZN => n2752);
   U2811 : INV_X1 port map( A => n2969, ZN => n2966);
   U2812 : AOI211_X1 port map( C1 => n750, C2 => n2938, A => n2945, B => n2966,
                           ZN => n2751);
   U2813 : OR2_X1 port map( A1 => n2752, A2 => n2751, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U2814 : AOI211_X1 port map( C1 => n2753, C2 => n2930, A => n2920, B => n2937
                           , ZN => n2755);
   U2815 : AOI211_X1 port map( C1 => n749, C2 => n2932, A => n2939, B => n2966,
                           ZN => n2754);
   U2816 : OR2_X1 port map( A1 => n2755, A2 => n2754, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U2817 : AOI211_X1 port map( C1 => n2756, C2 => n2924, A => n2920, B => n2931
                           , ZN => n2758);
   U2818 : AOI211_X1 port map( C1 => n748, C2 => n2926, A => n2933, B => n2966,
                           ZN => n2757);
   U2819 : OR2_X1 port map( A1 => n2758, A2 => n2757, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U2820 : AOI211_X1 port map( C1 => n2759, C2 => n2917, A => n2920, B => n2925
                           , ZN => n2761);
   U2821 : AOI211_X1 port map( C1 => n747, C2 => n2919, A => n2927, B => n2966,
                           ZN => n2760);
   U2822 : OR2_X1 port map( A1 => n2761, A2 => n2760, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U2823 : AOI211_X1 port map( C1 => n2762, C2 => n2911, A => n2920, B => n2918
                           , ZN => n2764);
   U2824 : AOI211_X1 port map( C1 => n746, C2 => n2913, A => n2921, B => n2872,
                           ZN => n2763);
   U2825 : OR2_X1 port map( A1 => n2764, A2 => n2763, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U2826 : AOI211_X1 port map( C1 => n2765, C2 => n2905, A => n2969, B => n2912
                           , ZN => n2767);
   U2827 : AOI211_X1 port map( C1 => n745, C2 => n2907, A => n2914, B => n2872,
                           ZN => n2766);
   U2828 : OR2_X1 port map( A1 => n2767, A2 => n2766, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U2829 : AOI211_X1 port map( C1 => n2768, C2 => n2899, A => n2969, B => n2906
                           , ZN => n2770);
   U2830 : AOI211_X1 port map( C1 => n752, C2 => n2901, A => n2908, B => n2872,
                           ZN => n2769);
   U2831 : OR2_X1 port map( A1 => n2770, A2 => n2769, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U2832 : AOI211_X1 port map( C1 => n2771, C2 => n2893, A => n2969, B => n2900
                           , ZN => n2773);
   U2833 : AOI211_X1 port map( C1 => n744, C2 => n2895, A => n2902, B => n2966,
                           ZN => n2772);
   U2834 : OR2_X1 port map( A1 => n2773, A2 => n2772, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U2835 : AOI211_X1 port map( C1 => n2774, C2 => n2887, A => n2920, B => n2894
                           , ZN => n2776);
   U2836 : AOI211_X1 port map( C1 => n743, C2 => n2889, A => n2896, B => n2966,
                           ZN => n2775);
   U2837 : OR2_X1 port map( A1 => n2776, A2 => n2775, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U2838 : AOI211_X1 port map( C1 => n2777, C2 => n2881, A => n2920, B => n2888
                           , ZN => n2779);
   U2839 : AOI211_X1 port map( C1 => n742, C2 => n2883, A => n2890, B => n2872,
                           ZN => n2778);
   U2840 : OR2_X1 port map( A1 => n2779, A2 => n2778, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U2841 : AOI211_X1 port map( C1 => n2780, C2 => n2875, A => n2920, B => n2882
                           , ZN => n2782);
   U2842 : AOI211_X1 port map( C1 => n741, C2 => n2877, A => n2884, B => n2966,
                           ZN => n2781);
   U2843 : OR2_X1 port map( A1 => n2782, A2 => n2781, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U2844 : NOR3_X1 port map( A1 => n3017, A2 => n2833, A3 => n3086, ZN => 
                           cu_i_cmd_word_7_port);
   U2845 : NOR3_X1 port map( A1 => n3085, A2 => n3089, A3 => n2784, ZN => n2835
                           );
   U2846 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => n737
                           , ZN => n2826);
   U2847 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n2826, A3 => n3091, ZN => n2810);
   U2848 : AOI21_X1 port map( B1 => n3085, B2 => n3086, A => n2810, ZN => n2818
                           );
   U2849 : NAND2_X1 port map( A1 => n2826, A2 => n3089, ZN => n2832);
   U2850 : AOI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n2833, A => n2832, ZN => n2783);
   U2851 : NOR3_X1 port map( A1 => n2835, A2 => n2818, A3 => n2783, ZN => n2853
                           );
   U2852 : OAI21_X1 port map( B1 => n2833, B2 => n2784, A => n2853, ZN => n2851
                           );
   U2853 : AND2_X1 port map( A1 => n2794, A2 => n3015, ZN => n3042);
   U2854 : INV_X1 port map( A => n3042, ZN => n3105);
   U2855 : INV_X1 port map( A => n3015, ZN => n3104);
   U2856 : NAND2_X1 port map( A1 => n2792, A2 => n2856, ZN => n2849);
   U2857 : INV_X1 port map( A => n2972, ZN => n2971);
   U2858 : AOI221_X1 port map( B1 => n2971, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n2972, C2 =>
                           curr_instruction_to_cu_i_15_port, A => n3104, ZN => 
                           n2786);
   U2859 : INV_X1 port map( A => n2786, ZN => n2708);
   U2860 : AOI221_X1 port map( B1 => n2971, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n2972, C2 =>
                           curr_instruction_to_cu_i_14_port, A => n3104, ZN => 
                           n2787);
   U2861 : INV_X1 port map( A => n2787, ZN => n2707);
   U2862 : AOI221_X1 port map( B1 => n2971, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n2972, C2 =>
                           curr_instruction_to_cu_i_12_port, A => n3104, ZN => 
                           n2788);
   U2863 : INV_X1 port map( A => n2788, ZN => n2706);
   U2864 : AOI221_X1 port map( B1 => n2971, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n2972, C2 =>
                           curr_instruction_to_cu_i_11_port, A => n3104, ZN => 
                           n2789);
   U2865 : INV_X1 port map( A => n2789, ZN => n2705);
   U2866 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_1_port, B1
                           => cu_i_cw1_1_port, B2 => n3093, ZN => n2801);
   U2867 : INV_X1 port map( A => n704, ZN => n2866);
   U2868 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_3_port, B1
                           => cu_i_cw1_3_port, B2 => n2866, ZN => n2798);
   U2869 : AOI21_X1 port map( B1 => n2807, B2 => n2801, A => n2798, ZN => n2790
                           );
   U2870 : NOR2_X1 port map( A1 => n2799, A2 => n2790, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U2871 : INV_X1 port map( A => n2798, ZN => n2806);
   U2872 : OAI211_X1 port map( C1 => n2799, C2 => n2801, A => n2806, B => n2807
                           , ZN => n2791);
   U2873 : INV_X1 port map( A => n2791, ZN => n2704);
   U2874 : INV_X1 port map( A => n2792, ZN => n2862);
   U2875 : OAI222_X1 port map( A1 => n3086, A2 => n3015, B1 => n2849, B2 => 
                           n2796, C1 => n2862, C2 => n2853, ZN => n311);
   U2876 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n311, ZN => 
                           cu_i_cmd_word_1_port);
   U2877 : OAI22_X1 port map( A1 => n3093, A2 => cu_i_cw3_6_port, B1 => 
                           cu_i_cw2_6_port, B2 => n704, ZN => n2793);
   U2878 : INV_X1 port map( A => n2793, ZN => n2712);
   U2879 : NAND2_X1 port map( A1 => n2794, A2 => n2971, ZN => enable_rf_i);
   U2880 : INV_X1 port map( A => n2849, ZN => n2795);
   U2881 : NAND2_X1 port map( A1 => n2796, A2 => n2795, ZN => n2844);
   U2882 : INV_X1 port map( A => n3042, ZN => n3106);
   U2883 : AND2_X1 port map( A1 => n3106, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U2884 : INV_X1 port map( A => n2797, ZN => DRAM_READNOTWRITE);
   U2885 : AOI22_X1 port map( A1 => n704, A2 => n3042, B1 => n2319, B2 => n2866
                           , ZN => n3045);
   U2886 : MUX2_X1 port map( A => datapath_i_val_b_i_0_port, B => 
                           datapath_i_val_immediate_i_0_port, S => n3045, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U2887 : CLKBUF_X1 port map( A => n3045, Z => n3047);
   U2888 : MUX2_X1 port map( A => datapath_i_val_b_i_1_port, B => 
                           datapath_i_val_immediate_i_1_port, S => n3047, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U2889 : AOI21_X1 port map( B1 => n2807, B2 => n2799, A => n2798, ZN => n2800
                           );
   U2890 : NOR2_X1 port map( A1 => n2801, A2 => n2800, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U2891 : NOR2_X1 port map( A1 => n3088, A2 => n2844, ZN => cu_i_N273);
   U2892 : INV_X1 port map( A => n2844, ZN => n2974);
   U2893 : AOI221_X1 port map( B1 => cu_i_n25, B2 => n2974, C1 => cu_i_n26, C2 
                           => n2974, A => cu_i_N273, ZN => n2802);
   U2894 : INV_X1 port map( A => n2802, ZN => n2805);
   U2895 : NOR2_X1 port map( A1 => cu_i_n125, A2 => n2844, ZN => n2803);
   U2896 : NAND2_X1 port map( A1 => n2803, A2 => n3095, ZN => n2842);
   U2897 : NOR2_X1 port map( A1 => cu_i_n25, A2 => n2842, ZN => n2804);
   U2898 : MUX2_X1 port map( A => n2805, B => n2804, S => cu_i_n124, Z => 
                           cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U2900 : MUX2_X1 port map( A => datapath_i_val_b_i_2_port, B => 
                           datapath_i_val_immediate_i_2_port, S => n3047, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U2901 : NOR2_X1 port map( A1 => n2807, A2 => n2806, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U2902 : NAND2_X1 port map( A1 => n3042, A2 => n2849, ZN => cu_i_N278);
   U2903 : NOR2_X1 port map( A1 => n2833, A2 => 
                           curr_instruction_to_cu_i_26_port, ZN => n2827);
   U2904 : INV_X1 port map( A => n2827, ZN => n3016);
   U2905 : INV_X1 port map( A => n2856, ZN => n2858);
   U2906 : NAND2_X1 port map( A1 => n3098, A2 => n3090, ZN => n2808);
   U2907 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => n3094
                           , A3 => n2858, A4 => n2808, ZN => n2837);
   U2908 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_5_port, A2 => 
                           n2856, A3 => n3090, A4 => n3097, ZN => n2825);
   U2909 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n2809
                           , A3 => n2825, ZN => n2815);
   U2910 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n3086, ZN => n2812);
   U2911 : INV_X1 port map( A => n2810, ZN => n2811);
   U2912 : AOI21_X1 port map( B1 => n2812, B2 => n2811, A => n2835, ZN => n2813
                           );
   U2913 : INV_X1 port map( A => n2813, ZN => n2814);
   U2914 : AOI211_X1 port map( C1 => n2837, C2 => n2824, A => n2815, B => n2814
                           , ZN => n2817);
   U2915 : OAI211_X1 port map( C1 => n2832, C2 => n3016, A => n2817, B => n2816
                           , ZN => cu_i_N265);
   U2916 : MUX2_X1 port map( A => datapath_i_val_b_i_3_port, B => 
                           datapath_i_val_immediate_i_3_port, S => n3045, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U2917 : OR2_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           curr_instruction_to_cu_i_2_port, ZN => n2848);
   U2918 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           n2848, ZN => n2820);
   U2919 : INV_X1 port map( A => n2818, ZN => n2819);
   U2920 : OAI21_X1 port map( B1 => n2825, B2 => n2820, A => n2819, ZN => 
                           cu_i_N267);
   U2921 : NOR2_X1 port map( A1 => n3093, A2 => n1152, ZN => n2821);
   U2922 : NOR2_X1 port map( A1 => n704, A2 => cu_i_cw1_4_port, ZN => n2850);
   U2923 : NOR2_X1 port map( A1 => n2821, A2 => n2850, ZN => n2822);
   U2924 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n2822, ZN => n3084);
   U2925 : INV_X1 port map( A => n2822, ZN => n3069);
   U2926 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n3069, ZN => n3082);
   U2927 : CLKBUF_X1 port map( A => n3082, Z => n3071);
   U2928 : CLKBUF_X1 port map( A => n3069, Z => n3081);
   U2929 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n3081, ZN => n2823);
   U2930 : OAI21_X1 port map( B1 => n691, B2 => n3073, A => n2823, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U2931 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_4_port, A3 => n2824, ZN => 
                           n2845);
   U2932 : NOR2_X1 port map( A1 => n3094, A2 => n2825, ZN => n2838);
   U2933 : AOI21_X1 port map( B1 => n2845, B2 => n2856, A => n2838, ZN => n2830
                           );
   U2934 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => 
                           n3091, A3 => n2832, ZN => n2831);
   U2935 : AOI21_X1 port map( B1 => n2827, B2 => n2826, A => n2831, ZN => n2829
                           );
   U2936 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n2835, B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           n2837, ZN => n2828);
   U2937 : OAI211_X1 port map( C1 => curr_instruction_to_cu_i_0_port, C2 => 
                           n2830, A => n2829, B => n2828, ZN => cu_i_N264);
   U2938 : INV_X1 port map( A => n2831, ZN => n2846);
   U2939 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_5_port, A2 => 
                           n3097, ZN => n2836);
   U2940 : NOR3_X1 port map( A1 => n2833, A2 => n3086, A3 => n2832, ZN => n2834
                           );
   U2941 : AOI211_X1 port map( C1 => n2837, C2 => n2836, A => n2835, B => n2834
                           , ZN => n2840);
   U2942 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           n2838, A3 => n3098, ZN => n2839);
   U2943 : OAI211_X1 port map( C1 => n2846, C2 => n3085, A => n2840, B => n2839
                           , ZN => cu_i_N266);
   U2944 : NAND2_X1 port map( A1 => n704, A2 => n2844, ZN => cu_i_N274);
   U2945 : AOI221_X1 port map( B1 => cu_i_n125, B2 => cu_i_n26, C1 => n3088, C2
                           => n3095, A => n2844, ZN => cu_i_N275);
   U2946 : OAI21_X1 port map( B1 => cu_i_n26, B2 => cu_i_n125, A => n2974, ZN 
                           => n2841);
   U2947 : AOI22_X1 port map( A1 => cu_i_n25, A2 => n2842, B1 => n2841, B2 => 
                           n3102, ZN => cu_i_N276);
   U2948 : INV_X1 port map( A => n2843, ZN => n2975);
   U2949 : AOI211_X1 port map( C1 => n704, C2 => cu_i_n145, A => n2975, B => 
                           n2844, ZN => cu_i_N279);
   U2950 : INV_X1 port map( A => n2845, ZN => n2847);
   U2951 : OAI33_X1 port map( A1 => n2849, A2 => n2848, A3 => n2847, B1 => 
                           n2862, B2 => n2846, B3 => 
                           curr_instruction_to_cu_i_28_port, ZN => 
                           cu_i_cmd_word_8_port);
   U2952 : MUX2_X1 port map( A => cu_i_cmd_word_8_port, B => cu_i_cw1_12_port, 
                           S => n2866, Z => alu_cin_i);
   U2953 : AOI21_X1 port map( B1 => n756, B2 => n704, A => n2850, ZN => 
                           cu_i_cw1_i_4_port);
   U2954 : MUX2_X1 port map( A => cu_i_cw2_7_port, B => cu_i_cw1_7_port, S => 
                           n3093, Z => cu_i_cw1_i_7_port);
   U2955 : MUX2_X1 port map( A => cu_i_cw2_8_port, B => cu_i_cw1_8_port, S => 
                           n3093, Z => cu_i_cw1_i_8_port);
   U2956 : INV_X1 port map( A => n2851, ZN => n2859);
   U2957 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_14_port, A2 => 
                           curr_instruction_to_cu_i_15_port, A3 => 
                           curr_instruction_to_cu_i_11_port, A4 => 
                           curr_instruction_to_cu_i_12_port, ZN => n2852);
   U2958 : NAND2_X1 port map( A1 => n740, A2 => n2852, ZN => n2857);
   U2959 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_19_port, A2 => 
                           curr_instruction_to_cu_i_20_port, A3 => 
                           curr_instruction_to_cu_i_16_port, A4 => 
                           curr_instruction_to_cu_i_17_port, ZN => n2854);
   U2960 : AOI21_X1 port map( B1 => n697, B2 => n2854, A => n2853, ZN => n2855)
                           ;
   U2961 : AOI221_X1 port map( B1 => n2859, B2 => n2858, C1 => n2857, C2 => 
                           n2856, A => n2855, ZN => n2863);
   U2962 : OAI211_X1 port map( C1 => n2863, C2 => n2862, A => n2861, B => n2860
                           , ZN => cu_i_n209);
   U2963 : NOR2_X1 port map( A1 => cu_i_n123, A2 => cu_i_n23, ZN => cu_i_n210);
   U2964 : AOI22_X1 port map( A1 => n704, A2 => n699, B1 => n3103, B2 => n3093,
                           ZN => cu_i_n131);
   U2965 : MUX2_X1 port map( A => cu_i_cw2_6_port, B => cu_i_cw1_6_port, S => 
                           n2866, Z => cu_i_n127);
   U2966 : MUX2_X1 port map( A => cu_i_cw2_5_port, B => cu_i_cw1_5_port, S => 
                           n2866, Z => cu_i_n126);
   U2967 : MUX2_X1 port map( A => curr_instruction_to_cu_i_31_port, B => 
                           IRAM_DATA(31), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U2968 : MUX2_X1 port map( A => curr_instruction_to_cu_i_30_port, B => 
                           IRAM_DATA(30), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U2969 : MUX2_X1 port map( A => n3100, B => IRAM_DATA(29), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U2970 : MUX2_X1 port map( A => curr_instruction_to_cu_i_28_port, B => 
                           IRAM_DATA(28), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U2971 : MUX2_X1 port map( A => curr_instruction_to_cu_i_27_port, B => 
                           IRAM_DATA(27), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U2972 : MUX2_X1 port map( A => curr_instruction_to_cu_i_26_port, B => 
                           IRAM_DATA(26), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U2973 : MUX2_X1 port map( A => datapath_i_n9, B => IRAM_DATA(25), S => n2866
                           , Z => datapath_i_fetch_stage_dp_n63);
   U2974 : MUX2_X1 port map( A => datapath_i_n10, B => IRAM_DATA(24), S => 
                           n2866, Z => datapath_i_fetch_stage_dp_n62);
   U2975 : MUX2_X1 port map( A => datapath_i_n11, B => IRAM_DATA(23), S => 
                           n2866, Z => datapath_i_fetch_stage_dp_n61);
   U2976 : MUX2_X1 port map( A => datapath_i_n12, B => IRAM_DATA(22), S => 
                           n3093, Z => datapath_i_fetch_stage_dp_n60);
   U2977 : MUX2_X1 port map( A => datapath_i_n13, B => IRAM_DATA(21), S => 
                           n3093, Z => datapath_i_fetch_stage_dp_n59);
   U2978 : MUX2_X1 port map( A => curr_instruction_to_cu_i_20_port, B => 
                           IRAM_DATA(20), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U2979 : MUX2_X1 port map( A => curr_instruction_to_cu_i_19_port, B => 
                           IRAM_DATA(19), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U2980 : NAND2_X1 port map( A1 => n3093, A2 => IRAM_DATA(18), ZN => n2864);
   U2981 : OAI21_X1 port map( B1 => n3093, B2 => n697, A => n2864, ZN => 
                           datapath_i_fetch_stage_dp_n56);
   U2982 : MUX2_X1 port map( A => curr_instruction_to_cu_i_17_port, B => 
                           IRAM_DATA(17), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U2983 : MUX2_X1 port map( A => curr_instruction_to_cu_i_16_port, B => 
                           IRAM_DATA(16), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U2984 : MUX2_X1 port map( A => curr_instruction_to_cu_i_15_port, B => 
                           IRAM_DATA(15), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U2985 : MUX2_X1 port map( A => curr_instruction_to_cu_i_14_port, B => 
                           IRAM_DATA(14), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U2986 : NAND2_X1 port map( A1 => n3093, A2 => IRAM_DATA(13), ZN => n2865);
   U2987 : OAI21_X1 port map( B1 => n2866, B2 => n740, A => n2865, ZN => 
                           datapath_i_fetch_stage_dp_n51);
   U2988 : MUX2_X1 port map( A => curr_instruction_to_cu_i_12_port, B => 
                           IRAM_DATA(12), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U2989 : MUX2_X1 port map( A => curr_instruction_to_cu_i_11_port, B => 
                           IRAM_DATA(11), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U2990 : MUX2_X1 port map( A => datapath_i_n14, B => IRAM_DATA(10), S => 
                           n2866, Z => datapath_i_fetch_stage_dp_n48);
   U2991 : MUX2_X1 port map( A => datapath_i_n15, B => IRAM_DATA(9), S => n2866
                           , Z => datapath_i_fetch_stage_dp_n47);
   U2992 : MUX2_X1 port map( A => datapath_i_n16, B => IRAM_DATA(8), S => n3093
                           , Z => datapath_i_fetch_stage_dp_n46);
   U2993 : MUX2_X1 port map( A => datapath_i_n17, B => IRAM_DATA(7), S => n2866
                           , Z => datapath_i_fetch_stage_dp_n45);
   U2994 : MUX2_X1 port map( A => datapath_i_n18, B => IRAM_DATA(6), S => n2866
                           , Z => datapath_i_fetch_stage_dp_n44);
   U2995 : MUX2_X1 port map( A => curr_instruction_to_cu_i_5_port, B => 
                           IRAM_DATA(5), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U2996 : MUX2_X1 port map( A => curr_instruction_to_cu_i_4_port, B => 
                           IRAM_DATA(4), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U2997 : MUX2_X1 port map( A => curr_instruction_to_cu_i_3_port, B => 
                           IRAM_DATA(3), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U2998 : MUX2_X1 port map( A => curr_instruction_to_cu_i_2_port, B => 
                           IRAM_DATA(2), S => n3093, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U2999 : MUX2_X1 port map( A => curr_instruction_to_cu_i_1_port, B => 
                           IRAM_DATA(1), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U3000 : MUX2_X1 port map( A => curr_instruction_to_cu_i_0_port, B => 
                           IRAM_DATA(0), S => n2866, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U3001 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_0_port, ZN => 
                           n2867);
   U3002 : OAI21_X1 port map( B1 => n733, B2 => n2963, A => n2867, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U3003 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N39_port, B => 
                           datapath_i_fetch_stage_dp_N5, S => n2872, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U3004 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_1_port, B1 => n2954, B2 
                           => datapath_i_new_pc_value_decode_1_port, ZN => 
                           n2868);
   U3005 : OAI21_X1 port map( B1 => n734, B2 => n2963, A => n2868, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U3006 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N40_port, B => 
                           datapath_i_fetch_stage_dp_N6, S => n2872, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U3007 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n2869, ZN => n2870);
   U3008 : AOI22_X1 port map( A1 => n2969, A2 => n2870, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n2966, ZN => datapath_i_fetch_stage_dp_n35);
   U3009 : OAI21_X1 port map( B1 => n2871, B2 => IRAM_ADDRESS_3_port, A => 
                           n2920, ZN => n2874);
   U3010 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n2876);
   U3011 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           B2 => datapath_i_new_pc_value_mem_stage_i_3_port, A 
                           => n2872, ZN => n2873);
   U3012 : OAI22_X1 port map( A1 => n2878, A2 => n2874, B1 => n2876, B2 => 
                           n2873, ZN => datapath_i_fetch_stage_dp_n34);
   U3013 : OAI211_X1 port map( C1 => n2876, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n2966, B => n2875, ZN => n2880);
   U3014 : OAI211_X1 port map( C1 => n2878, C2 => IRAM_ADDRESS_4_port, A => 
                           n2969, B => n2877, ZN => n2879);
   U3015 : NAND2_X1 port map( A1 => n2880, A2 => n2879, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U3016 : OAI211_X1 port map( C1 => n2882, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n2966, B => n2881, ZN => n2886);
   U3017 : OAI211_X1 port map( C1 => n2884, C2 => IRAM_ADDRESS_6_port, A => 
                           n2969, B => n2883, ZN => n2885);
   U3018 : NAND2_X1 port map( A1 => n2886, A2 => n2885, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U3019 : OAI211_X1 port map( C1 => n2888, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n2966, B => n2887, ZN => n2892);
   U3020 : OAI211_X1 port map( C1 => n2890, C2 => IRAM_ADDRESS_8_port, A => 
                           n2969, B => n2889, ZN => n2891);
   U3021 : NAND2_X1 port map( A1 => n2892, A2 => n2891, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U3022 : OAI211_X1 port map( C1 => n2894, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n2966, B => n2893, ZN => n2898);
   U3023 : OAI211_X1 port map( C1 => n2896, C2 => IRAM_ADDRESS_10_port, A => 
                           n2969, B => n2895, ZN => n2897);
   U3024 : NAND2_X1 port map( A1 => n2898, A2 => n2897, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U3025 : OAI211_X1 port map( C1 => n2900, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n2966, B => n2899, ZN => n2904);
   U3026 : OAI211_X1 port map( C1 => n2902, C2 => IRAM_ADDRESS_12_port, A => 
                           n2920, B => n2901, ZN => n2903);
   U3027 : NAND2_X1 port map( A1 => n2904, A2 => n2903, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U3028 : OAI211_X1 port map( C1 => n2906, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n2966, B => n2905, ZN => n2910);
   U3029 : OAI211_X1 port map( C1 => n2908, C2 => IRAM_ADDRESS_14_port, A => 
                           n2920, B => n2907, ZN => n2909);
   U3030 : NAND2_X1 port map( A1 => n2910, A2 => n2909, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U3031 : OAI211_X1 port map( C1 => n2912, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n2966, B => n2911, ZN => n2916);
   U3032 : OAI211_X1 port map( C1 => n2914, C2 => IRAM_ADDRESS_16_port, A => 
                           n2920, B => n2913, ZN => n2915);
   U3033 : NAND2_X1 port map( A1 => n2916, A2 => n2915, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U3034 : OAI211_X1 port map( C1 => n2918, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n2966, B => n2917, ZN => n2923);
   U3035 : OAI211_X1 port map( C1 => n2921, C2 => IRAM_ADDRESS_18_port, A => 
                           n2920, B => n2919, ZN => n2922);
   U3036 : NAND2_X1 port map( A1 => n2923, A2 => n2922, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U3037 : OAI211_X1 port map( C1 => n2925, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n2966, B => n2924, ZN => n2929);
   U3038 : OAI211_X1 port map( C1 => n2927, C2 => IRAM_ADDRESS_20_port, A => 
                           n2969, B => n2926, ZN => n2928);
   U3039 : NAND2_X1 port map( A1 => n2929, A2 => n2928, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U3040 : OAI211_X1 port map( C1 => n2931, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n2966, B => n2930, ZN => n2935);
   U3041 : OAI211_X1 port map( C1 => n2933, C2 => IRAM_ADDRESS_22_port, A => 
                           n2969, B => n2932, ZN => n2934);
   U3042 : NAND2_X1 port map( A1 => n2935, A2 => n2934, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U3043 : OAI211_X1 port map( C1 => n2937, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n2966, B => n2936, ZN => n2941);
   U3044 : OAI211_X1 port map( C1 => n2939, C2 => IRAM_ADDRESS_24_port, A => 
                           n2969, B => n2938, ZN => n2940);
   U3045 : NAND2_X1 port map( A1 => n2941, A2 => n2940, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U3046 : OAI211_X1 port map( C1 => n2943, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n2966, B => n2942, ZN => n2947);
   U3047 : OAI211_X1 port map( C1 => n2945, C2 => IRAM_ADDRESS_26_port, A => 
                           n2969, B => n2944, ZN => n2946);
   U3048 : NAND2_X1 port map( A1 => n2947, A2 => n2946, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U3049 : OAI211_X1 port map( C1 => n2949, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n2966, B => n2948, ZN => n2953);
   U3050 : OAI211_X1 port map( C1 => n2951, C2 => IRAM_ADDRESS_28_port, A => 
                           n2969, B => n2950, ZN => n2952);
   U3051 : NAND2_X1 port map( A1 => n2953, A2 => n2952, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U3052 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_30_port, B1 => n2954, B2
                           => datapath_i_new_pc_value_decode_30_port, ZN => 
                           n2955);
   U3053 : OAI21_X1 port map( B1 => n727, B2 => n2963, A => n2955, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   U3054 : NAND2_X1 port map( A1 => n2956, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n2965);
   U3055 : OAI211_X1 port map( C1 => n2956, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n2966, B => n2965, ZN => n2959);
   U3056 : NAND2_X1 port map( A1 => n2957, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n2964);
   U3057 : OAI211_X1 port map( C1 => n2957, C2 => IRAM_ADDRESS_30_port, A => 
                           n2969, B => n2964, ZN => n2958);
   U3058 : NAND2_X1 port map( A1 => n2959, A2 => n2958, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U3059 : AOI22_X1 port map( A1 => n2961, A2 => 
                           datapath_i_alu_output_val_i_31_port, B1 => 
                           datapath_i_new_pc_value_decode_31_port, B2 => n2960,
                           ZN => n2962);
   U3060 : OAI21_X1 port map( B1 => n703, B2 => n2963, A => n2962, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U3061 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n2964, Z => n2968)
                           ;
   U3062 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n2965, Z => n2967);
   U3063 : AOI22_X1 port map( A1 => n2969, A2 => n2968, B1 => n2967, B2 => 
                           n2966, ZN => datapath_i_fetch_stage_dp_n2);
   U3064 : OAI21_X1 port map( B1 => n737, B2 => n2970, A => n2971, ZN => 
                           read_rf_p2_i);
   U3065 : OAI221_X1 port map( B1 => n2972, B2 => n697, C1 => n2971, C2 => n740
                           , A => n3015, ZN => datapath_i_decode_stage_dp_n78);
   U3066 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ZN => n2973);
   U3067 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n2973, ZN => n2989);
   U3068 : INV_X1 port map( A => n2989, ZN => n2998);
   U3069 : AND2_X2 port map( A1 => n2998, A2 => n2976, ZN => n3012);
   U3070 : NOR2_X1 port map( A1 => n2989, A2 => n2976, ZN => n3011);
   U3071 : CLKBUF_X1 port map( A => n3011, Z => n3002);
   U3072 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_0_port, ZN => n2977
                           );
   U3073 : OAI21_X1 port map( B1 => n733, B2 => n2998, A => n2977, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U3074 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_1_port, ZN => n2978
                           );
   U3075 : OAI21_X1 port map( B1 => n734, B2 => n2998, A => n2978, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U3076 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_2_port, ZN => n2979
                           );
   U3077 : OAI21_X1 port map( B1 => n728, B2 => n2998, A => n2979, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U3078 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_3_port, ZN => n2980
                           );
   U3079 : OAI21_X1 port map( B1 => n729, B2 => n2998, A => n2980, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U3080 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_4_port, ZN => n2981
                           );
   U3081 : OAI21_X1 port map( B1 => n730, B2 => n2998, A => n2981, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U3082 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_5_port, ZN => n2982
                           );
   U3083 : OAI21_X1 port map( B1 => n731, B2 => n2998, A => n2982, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U3084 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_6_port, ZN => n2983
                           );
   U3085 : OAI21_X1 port map( B1 => n732, B2 => n2998, A => n2983, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U3086 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_7_port, ZN => n2984
                           );
   U3087 : OAI21_X1 port map( B1 => n705, B2 => n2998, A => n2984, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U3088 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_8_port, ZN => n2985
                           );
   U3089 : OAI21_X1 port map( B1 => n706, B2 => n2998, A => n2985, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U3090 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_9_port, ZN => n2986
                           );
   U3091 : OAI21_X1 port map( B1 => n707, B2 => n2998, A => n2986, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U3092 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => 
                           n2987);
   U3093 : OAI21_X1 port map( B1 => n708, B2 => n2998, A => n2987, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U3094 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => 
                           n2988);
   U3095 : OAI21_X1 port map( B1 => n709, B2 => n2998, A => n2988, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U3096 : INV_X1 port map( A => n2989, ZN => n3014);
   U3097 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => 
                           n2990);
   U3098 : OAI21_X1 port map( B1 => n710, B2 => n3014, A => n2990, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U3099 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => 
                           n2991);
   U3100 : OAI21_X1 port map( B1 => n711, B2 => n2998, A => n2991, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U3101 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => 
                           n2992);
   U3102 : OAI21_X1 port map( B1 => n712, B2 => n3014, A => n2992, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U3103 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => 
                           n2993);
   U3104 : OAI21_X1 port map( B1 => n713, B2 => n2998, A => n2993, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U3105 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => 
                           n2994);
   U3106 : OAI21_X1 port map( B1 => n714, B2 => n3014, A => n2994, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U3107 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => 
                           n2995);
   U3108 : OAI21_X1 port map( B1 => n715, B2 => n2998, A => n2995, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U3109 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => 
                           n2996);
   U3110 : OAI21_X1 port map( B1 => n716, B2 => n3014, A => n2996, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U3111 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => 
                           n2997);
   U3112 : OAI21_X1 port map( B1 => n717, B2 => n2998, A => n2997, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U3113 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => 
                           n2999);
   U3114 : OAI21_X1 port map( B1 => n718, B2 => n3014, A => n2999, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U3115 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => 
                           n3000);
   U3116 : OAI21_X1 port map( B1 => n719, B2 => n3014, A => n3000, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U3117 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => 
                           n3001);
   U3118 : OAI21_X1 port map( B1 => n720, B2 => n3014, A => n3001, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U3119 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n3002, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => 
                           n3003);
   U3120 : OAI21_X1 port map( B1 => n721, B2 => n3014, A => n3003, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U3121 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => 
                           n3004);
   U3122 : OAI21_X1 port map( B1 => n722, B2 => n3014, A => n3004, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U3123 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => 
                           n3005);
   U3124 : OAI21_X1 port map( B1 => n723, B2 => n3014, A => n3005, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U3125 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => 
                           n3006);
   U3126 : OAI21_X1 port map( B1 => n691, B2 => n3014, A => n3006, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U3127 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => 
                           n3007);
   U3128 : OAI21_X1 port map( B1 => n724, B2 => n3014, A => n3007, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U3129 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => 
                           n3008);
   U3130 : OAI21_X1 port map( B1 => n725, B2 => n3014, A => n3008, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U3131 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => 
                           n3009);
   U3132 : OAI21_X1 port map( B1 => n726, B2 => n3014, A => n3009, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U3133 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => 
                           n3010);
   U3134 : OAI21_X1 port map( B1 => n727, B2 => n3014, A => n3010, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U3135 : AOI22_X1 port map( A1 => n3012, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n3011, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => 
                           n3013);
   U3136 : OAI21_X1 port map( B1 => n703, B2 => n3014, A => n3013, ZN => 
                           datapath_i_decode_stage_dp_n12);
   U3137 : OAI21_X1 port map( B1 => n3017, B2 => n3016, A => n3015, ZN => 
                           cu_i_cmd_word_6_port);
   U3138 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_6_port, B1 => 
                           cu_i_cw1_10_port, B2 => n3093, ZN => n3031);
   U3139 : NOR4_X1 port map( A1 => datapath_i_val_a_i_14_port, A2 => 
                           datapath_i_val_a_i_15_port, A3 => 
                           datapath_i_val_a_i_16_port, A4 => 
                           datapath_i_val_a_i_17_port, ZN => n3021);
   U3140 : NOR4_X1 port map( A1 => datapath_i_val_a_i_18_port, A2 => 
                           datapath_i_val_a_i_19_port, A3 => 
                           datapath_i_val_a_i_20_port, A4 => 
                           datapath_i_val_a_i_21_port, ZN => n3020);
   U3141 : NOR4_X1 port map( A1 => datapath_i_val_a_i_26_port, A2 => 
                           datapath_i_val_a_i_7_port, A3 => 
                           datapath_i_val_a_i_8_port, A4 => 
                           datapath_i_val_a_i_9_port, ZN => n3019);
   U3142 : NOR4_X1 port map( A1 => datapath_i_val_a_i_10_port, A2 => 
                           datapath_i_val_a_i_11_port, A3 => 
                           datapath_i_val_a_i_12_port, A4 => 
                           datapath_i_val_a_i_13_port, ZN => n3018);
   U3143 : NAND4_X1 port map( A1 => n3021, A2 => n3020, A3 => n3019, A4 => 
                           n3018, ZN => n3027);
   U3144 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n3025);
   U3145 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n3024);
   U3146 : NOR4_X1 port map( A1 => datapath_i_val_a_i_22_port, A2 => 
                           datapath_i_val_a_i_23_port, A3 => 
                           datapath_i_val_a_i_24_port, A4 => 
                           datapath_i_val_a_i_25_port, ZN => n3023);
   U3147 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n3022);
   U3148 : NAND4_X1 port map( A1 => n3025, A2 => n3024, A3 => n3023, A4 => 
                           n3022, ZN => n3026);
   U3149 : NOR2_X1 port map( A1 => n3027, A2 => n3026, ZN => n3029);
   U3150 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_7_port, B1 => 
                           cu_i_cw1_11_port, B2 => n3093, ZN => n3028);
   U3151 : NAND2_X1 port map( A1 => n3029, A2 => n3028, ZN => n3030);
   U3152 : OAI22_X1 port map( A1 => n3031, A2 => n3030, B1 => n3029, B2 => 
                           n3028, ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U3153 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, S 
                           => n3106, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U3154 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U3155 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, S 
                           => n3106, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U3156 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U3157 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, S 
                           => n3106, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U3158 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U3159 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U3160 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U3161 : NAND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
                           A2 => n3106, ZN => n3044);
   U3162 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
                           ZN => n3032);
   U3163 : NAND2_X1 port map( A1 => n3044, A2 => n3032, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U3164 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
                           ZN => n3033);
   U3165 : NAND2_X1 port map( A1 => n3044, A2 => n3033, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U3166 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
                           ZN => n3034);
   U3167 : NAND2_X1 port map( A1 => n3044, A2 => n3034, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U3168 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
                           ZN => n3035);
   U3169 : NAND2_X1 port map( A1 => n3044, A2 => n3035, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U3170 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
                           ZN => n3036);
   U3171 : NAND2_X1 port map( A1 => n3044, A2 => n3036, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U3172 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
                           ZN => n3037);
   U3173 : NAND2_X1 port map( A1 => n3044, A2 => n3037, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U3174 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
                           ZN => n3038);
   U3175 : NAND2_X1 port map( A1 => n3044, A2 => n3038, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U3176 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
                           ZN => n3039);
   U3177 : NAND2_X1 port map( A1 => n3044, A2 => n3039, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U3178 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
                           ZN => n3040);
   U3179 : NAND2_X1 port map( A1 => n3044, A2 => n3040, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U3180 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
                           ZN => n3041);
   U3181 : NAND2_X1 port map( A1 => n3044, A2 => n3041, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U3182 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U3183 : NAND2_X1 port map( A1 => n3042, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
                           ZN => n3043);
   U3184 : NAND2_X1 port map( A1 => n3044, A2 => n3043, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U3185 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U3186 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U3187 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U3188 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U3189 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U3190 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, S 
                           => n3105, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U3191 : MUX2_X1 port map( A => datapath_i_val_b_i_7_port, B => 
                           datapath_i_val_immediate_i_7_port, S => n3045, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U3192 : MUX2_X1 port map( A => datapath_i_val_b_i_8_port, B => 
                           datapath_i_val_immediate_i_8_port, S => n3045, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U3193 : MUX2_X1 port map( A => datapath_i_val_b_i_9_port, B => 
                           datapath_i_val_immediate_i_9_port, S => n3045, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U3194 : MUX2_X1 port map( A => datapath_i_val_b_i_10_port, B => 
                           datapath_i_val_immediate_i_10_port, S => n3045, Z =>
                           datapath_i_execute_stage_dp_opb_10_port);
   U3195 : MUX2_X1 port map( A => datapath_i_val_b_i_11_port, B => 
                           datapath_i_val_immediate_i_11_port, S => n3045, Z =>
                           datapath_i_execute_stage_dp_opb_11_port);
   U3196 : MUX2_X1 port map( A => datapath_i_val_b_i_12_port, B => 
                           datapath_i_val_immediate_i_12_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_12_port);
   U3197 : MUX2_X1 port map( A => datapath_i_val_b_i_13_port, B => 
                           datapath_i_val_immediate_i_13_port, S => n3045, Z =>
                           datapath_i_execute_stage_dp_opb_13_port);
   U3198 : MUX2_X1 port map( A => datapath_i_val_b_i_14_port, B => 
                           datapath_i_val_immediate_i_14_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_14_port);
   U3199 : MUX2_X1 port map( A => datapath_i_val_b_i_15_port, B => 
                           datapath_i_val_immediate_i_15_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_15_port);
   U3200 : MUX2_X1 port map( A => datapath_i_val_b_i_16_port, B => 
                           datapath_i_val_immediate_i_16_port, S => n3045, Z =>
                           datapath_i_execute_stage_dp_opb_16_port);
   U3201 : MUX2_X1 port map( A => datapath_i_val_b_i_17_port, B => 
                           datapath_i_val_immediate_i_17_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_17_port);
   U3202 : MUX2_X1 port map( A => datapath_i_val_b_i_18_port, B => 
                           datapath_i_val_immediate_i_18_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_18_port);
   U3203 : MUX2_X1 port map( A => datapath_i_val_b_i_19_port, B => 
                           datapath_i_val_immediate_i_19_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_19_port);
   U3204 : MUX2_X1 port map( A => datapath_i_val_b_i_20_port, B => 
                           datapath_i_val_immediate_i_20_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_20_port);
   U3205 : MUX2_X1 port map( A => datapath_i_val_b_i_21_port, B => 
                           datapath_i_val_immediate_i_21_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_21_port);
   U3206 : MUX2_X1 port map( A => datapath_i_val_b_i_22_port, B => 
                           datapath_i_val_immediate_i_22_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_22_port);
   U3207 : MUX2_X1 port map( A => datapath_i_val_b_i_23_port, B => 
                           datapath_i_val_immediate_i_23_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_23_port);
   U3208 : MUX2_X1 port map( A => datapath_i_val_b_i_24_port, B => 
                           datapath_i_val_immediate_i_24_port, S => n3047, Z =>
                           datapath_i_execute_stage_dp_opb_24_port);
   U3209 : NAND2_X1 port map( A1 => n3047, A2 => 
                           datapath_i_val_immediate_i_25_port, ZN => n3046);
   U3210 : OAI21_X1 port map( B1 => n3047, B2 => n758, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U3211 : OAI21_X1 port map( B1 => n3047, B2 => n759, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U3212 : OAI21_X1 port map( B1 => n3047, B2 => n760, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U3213 : OAI21_X1 port map( B1 => n3047, B2 => n761, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U3214 : OAI21_X1 port map( B1 => n3047, B2 => n762, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U3215 : OAI21_X1 port map( B1 => n3047, B2 => n763, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U3216 : OAI21_X1 port map( B1 => n3047, B2 => n764, A => n3046, ZN => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U3217 : MUX2_X1 port map( A => datapath_i_val_b_i_4_port, B => 
                           datapath_i_val_immediate_i_4_port, S => n3047, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U3218 : MUX2_X1 port map( A => datapath_i_val_b_i_5_port, B => 
                           datapath_i_val_immediate_i_5_port, S => n3047, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U3219 : MUX2_X1 port map( A => datapath_i_val_b_i_6_port, B => 
                           datapath_i_val_immediate_i_6_port, S => n3047, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U3220 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_7_port, B2 => 
                           n3069, ZN => n3048);
   U3221 : OAI21_X1 port map( B1 => n705, B2 => n3084, A => n3048, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U3222 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_8_port, B2 => 
                           n3081, ZN => n3049);
   U3223 : OAI21_X1 port map( B1 => n706, B2 => n3073, A => n3049, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U3224 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_9_port, B2 => 
                           n3069, ZN => n3050);
   U3225 : OAI21_X1 port map( B1 => n707, B2 => n3084, A => n3050, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U3226 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n3081, ZN => n3051);
   U3227 : OAI21_X1 port map( B1 => n708, B2 => n3073, A => n3051, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U3228 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n3069, ZN => n3052);
   U3229 : OAI21_X1 port map( B1 => n709, B2 => n3084, A => n3052, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U3230 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n3081, ZN => n3053);
   U3231 : OAI21_X1 port map( B1 => n710, B2 => n3073, A => n3053, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U3232 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n3069, ZN => n3054);
   U3233 : OAI21_X1 port map( B1 => n711, B2 => n3084, A => n3054, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U3234 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n3081, ZN => n3055);
   U3235 : OAI21_X1 port map( B1 => n712, B2 => n3073, A => n3055, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U3236 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n3069, ZN => n3056);
   U3237 : OAI21_X1 port map( B1 => n713, B2 => n3084, A => n3056, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U3238 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n3069, ZN => n3057);
   U3239 : OAI21_X1 port map( B1 => n714, B2 => n3084, A => n3057, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U3240 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n3081, ZN => n3058);
   U3241 : OAI21_X1 port map( B1 => n715, B2 => n3084, A => n3058, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U3242 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n3069, ZN => n3059);
   U3243 : OAI21_X1 port map( B1 => n716, B2 => n3073, A => n3059, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U3244 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n3081, ZN => n3060);
   U3245 : OAI21_X1 port map( B1 => n717, B2 => n3073, A => n3060, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U3246 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n3069, ZN => n3061);
   U3247 : OAI21_X1 port map( B1 => n718, B2 => n3073, A => n3061, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U3248 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n3081, ZN => n3062);
   U3249 : OAI21_X1 port map( B1 => n719, B2 => n3073, A => n3062, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U3250 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n3069, ZN => n3063);
   U3251 : OAI21_X1 port map( B1 => n720, B2 => n3073, A => n3063, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U3252 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n3069, ZN => n3064);
   U3253 : OAI21_X1 port map( B1 => n721, B2 => n3073, A => n3064, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U3254 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n3069, ZN => n3065);
   U3255 : OAI21_X1 port map( B1 => n722, B2 => n3073, A => n3065, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U3256 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n3069, ZN => n3066);
   U3257 : OAI21_X1 port map( B1 => n723, B2 => n3073, A => n3066, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U3258 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_0_port, B2 => 
                           n3069, ZN => n3067);
   U3259 : OAI21_X1 port map( B1 => n733, B2 => n3073, A => n3067, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U3260 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n3069, ZN => n3068);
   U3261 : OAI21_X1 port map( B1 => n724, B2 => n3073, A => n3068, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U3262 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n3069, ZN => n3070);
   U3263 : OAI21_X1 port map( B1 => n725, B2 => n3073, A => n3070, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U3264 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n3071, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n3081, ZN => n3072);
   U3265 : OAI21_X1 port map( B1 => n726, B2 => n3073, A => n3072, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U3266 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n3081, ZN => n3074);
   U3267 : OAI21_X1 port map( B1 => n727, B2 => n3084, A => n3074, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U3268 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n3081, ZN => n3075);
   U3269 : OAI21_X1 port map( B1 => n703, B2 => n3084, A => n3075, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U3270 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_1_port, B2 => 
                           n3081, ZN => n3076);
   U3271 : OAI21_X1 port map( B1 => n734, B2 => n3084, A => n3076, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U3272 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_2_port, B2 => 
                           n3081, ZN => n3077);
   U3273 : OAI21_X1 port map( B1 => n728, B2 => n3084, A => n3077, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U3274 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_3_port, B2 => 
                           n3081, ZN => n3078);
   U3275 : OAI21_X1 port map( B1 => n729, B2 => n3084, A => n3078, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U3276 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_4_port, B2 => 
                           n3081, ZN => n3079);
   U3277 : OAI21_X1 port map( B1 => n730, B2 => n3084, A => n3079, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U3278 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_5_port, B2 => 
                           n3081, ZN => n3080);
   U3279 : OAI21_X1 port map( B1 => n731, B2 => n3084, A => n3080, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U3280 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n3082, B1 => datapath_i_val_a_i_6_port, B2 => 
                           n3081, ZN => n3083);
   U3281 : OAI21_X1 port map( B1 => n732, B2 => n3084, A => n3083, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);

end SYN_dlx_rtl;
